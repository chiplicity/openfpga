magic
tech EFS8A
magscale 1 2
timestamp 1602523950
<< locali >>
rect 29101 12733 29307 12767
rect 29101 12631 29135 12733
rect 12219 12393 12357 12427
rect 12115 12257 12150 12291
rect 23063 12257 23098 12291
rect 28123 11169 28250 11203
rect 35943 11169 35978 11203
rect 7935 10217 7941 10251
rect 11339 10217 11345 10251
rect 15847 10217 15853 10251
rect 17595 10217 17601 10251
rect 21275 10217 21281 10251
rect 30659 10217 30665 10251
rect 7935 10149 7969 10217
rect 11339 10149 11373 10217
rect 13035 10149 13080 10183
rect 15847 10149 15881 10217
rect 17595 10149 17629 10217
rect 21275 10149 21309 10217
rect 30659 10149 30693 10217
rect 25047 9129 25053 9163
rect 25047 9061 25081 9129
rect 32505 8993 32666 9027
rect 32505 8823 32539 8993
rect 9597 8279 9631 8449
rect 21097 8313 21281 8347
rect 33419 8041 33425 8075
rect 33419 7973 33453 8041
rect 33419 7191 33453 7259
rect 34529 7191 34563 7497
rect 33419 7157 33425 7191
rect 21275 6953 21281 6987
rect 34063 6953 34069 6987
rect 21275 6885 21309 6953
rect 34063 6885 34097 6953
rect 7389 6715 7423 6885
rect 11287 6817 11322 6851
rect 19843 6817 19878 6851
rect 29837 6647 29871 6817
rect 26893 6239 26927 6341
rect 13277 5151 13311 5321
rect 26985 5015 27019 5253
rect 23075 4777 23213 4811
rect 18739 4641 18774 4675
rect 21315 4641 21350 4675
rect 2651 4233 2789 4267
rect 19107 4029 19142 4063
rect 26249 3995 26283 4165
rect 29561 3995 29595 4165
<< viali >>
rect 21224 13345 21258 13379
rect 11529 13277 11563 13311
rect 20085 13277 20119 13311
rect 16129 13141 16163 13175
rect 21327 13141 21361 13175
rect 7067 12937 7101 12971
rect 10931 12937 10965 12971
rect 22109 12937 22143 12971
rect 25237 12937 25271 12971
rect 35633 12937 35667 12971
rect 29469 12869 29503 12903
rect 7481 12801 7515 12835
rect 16681 12801 16715 12835
rect 25697 12801 25731 12835
rect 2605 12733 2639 12767
rect 3065 12733 3099 12767
rect 6996 12733 7030 12767
rect 8769 12733 8803 12767
rect 10860 12733 10894 12767
rect 11253 12733 11287 12767
rect 14933 12733 14967 12767
rect 15393 12733 15427 12767
rect 19993 12733 20027 12767
rect 20453 12733 20487 12767
rect 21925 12733 21959 12767
rect 22477 12733 22511 12767
rect 25053 12733 25087 12767
rect 26192 12733 26226 12767
rect 26617 12733 26651 12767
rect 35449 12733 35483 12767
rect 36001 12733 36035 12767
rect 16221 12665 16255 12699
rect 16313 12665 16347 12699
rect 20729 12665 20763 12699
rect 2789 12597 2823 12631
rect 8585 12597 8619 12631
rect 8953 12597 8987 12631
rect 15117 12597 15151 12631
rect 16037 12597 16071 12631
rect 19809 12597 19843 12631
rect 21189 12597 21223 12631
rect 26295 12597 26329 12631
rect 29101 12597 29135 12631
rect 29837 12597 29871 12631
rect 12357 12393 12391 12427
rect 4215 12325 4249 12359
rect 16221 12325 16255 12359
rect 2789 12257 2823 12291
rect 4128 12257 4162 12291
rect 6561 12257 6595 12291
rect 7608 12257 7642 12291
rect 10793 12257 10827 12291
rect 10977 12257 11011 12291
rect 12081 12257 12115 12291
rect 13093 12257 13127 12291
rect 19844 12257 19878 12291
rect 22084 12257 22118 12291
rect 23029 12257 23063 12291
rect 25145 12257 25179 12291
rect 26592 12257 26626 12291
rect 27997 12257 28031 12291
rect 33736 12257 33770 12291
rect 34780 12257 34814 12291
rect 2881 12189 2915 12223
rect 8585 12189 8619 12223
rect 11069 12189 11103 12223
rect 16129 12189 16163 12223
rect 21005 12189 21039 12223
rect 16681 12121 16715 12155
rect 23167 12121 23201 12155
rect 2053 12053 2087 12087
rect 3801 12053 3835 12087
rect 6745 12053 6779 12087
rect 7711 12053 7745 12087
rect 12541 12053 12575 12087
rect 13277 12053 13311 12087
rect 19947 12053 19981 12087
rect 22155 12053 22189 12087
rect 24685 12053 24719 12087
rect 25329 12053 25363 12087
rect 26663 12053 26697 12087
rect 28181 12053 28215 12087
rect 33839 12053 33873 12087
rect 34851 12053 34885 12087
rect 8953 11849 8987 11883
rect 10609 11849 10643 11883
rect 14243 11849 14277 11883
rect 16037 11849 16071 11883
rect 21189 11849 21223 11883
rect 24501 11849 24535 11883
rect 31309 11849 31343 11883
rect 33609 11849 33643 11883
rect 35495 11849 35529 11883
rect 1685 11781 1719 11815
rect 2053 11781 2087 11815
rect 2237 11781 2271 11815
rect 3801 11781 3835 11815
rect 13461 11781 13495 11815
rect 16773 11781 16807 11815
rect 2789 11713 2823 11747
rect 9229 11713 9263 11747
rect 9873 11713 9907 11747
rect 11897 11713 11931 11747
rect 15255 11713 15289 11747
rect 16221 11713 16255 11747
rect 17509 11713 17543 11747
rect 21373 11713 21407 11747
rect 24133 11713 24167 11747
rect 2145 11645 2179 11679
rect 2421 11645 2455 11679
rect 3709 11645 3743 11679
rect 3985 11645 4019 11679
rect 7665 11645 7699 11679
rect 10977 11645 11011 11679
rect 11253 11645 11287 11679
rect 14172 11645 14206 11679
rect 15152 11645 15186 11679
rect 15577 11645 15611 11679
rect 19533 11645 19567 11679
rect 19809 11645 19843 11679
rect 20177 11645 20211 11679
rect 23740 11645 23774 11679
rect 24685 11645 24719 11679
rect 25145 11645 25179 11679
rect 26065 11645 26099 11679
rect 26525 11645 26559 11679
rect 26709 11645 26743 11679
rect 30824 11645 30858 11679
rect 33860 11645 33894 11679
rect 34253 11645 34287 11679
rect 35392 11645 35426 11679
rect 35817 11645 35851 11679
rect 6561 11577 6595 11611
rect 8309 11577 8343 11611
rect 9321 11577 9355 11611
rect 11529 11577 11563 11611
rect 12541 11577 12575 11611
rect 12633 11577 12667 11611
rect 13185 11577 13219 11611
rect 16313 11577 16347 11611
rect 18889 11577 18923 11611
rect 20453 11577 20487 11611
rect 21465 11577 21499 11611
rect 22017 11577 22051 11611
rect 23029 11577 23063 11611
rect 25421 11577 25455 11611
rect 25789 11577 25823 11611
rect 26985 11577 27019 11611
rect 3157 11509 3191 11543
rect 3525 11509 3559 11543
rect 4169 11509 4203 11543
rect 4813 11509 4847 11543
rect 5273 11509 5307 11543
rect 7481 11509 7515 11543
rect 10241 11509 10275 11543
rect 12265 11509 12299 11543
rect 14657 11509 14691 11543
rect 17141 11509 17175 11543
rect 19257 11509 19291 11543
rect 22293 11509 22327 11543
rect 23811 11509 23845 11543
rect 27353 11509 27387 11543
rect 27813 11509 27847 11543
rect 28273 11509 28307 11543
rect 30895 11509 30929 11543
rect 31769 11509 31803 11543
rect 33931 11509 33965 11543
rect 35173 11509 35207 11543
rect 3709 11305 3743 11339
rect 7665 11305 7699 11339
rect 9229 11305 9263 11339
rect 19947 11305 19981 11339
rect 23719 11305 23753 11339
rect 30389 11305 30423 11339
rect 32321 11305 32355 11339
rect 8125 11237 8159 11271
rect 8217 11237 8251 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 11989 11237 12023 11271
rect 13553 11237 13587 11271
rect 16681 11237 16715 11271
rect 17233 11237 17267 11271
rect 18245 11237 18279 11271
rect 18797 11237 18831 11271
rect 21925 11237 21959 11271
rect 26249 11237 26283 11271
rect 26617 11237 26651 11271
rect 26709 11237 26743 11271
rect 28319 11237 28353 11271
rect 34437 11237 34471 11271
rect 34529 11237 34563 11271
rect 1961 11169 1995 11203
rect 2053 11169 2087 11203
rect 2237 11169 2271 11203
rect 4077 11169 4111 11203
rect 4353 11169 4387 11203
rect 6745 11169 6779 11203
rect 6929 11169 6963 11203
rect 15520 11169 15554 11203
rect 16313 11169 16347 11203
rect 19876 11169 19910 11203
rect 23648 11169 23682 11203
rect 24777 11169 24811 11203
rect 25053 11169 25087 11203
rect 28089 11169 28123 11203
rect 30113 11169 30147 11203
rect 30573 11169 30607 11203
rect 32137 11169 32171 11203
rect 33368 11169 33402 11203
rect 35909 11169 35943 11203
rect 2421 11101 2455 11135
rect 4537 11101 4571 11135
rect 7205 11101 7239 11135
rect 8769 11101 8803 11135
rect 9781 11101 9815 11135
rect 11897 11101 11931 11135
rect 13461 11101 13495 11135
rect 13737 11101 13771 11135
rect 15623 11101 15657 11135
rect 16589 11101 16623 11135
rect 18153 11101 18187 11135
rect 21833 11101 21867 11135
rect 22477 11101 22511 11135
rect 25329 11101 25363 11135
rect 26893 11101 26927 11135
rect 4169 11033 4203 11067
rect 12449 11033 12483 11067
rect 24133 11033 24167 11067
rect 34989 11033 35023 11067
rect 35725 11033 35759 11067
rect 1685 10965 1719 10999
rect 2973 10965 3007 10999
rect 5089 10965 5123 10999
rect 10885 10965 10919 10999
rect 11161 10965 11195 10999
rect 15945 10965 15979 10999
rect 21373 10965 21407 10999
rect 25789 10965 25823 10999
rect 29837 10965 29871 10999
rect 33471 10965 33505 10999
rect 35357 10965 35391 10999
rect 36047 10965 36081 10999
rect 2329 10761 2363 10795
rect 4445 10761 4479 10795
rect 6561 10761 6595 10795
rect 9321 10761 9355 10795
rect 10517 10761 10551 10795
rect 13369 10761 13403 10795
rect 13645 10761 13679 10795
rect 14519 10761 14553 10795
rect 16313 10761 16347 10795
rect 16589 10761 16623 10795
rect 17877 10761 17911 10795
rect 19073 10761 19107 10795
rect 19763 10761 19797 10795
rect 21557 10761 21591 10795
rect 22201 10761 22235 10795
rect 31033 10761 31067 10795
rect 32965 10761 32999 10795
rect 36921 10761 36955 10795
rect 2697 10693 2731 10727
rect 2973 10693 3007 10727
rect 5365 10693 5399 10727
rect 7113 10693 7147 10727
rect 8953 10693 8987 10727
rect 10149 10693 10183 10727
rect 14013 10693 14047 10727
rect 15301 10693 15335 10727
rect 18705 10693 18739 10727
rect 19533 10693 19567 10727
rect 22707 10693 22741 10727
rect 32597 10693 32631 10727
rect 3617 10625 3651 10659
rect 4813 10625 4847 10659
rect 9597 10625 9631 10659
rect 12449 10625 12483 10659
rect 15393 10625 15427 10659
rect 16957 10625 16991 10659
rect 20637 10625 20671 10659
rect 26065 10625 26099 10659
rect 27353 10625 27387 10659
rect 27629 10625 27663 10659
rect 29837 10625 29871 10659
rect 31493 10625 31527 10659
rect 31677 10625 31711 10659
rect 32321 10625 32355 10659
rect 34989 10625 35023 10659
rect 35265 10625 35299 10659
rect 37933 10625 37967 10659
rect 1409 10557 1443 10591
rect 2881 10557 2915 10591
rect 3157 10557 3191 10591
rect 7757 10557 7791 10591
rect 11136 10557 11170 10591
rect 11621 10557 11655 10591
rect 14448 10557 14482 10591
rect 17417 10557 17451 10591
rect 19692 10557 19726 10591
rect 20085 10557 20119 10591
rect 22604 10557 22638 10591
rect 23029 10557 23063 10591
rect 23949 10557 23983 10591
rect 24133 10557 24167 10591
rect 24593 10557 24627 10591
rect 30757 10557 30791 10591
rect 33216 10557 33250 10591
rect 33977 10557 34011 10591
rect 36528 10557 36562 10591
rect 37524 10557 37558 10591
rect 4905 10489 4939 10523
rect 8078 10489 8112 10523
rect 9689 10489 9723 10523
rect 10977 10489 11011 10523
rect 12770 10489 12804 10523
rect 15755 10489 15789 10523
rect 18153 10489 18187 10523
rect 18245 10489 18279 10523
rect 20545 10489 20579 10523
rect 20999 10489 21033 10523
rect 24869 10489 24903 10523
rect 25789 10489 25823 10523
rect 25881 10489 25915 10523
rect 27077 10489 27111 10523
rect 27445 10489 27479 10523
rect 30158 10489 30192 10523
rect 31769 10489 31803 10523
rect 34345 10489 34379 10523
rect 35081 10489 35115 10523
rect 36001 10489 36035 10523
rect 37611 10489 37645 10523
rect 1593 10421 1627 10455
rect 1961 10421 1995 10455
rect 4077 10421 4111 10455
rect 7573 10421 7607 10455
rect 8677 10421 8711 10455
rect 11207 10421 11241 10455
rect 12173 10421 12207 10455
rect 14841 10421 14875 10455
rect 21833 10421 21867 10455
rect 25237 10421 25271 10455
rect 25605 10421 25639 10455
rect 26709 10421 26743 10455
rect 28273 10421 28307 10455
rect 29745 10421 29779 10455
rect 33287 10421 33321 10455
rect 33609 10421 33643 10455
rect 36599 10421 36633 10455
rect 2973 10217 3007 10251
rect 4261 10217 4295 10251
rect 4813 10217 4847 10251
rect 5825 10217 5859 10251
rect 6929 10217 6963 10251
rect 7941 10217 7975 10251
rect 8769 10217 8803 10251
rect 9505 10217 9539 10251
rect 10241 10217 10275 10251
rect 10885 10217 10919 10251
rect 11345 10217 11379 10251
rect 11897 10217 11931 10251
rect 12541 10217 12575 10251
rect 13645 10217 13679 10251
rect 15853 10217 15887 10251
rect 16405 10217 16439 10251
rect 17049 10217 17083 10251
rect 17601 10217 17635 10251
rect 18797 10217 18831 10251
rect 20637 10217 20671 10251
rect 21281 10217 21315 10251
rect 21833 10217 21867 10251
rect 24133 10217 24167 10251
rect 24593 10217 24627 10251
rect 26341 10217 26375 10251
rect 27537 10217 27571 10251
rect 30113 10217 30147 10251
rect 30665 10217 30699 10251
rect 31677 10217 31711 10251
rect 34253 10217 34287 10251
rect 35449 10217 35483 10251
rect 2329 10149 2363 10183
rect 3249 10149 3283 10183
rect 5226 10149 5260 10183
rect 13001 10149 13035 10183
rect 22845 10149 22879 10183
rect 25053 10149 25087 10183
rect 25973 10149 26007 10183
rect 26617 10149 26651 10183
rect 26709 10149 26743 10183
rect 28273 10149 28307 10183
rect 33066 10149 33100 10183
rect 34621 10149 34655 10183
rect 35173 10149 35207 10183
rect 35909 10149 35943 10183
rect 36093 10149 36127 10183
rect 36185 10149 36219 10183
rect 1685 10081 1719 10115
rect 8493 10081 8527 10115
rect 9689 10081 9723 10115
rect 10977 10081 11011 10115
rect 12173 10081 12207 10115
rect 18153 10081 18187 10115
rect 19349 10081 19383 10115
rect 19717 10081 19751 10115
rect 20913 10081 20947 10115
rect 30297 10081 30331 10115
rect 4905 10013 4939 10047
rect 7573 10013 7607 10047
rect 12725 10013 12759 10047
rect 15485 10013 15519 10047
rect 17233 10013 17267 10047
rect 19993 10013 20027 10047
rect 22753 10013 22787 10047
rect 23029 10013 23063 10047
rect 24961 10013 24995 10047
rect 25237 10013 25271 10047
rect 26893 10013 26927 10047
rect 28181 10013 28215 10047
rect 28457 10013 28491 10047
rect 32781 10013 32815 10047
rect 32965 10013 32999 10047
rect 33609 10013 33643 10047
rect 33977 10013 34011 10047
rect 34529 10013 34563 10047
rect 36369 10013 36403 10047
rect 7205 9877 7239 9911
rect 9873 9877 9907 9911
rect 14381 9877 14415 9911
rect 16681 9877 16715 9911
rect 18429 9877 18463 9911
rect 31217 9877 31251 9911
rect 2973 9673 3007 9707
rect 9781 9673 9815 9707
rect 15393 9673 15427 9707
rect 15761 9673 15795 9707
rect 17233 9673 17267 9707
rect 19855 9673 19889 9707
rect 21649 9673 21683 9707
rect 21925 9673 21959 9707
rect 22477 9673 22511 9707
rect 23397 9673 23431 9707
rect 23995 9673 24029 9707
rect 25789 9673 25823 9707
rect 26157 9673 26191 9707
rect 28181 9673 28215 9707
rect 29009 9673 29043 9707
rect 34345 9673 34379 9707
rect 36093 9673 36127 9707
rect 1961 9605 1995 9639
rect 9321 9605 9355 9639
rect 16865 9605 16899 9639
rect 19349 9605 19383 9639
rect 24409 9605 24443 9639
rect 27537 9605 27571 9639
rect 28457 9605 28491 9639
rect 31953 9605 31987 9639
rect 5549 9537 5583 9571
rect 5825 9537 5859 9571
rect 12633 9537 12667 9571
rect 13553 9537 13587 9571
rect 15117 9537 15151 9571
rect 17601 9537 17635 9571
rect 18521 9537 18555 9571
rect 20729 9537 20763 9571
rect 24869 9537 24903 9571
rect 26617 9537 26651 9571
rect 29837 9537 29871 9571
rect 33057 9537 33091 9571
rect 35265 9537 35299 9571
rect 36553 9537 36587 9571
rect 37473 9537 37507 9571
rect 1869 9469 1903 9503
rect 2145 9469 2179 9503
rect 2605 9469 2639 9503
rect 3433 9469 3467 9503
rect 3893 9469 3927 9503
rect 5089 9469 5123 9503
rect 5365 9469 5399 9503
rect 7205 9469 7239 9503
rect 7665 9469 7699 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 9137 9469 9171 9503
rect 10701 9469 10735 9503
rect 10885 9469 10919 9503
rect 12265 9469 12299 9503
rect 13093 9469 13127 9503
rect 13369 9469 13403 9503
rect 14381 9469 14415 9503
rect 14841 9469 14875 9503
rect 15945 9469 15979 9503
rect 19784 9469 19818 9503
rect 20269 9469 20303 9503
rect 22620 9469 22654 9503
rect 23924 9469 23958 9503
rect 29285 9469 29319 9503
rect 29745 9469 29779 9503
rect 31033 9469 31067 9503
rect 4353 9401 4387 9435
rect 6653 9401 6687 9435
rect 14289 9401 14323 9435
rect 16266 9401 16300 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 20637 9401 20671 9435
rect 21091 9401 21125 9435
rect 22707 9401 22741 9435
rect 25190 9401 25224 9435
rect 26938 9401 26972 9435
rect 30389 9401 30423 9435
rect 30941 9401 30975 9435
rect 31395 9401 31429 9435
rect 33149 9401 33183 9435
rect 33701 9401 33735 9435
rect 34989 9401 35023 9435
rect 35081 9401 35115 9435
rect 36645 9401 36679 9435
rect 37197 9401 37231 9435
rect 1777 9333 1811 9367
rect 3617 9333 3651 9367
rect 4721 9333 4755 9367
rect 7021 9333 7055 9367
rect 7297 9333 7331 9367
rect 9045 9333 9079 9367
rect 10241 9333 10275 9367
rect 10701 9333 10735 9367
rect 11437 9333 11471 9367
rect 11805 9333 11839 9367
rect 13921 9333 13955 9367
rect 23121 9333 23155 9367
rect 24685 9333 24719 9367
rect 26525 9333 26559 9367
rect 32413 9333 32447 9367
rect 32781 9333 32815 9367
rect 34713 9333 34747 9367
rect 1869 9129 1903 9163
rect 2237 9129 2271 9163
rect 7021 9129 7055 9163
rect 7205 9129 7239 9163
rect 8493 9129 8527 9163
rect 10517 9129 10551 9163
rect 14381 9129 14415 9163
rect 16221 9129 16255 9163
rect 21465 9129 21499 9163
rect 23857 9129 23891 9163
rect 24593 9129 24627 9163
rect 25053 9129 25087 9163
rect 25605 9129 25639 9163
rect 25881 9129 25915 9163
rect 26341 9129 26375 9163
rect 27077 9129 27111 9163
rect 29285 9129 29319 9163
rect 31125 9129 31159 9163
rect 34529 9129 34563 9163
rect 34989 9129 35023 9163
rect 36277 9129 36311 9163
rect 36645 9129 36679 9163
rect 4261 9061 4295 9095
rect 4813 9061 4847 9095
rect 11206 9061 11240 9095
rect 12817 9061 12851 9095
rect 15663 9061 15697 9095
rect 17509 9061 17543 9095
rect 19441 9061 19475 9095
rect 21925 9061 21959 9095
rect 27813 9061 27847 9095
rect 27905 9061 27939 9095
rect 30291 9061 30325 9095
rect 33971 9061 34005 9095
rect 35719 9061 35753 9095
rect 1409 8993 1443 9027
rect 2421 8993 2455 9027
rect 2973 8993 3007 9027
rect 5733 8993 5767 9027
rect 5917 8993 5951 9027
rect 7205 8993 7239 9027
rect 7573 8993 7607 9027
rect 7941 8993 7975 9027
rect 11805 8993 11839 9027
rect 14197 8993 14231 9027
rect 23673 8993 23707 9027
rect 26560 8993 26594 9027
rect 27445 8993 27479 9027
rect 30849 8993 30883 9027
rect 36921 8993 36955 9027
rect 3157 8925 3191 8959
rect 4169 8925 4203 8959
rect 9873 8925 9907 8959
rect 10885 8925 10919 8959
rect 12725 8925 12759 8959
rect 15301 8925 15335 8959
rect 17417 8925 17451 8959
rect 17693 8925 17727 8959
rect 19349 8925 19383 8959
rect 21833 8925 21867 8959
rect 24685 8925 24719 8959
rect 28089 8925 28123 8959
rect 29929 8925 29963 8959
rect 1593 8857 1627 8891
rect 13277 8857 13311 8891
rect 19901 8857 19935 8891
rect 22385 8857 22419 8891
rect 33609 8925 33643 8959
rect 35357 8925 35391 8959
rect 3893 8789 3927 8823
rect 5181 8789 5215 8823
rect 6009 8789 6043 8823
rect 15117 8789 15151 8823
rect 16497 8789 16531 8823
rect 17233 8789 17267 8823
rect 18613 8789 18647 8823
rect 19073 8789 19107 8823
rect 21189 8789 21223 8823
rect 24133 8789 24167 8823
rect 26663 8789 26697 8823
rect 31493 8789 31527 8823
rect 32505 8789 32539 8823
rect 32735 8789 32769 8823
rect 33333 8789 33367 8823
rect 1593 8585 1627 8619
rect 3985 8585 4019 8619
rect 7021 8585 7055 8619
rect 8033 8585 8067 8619
rect 11253 8585 11287 8619
rect 11805 8585 11839 8619
rect 12173 8585 12207 8619
rect 14473 8585 14507 8619
rect 17509 8585 17543 8619
rect 17785 8585 17819 8619
rect 21465 8585 21499 8619
rect 23029 8585 23063 8619
rect 26525 8585 26559 8619
rect 28273 8585 28307 8619
rect 29009 8585 29043 8619
rect 32321 8585 32355 8619
rect 32689 8585 32723 8619
rect 36277 8585 36311 8619
rect 5365 8517 5399 8551
rect 10977 8517 11011 8551
rect 14197 8517 14231 8551
rect 17141 8517 17175 8551
rect 19533 8517 19567 8551
rect 21741 8517 21775 8551
rect 22569 8517 22603 8551
rect 23489 8517 23523 8551
rect 34345 8517 34379 8551
rect 35541 8517 35575 8551
rect 8125 8449 8159 8483
rect 9597 8449 9631 8483
rect 9965 8449 9999 8483
rect 10241 8449 10275 8483
rect 15393 8449 15427 8483
rect 16221 8449 16255 8483
rect 19809 8449 19843 8483
rect 23765 8449 23799 8483
rect 24041 8449 24075 8483
rect 25329 8449 25363 8483
rect 27077 8449 27111 8483
rect 30573 8449 30607 8483
rect 33333 8449 33367 8483
rect 34989 8449 35023 8483
rect 36829 8449 36863 8483
rect 1409 8381 1443 8415
rect 2697 8381 2731 8415
rect 4445 8381 4479 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 9045 8381 9079 8415
rect 2605 8313 2639 8347
rect 3059 8313 3093 8347
rect 4766 8313 4800 8347
rect 5825 8313 5859 8347
rect 8446 8313 8480 8347
rect 13001 8381 13035 8415
rect 13369 8381 13403 8415
rect 13553 8381 13587 8415
rect 14657 8381 14691 8415
rect 15117 8381 15151 8415
rect 18613 8381 18647 8415
rect 29837 8381 29871 8415
rect 30297 8381 30331 8415
rect 30941 8381 30975 8415
rect 31401 8381 31435 8415
rect 10057 8313 10091 8347
rect 13829 8313 13863 8347
rect 15761 8313 15795 8347
rect 16129 8313 16163 8347
rect 16583 8313 16617 8347
rect 18934 8313 18968 8347
rect 20453 8313 20487 8347
rect 20545 8313 20579 8347
rect 21281 8313 21315 8347
rect 22017 8313 22051 8347
rect 22109 8313 22143 8347
rect 23857 8313 23891 8347
rect 24777 8313 24811 8347
rect 25237 8313 25271 8347
rect 25691 8313 25725 8347
rect 27398 8313 27432 8347
rect 31763 8313 31797 8347
rect 33425 8313 33459 8347
rect 33977 8313 34011 8347
rect 34713 8313 34747 8347
rect 35081 8313 35115 8347
rect 36553 8313 36587 8347
rect 36645 8313 36679 8347
rect 2053 8245 2087 8279
rect 3617 8245 3651 8279
rect 4353 8245 4387 8279
rect 6193 8245 6227 8279
rect 7389 8245 7423 8279
rect 9321 8245 9355 8279
rect 9597 8245 9631 8279
rect 9781 8245 9815 8279
rect 18521 8245 18555 8279
rect 20269 8245 20303 8279
rect 26249 8245 26283 8279
rect 26985 8245 27019 8279
rect 27997 8245 28031 8279
rect 29745 8245 29779 8279
rect 31309 8245 31343 8279
rect 33057 8245 33091 8279
rect 35909 8245 35943 8279
rect 37473 8245 37507 8279
rect 1961 8041 1995 8075
rect 2697 8041 2731 8075
rect 3433 8041 3467 8075
rect 3893 8041 3927 8075
rect 5089 8041 5123 8075
rect 7205 8041 7239 8075
rect 12633 8041 12667 8075
rect 15485 8041 15519 8075
rect 19625 8041 19659 8075
rect 25421 8041 25455 8075
rect 27813 8041 27847 8075
rect 28825 8041 28859 8075
rect 30021 8041 30055 8075
rect 32965 8041 32999 8075
rect 33425 8041 33459 8075
rect 36645 8041 36679 8075
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 10149 7973 10183 8007
rect 11345 7973 11379 8007
rect 13230 7973 13264 8007
rect 14657 7973 14691 8007
rect 16589 7973 16623 8007
rect 19026 7973 19060 8007
rect 19993 7973 20027 8007
rect 21097 7973 21131 8007
rect 21925 7973 21959 8007
rect 22661 7973 22695 8007
rect 23765 7973 23799 8007
rect 24133 7973 24167 8007
rect 24225 7973 24259 8007
rect 26709 7973 26743 8007
rect 29653 7973 29687 8007
rect 30297 7973 30331 8007
rect 31217 7973 31251 8007
rect 35081 7973 35115 8007
rect 1409 7905 1443 7939
rect 2329 7905 2363 7939
rect 2697 7905 2731 7939
rect 2973 7905 3007 7939
rect 6193 7905 6227 7939
rect 7665 7905 7699 7939
rect 11529 7905 11563 7939
rect 11713 7905 11747 7939
rect 15853 7905 15887 7939
rect 16313 7905 16347 7939
rect 16865 7905 16899 7939
rect 17417 7905 17451 7939
rect 22293 7905 22327 7939
rect 28917 7905 28951 7939
rect 29377 7905 29411 7939
rect 30481 7905 30515 7939
rect 30941 7905 30975 7939
rect 36461 7905 36495 7939
rect 4169 7837 4203 7871
rect 6837 7837 6871 7871
rect 8033 7837 8067 7871
rect 8769 7837 8803 7871
rect 10057 7837 10091 7871
rect 10333 7837 10367 7871
rect 12909 7837 12943 7871
rect 18705 7837 18739 7871
rect 21005 7837 21039 7871
rect 21649 7837 21683 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 24409 7837 24443 7871
rect 26617 7837 26651 7871
rect 27261 7837 27295 7871
rect 33057 7837 33091 7871
rect 34437 7837 34471 7871
rect 34989 7837 35023 7871
rect 1593 7769 1627 7803
rect 7803 7769 7837 7803
rect 20453 7769 20487 7803
rect 35541 7769 35575 7803
rect 7481 7701 7515 7735
rect 7941 7701 7975 7735
rect 8309 7701 8343 7735
rect 9229 7701 9263 7735
rect 10977 7701 11011 7735
rect 11805 7701 11839 7735
rect 13829 7701 13863 7735
rect 17601 7701 17635 7735
rect 33977 7701 34011 7735
rect 34805 7701 34839 7735
rect 1777 7497 1811 7531
rect 3433 7497 3467 7531
rect 5549 7497 5583 7531
rect 5871 7497 5905 7531
rect 9689 7497 9723 7531
rect 15853 7497 15887 7531
rect 18245 7497 18279 7531
rect 19993 7497 20027 7531
rect 20913 7497 20947 7531
rect 22477 7497 22511 7531
rect 23121 7497 23155 7531
rect 26801 7497 26835 7531
rect 29101 7497 29135 7531
rect 30481 7497 30515 7531
rect 34529 7497 34563 7531
rect 34621 7497 34655 7531
rect 6193 7429 6227 7463
rect 7941 7429 7975 7463
rect 8677 7429 8711 7463
rect 9137 7429 9171 7463
rect 9505 7429 9539 7463
rect 14473 7429 14507 7463
rect 17785 7429 17819 7463
rect 23397 7429 23431 7463
rect 32045 7429 32079 7463
rect 33977 7429 34011 7463
rect 6653 7361 6687 7395
rect 8033 7361 8067 7395
rect 8401 7361 8435 7395
rect 9597 7361 9631 7395
rect 11529 7361 11563 7395
rect 11805 7361 11839 7395
rect 15209 7361 15243 7395
rect 17141 7361 17175 7395
rect 18613 7361 18647 7395
rect 18981 7361 19015 7395
rect 27445 7361 27479 7395
rect 27721 7361 27755 7395
rect 2237 7293 2271 7327
rect 3985 7293 4019 7327
rect 5181 7293 5215 7327
rect 5800 7293 5834 7327
rect 7812 7293 7846 7327
rect 9376 7293 9410 7327
rect 11069 7293 11103 7327
rect 11253 7293 11287 7327
rect 12449 7293 12483 7327
rect 13645 7293 13679 7327
rect 14657 7293 14691 7327
rect 15117 7293 15151 7327
rect 16313 7293 16347 7327
rect 16681 7293 16715 7327
rect 16865 7293 16899 7327
rect 18061 7293 18095 7327
rect 19073 7293 19107 7327
rect 24041 7293 24075 7327
rect 24501 7293 24535 7327
rect 25145 7293 25179 7327
rect 25605 7293 25639 7327
rect 29285 7293 29319 7327
rect 29745 7293 29779 7327
rect 31125 7293 31159 7327
rect 33057 7293 33091 7327
rect 34253 7293 34287 7327
rect 2145 7225 2179 7259
rect 2558 7225 2592 7259
rect 3801 7225 3835 7259
rect 4347 7225 4381 7259
rect 7665 7225 7699 7259
rect 9229 7225 9263 7259
rect 10241 7225 10275 7259
rect 12770 7225 12804 7259
rect 14013 7225 14047 7259
rect 19435 7225 19469 7259
rect 21189 7225 21223 7259
rect 21281 7225 21315 7259
rect 21833 7225 21867 7259
rect 25926 7225 25960 7259
rect 27537 7225 27571 7259
rect 31033 7225 31067 7259
rect 31487 7225 31521 7259
rect 35909 7429 35943 7463
rect 34989 7361 35023 7395
rect 36829 7361 36863 7395
rect 35081 7225 35115 7259
rect 35633 7225 35667 7259
rect 36553 7225 36587 7259
rect 36645 7225 36679 7259
rect 3157 7157 3191 7191
rect 4905 7157 4939 7191
rect 7205 7157 7239 7191
rect 7481 7157 7515 7191
rect 10701 7157 10735 7191
rect 12173 7157 12207 7191
rect 13369 7157 13403 7191
rect 17417 7157 17451 7191
rect 20637 7157 20671 7191
rect 22109 7157 22143 7191
rect 23949 7157 23983 7191
rect 24133 7157 24167 7191
rect 25513 7157 25547 7191
rect 26525 7157 26559 7191
rect 27169 7157 27203 7191
rect 28641 7157 28675 7191
rect 29561 7157 29595 7191
rect 32597 7157 32631 7191
rect 32965 7157 32999 7191
rect 33425 7157 33459 7191
rect 34529 7157 34563 7191
rect 36277 7157 36311 7191
rect 1869 6953 1903 6987
rect 14243 6953 14277 6987
rect 15945 6953 15979 6987
rect 19947 6953 19981 6987
rect 20361 6953 20395 6987
rect 21281 6953 21315 6987
rect 21833 6953 21867 6987
rect 22753 6953 22787 6987
rect 24409 6953 24443 6987
rect 26249 6953 26283 6987
rect 27537 6953 27571 6987
rect 31493 6953 31527 6987
rect 32229 6953 32263 6987
rect 33241 6953 33275 6987
rect 34069 6953 34103 6987
rect 34989 6953 35023 6987
rect 36369 6953 36403 6987
rect 2605 6885 2639 6919
rect 4261 6885 4295 6919
rect 7389 6885 7423 6919
rect 8769 6885 8803 6919
rect 10885 6885 10919 6919
rect 11713 6885 11747 6919
rect 12678 6885 12712 6919
rect 16450 6885 16484 6919
rect 18613 6885 18647 6919
rect 18889 6885 18923 6919
rect 25053 6885 25087 6919
rect 26709 6885 26743 6919
rect 27261 6885 27295 6919
rect 30849 6885 30883 6919
rect 35811 6885 35845 6919
rect 1409 6817 1443 6851
rect 5641 6817 5675 6851
rect 6193 6817 6227 6851
rect 2513 6749 2547 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 6009 6749 6043 6783
rect 7757 6817 7791 6851
rect 9965 6817 9999 6851
rect 11253 6817 11287 6851
rect 14172 6817 14206 6851
rect 17877 6817 17911 6851
rect 18337 6817 18371 6851
rect 19809 6817 19843 6851
rect 22845 6817 22879 6851
rect 23121 6817 23155 6851
rect 28825 6817 28859 6851
rect 29009 6817 29043 6851
rect 29561 6817 29595 6851
rect 29837 6817 29871 6851
rect 30389 6817 30423 6851
rect 30665 6817 30699 6851
rect 32137 6817 32171 6851
rect 32597 6817 32631 6851
rect 36645 6817 36679 6851
rect 8125 6749 8159 6783
rect 9229 6749 9263 6783
rect 12357 6749 12391 6783
rect 16129 6749 16163 6783
rect 20913 6749 20947 6783
rect 24041 6749 24075 6783
rect 24961 6749 24995 6783
rect 25605 6749 25639 6783
rect 26617 6749 26651 6783
rect 29285 6749 29319 6783
rect 3065 6681 3099 6715
rect 7389 6681 7423 6715
rect 7922 6681 7956 6715
rect 31125 6749 31159 6783
rect 33701 6749 33735 6783
rect 35449 6749 35483 6783
rect 33517 6681 33551 6715
rect 34621 6681 34655 6715
rect 35265 6681 35299 6715
rect 1593 6613 1627 6647
rect 2237 6613 2271 6647
rect 3433 6613 3467 6647
rect 3801 6613 3835 6647
rect 6929 6613 6963 6647
rect 7205 6613 7239 6647
rect 7573 6613 7607 6647
rect 8033 6613 8067 6647
rect 8401 6613 8435 6647
rect 10149 6613 10183 6647
rect 11391 6613 11425 6647
rect 12173 6613 12207 6647
rect 13277 6613 13311 6647
rect 14749 6613 14783 6647
rect 17049 6613 17083 6647
rect 19257 6613 19291 6647
rect 20637 6613 20671 6647
rect 22109 6613 22143 6647
rect 23765 6613 23799 6647
rect 29837 6613 29871 6647
rect 30021 6613 30055 6647
rect 1593 6409 1627 6443
rect 2513 6409 2547 6443
rect 3617 6409 3651 6443
rect 5641 6409 5675 6443
rect 7941 6409 7975 6443
rect 9413 6409 9447 6443
rect 12173 6409 12207 6443
rect 13645 6409 13679 6443
rect 15577 6409 15611 6443
rect 15945 6409 15979 6443
rect 17417 6409 17451 6443
rect 19947 6409 19981 6443
rect 21833 6409 21867 6443
rect 24961 6409 24995 6443
rect 26341 6409 26375 6443
rect 28181 6409 28215 6443
rect 28641 6409 28675 6443
rect 29745 6409 29779 6443
rect 32505 6409 32539 6443
rect 34253 6409 34287 6443
rect 35909 6409 35943 6443
rect 36645 6409 36679 6443
rect 37105 6409 37139 6443
rect 4077 6341 4111 6375
rect 4813 6341 4847 6375
rect 5917 6341 5951 6375
rect 26893 6341 26927 6375
rect 26985 6341 27019 6375
rect 32781 6341 32815 6375
rect 35541 6341 35575 6375
rect 2697 6273 2731 6307
rect 3341 6273 3375 6307
rect 6653 6273 6687 6307
rect 10057 6273 10091 6307
rect 11253 6273 11287 6307
rect 14105 6273 14139 6307
rect 14657 6273 14691 6307
rect 17785 6273 17819 6307
rect 18429 6273 18463 6307
rect 20361 6273 20395 6307
rect 21373 6273 21407 6307
rect 26617 6273 26651 6307
rect 28917 6273 28951 6307
rect 31217 6273 31251 6307
rect 33241 6273 33275 6307
rect 33701 6273 33735 6307
rect 36277 6273 36311 6307
rect 1409 6205 1443 6239
rect 5733 6205 5767 6239
rect 6837 6205 6871 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 8493 6205 8527 6239
rect 11897 6205 11931 6239
rect 12449 6205 12483 6239
rect 16037 6205 16071 6239
rect 19876 6205 19910 6239
rect 22636 6205 22670 6239
rect 23029 6205 23063 6239
rect 23857 6205 23891 6239
rect 24133 6205 24167 6239
rect 25421 6205 25455 6239
rect 26893 6205 26927 6239
rect 27169 6205 27203 6239
rect 27629 6205 27663 6239
rect 31493 6205 31527 6239
rect 31861 6205 31895 6239
rect 36461 6205 36495 6239
rect 37616 6205 37650 6239
rect 38025 6205 38059 6239
rect 2789 6137 2823 6171
rect 4261 6137 4295 6171
rect 4353 6137 4387 6171
rect 10149 6137 10183 6171
rect 10701 6137 10735 6171
rect 12770 6137 12804 6171
rect 14289 6137 14323 6171
rect 14381 6137 14415 6171
rect 16358 6137 16392 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 19073 6137 19107 6171
rect 20913 6137 20947 6171
rect 21005 6137 21039 6171
rect 23489 6137 23523 6171
rect 25329 6137 25363 6171
rect 25783 6137 25817 6171
rect 29929 6137 29963 6171
rect 30021 6137 30055 6171
rect 30573 6137 30607 6171
rect 32137 6137 32171 6171
rect 33333 6137 33367 6171
rect 34713 6137 34747 6171
rect 34989 6137 35023 6171
rect 35081 6137 35115 6171
rect 37703 6137 37737 6171
rect 2053 6069 2087 6103
rect 5181 6069 5215 6103
rect 6193 6069 6227 6103
rect 7297 6069 7331 6103
rect 8217 6069 8251 6103
rect 8677 6069 8711 6103
rect 9873 6069 9907 6103
rect 13369 6069 13403 6103
rect 16957 6069 16991 6103
rect 20637 6069 20671 6103
rect 22385 6069 22419 6103
rect 22707 6069 22741 6103
rect 23765 6069 23799 6103
rect 27261 6069 27295 6103
rect 30941 6069 30975 6103
rect 1593 5865 1627 5899
rect 2881 5865 2915 5899
rect 3249 5865 3283 5899
rect 3617 5865 3651 5899
rect 4215 5865 4249 5899
rect 4537 5865 4571 5899
rect 5641 5865 5675 5899
rect 6561 5865 6595 5899
rect 9505 5865 9539 5899
rect 11161 5865 11195 5899
rect 12449 5865 12483 5899
rect 14197 5865 14231 5899
rect 18613 5865 18647 5899
rect 24869 5865 24903 5899
rect 26709 5865 26743 5899
rect 34069 5865 34103 5899
rect 6837 5797 6871 5831
rect 8953 5797 8987 5831
rect 10241 5797 10275 5831
rect 10793 5797 10827 5831
rect 13185 5797 13219 5831
rect 15485 5797 15519 5831
rect 17785 5797 17819 5831
rect 19993 5797 20027 5831
rect 20637 5797 20671 5831
rect 21189 5797 21223 5831
rect 21827 5797 21861 5831
rect 23575 5797 23609 5831
rect 27439 5797 27473 5831
rect 29790 5797 29824 5831
rect 32642 5797 32676 5831
rect 34621 5797 34655 5831
rect 1961 5729 1995 5763
rect 4144 5729 4178 5763
rect 6009 5729 6043 5763
rect 7849 5729 7883 5763
rect 8401 5729 8435 5763
rect 11621 5729 11655 5763
rect 11805 5729 11839 5763
rect 19257 5729 19291 5763
rect 19809 5729 19843 5763
rect 21465 5729 21499 5763
rect 23213 5729 23247 5763
rect 25028 5729 25062 5763
rect 27077 5729 27111 5763
rect 29469 5729 29503 5763
rect 32321 5729 32355 5763
rect 36036 5729 36070 5763
rect 8309 5661 8343 5695
rect 8677 5661 8711 5695
rect 10149 5661 10183 5695
rect 13093 5661 13127 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17509 5661 17543 5695
rect 17693 5661 17727 5695
rect 34529 5661 34563 5695
rect 34805 5661 34839 5695
rect 2145 5593 2179 5627
rect 13645 5593 13679 5627
rect 18245 5593 18279 5627
rect 30665 5593 30699 5627
rect 4905 5525 4939 5559
rect 7389 5525 7423 5559
rect 9965 5525 9999 5559
rect 11897 5525 11931 5559
rect 12909 5525 12943 5559
rect 16313 5525 16347 5559
rect 16681 5525 16715 5559
rect 22385 5525 22419 5559
rect 24133 5525 24167 5559
rect 24409 5525 24443 5559
rect 25099 5525 25133 5559
rect 25513 5525 25547 5559
rect 27997 5525 28031 5559
rect 30389 5525 30423 5559
rect 31493 5525 31527 5559
rect 33241 5525 33275 5559
rect 33701 5525 33735 5559
rect 36139 5525 36173 5559
rect 3157 5321 3191 5355
rect 5457 5321 5491 5355
rect 6285 5321 6319 5355
rect 9229 5321 9263 5355
rect 10609 5321 10643 5355
rect 11989 5321 12023 5355
rect 13093 5321 13127 5355
rect 13277 5321 13311 5355
rect 14841 5321 14875 5355
rect 15117 5321 15151 5355
rect 17417 5321 17451 5355
rect 17877 5321 17911 5355
rect 19257 5321 19291 5355
rect 19717 5321 19751 5355
rect 20039 5321 20073 5355
rect 20821 5321 20855 5355
rect 21925 5321 21959 5355
rect 23305 5321 23339 5355
rect 25053 5321 25087 5355
rect 26801 5321 26835 5355
rect 28733 5321 28767 5355
rect 30389 5321 30423 5355
rect 34529 5321 34563 5355
rect 36047 5321 36081 5355
rect 36737 5321 36771 5355
rect 4997 5253 5031 5287
rect 10333 5253 10367 5287
rect 12679 5253 12713 5287
rect 4629 5185 4663 5219
rect 7297 5185 7331 5219
rect 8861 5185 8895 5219
rect 15485 5253 15519 5287
rect 21097 5253 21131 5287
rect 22661 5253 22695 5287
rect 26985 5253 27019 5287
rect 28273 5253 28307 5287
rect 36461 5253 36495 5287
rect 13645 5185 13679 5219
rect 14289 5185 14323 5219
rect 16773 5185 16807 5219
rect 18797 5185 18831 5219
rect 23765 5185 23799 5219
rect 25329 5185 25363 5219
rect 25605 5185 25639 5219
rect 2421 5117 2455 5151
rect 2697 5117 2731 5151
rect 3985 5117 4019 5151
rect 5733 5117 5767 5151
rect 7757 5117 7791 5151
rect 8125 5117 8159 5151
rect 8309 5117 8343 5151
rect 8585 5117 8619 5151
rect 9413 5117 9447 5151
rect 11212 5117 11246 5151
rect 12608 5117 12642 5151
rect 13277 5117 13311 5151
rect 15289 5117 15323 5151
rect 15853 5117 15887 5151
rect 18061 5117 18095 5151
rect 18521 5117 18555 5151
rect 19947 5117 19981 5151
rect 20913 5117 20947 5151
rect 21465 5117 21499 5151
rect 3709 5049 3743 5083
rect 6653 5049 6687 5083
rect 9734 5049 9768 5083
rect 11299 5049 11333 5083
rect 13737 5049 13771 5083
rect 16497 5049 16531 5083
rect 16589 5049 16623 5083
rect 20361 5049 20395 5083
rect 22109 5049 22143 5083
rect 22201 5049 22235 5083
rect 23857 5049 23891 5083
rect 24409 5049 24443 5083
rect 25421 5049 25455 5083
rect 29009 5185 29043 5219
rect 29469 5185 29503 5219
rect 30665 5185 30699 5219
rect 31125 5185 31159 5219
rect 33517 5185 33551 5219
rect 34897 5185 34931 5219
rect 27169 5117 27203 5151
rect 31217 5117 31251 5151
rect 31769 5117 31803 5151
rect 35976 5117 36010 5151
rect 27721 5049 27755 5083
rect 27813 5049 27847 5083
rect 29790 5049 29824 5083
rect 32321 5049 32355 5083
rect 33057 5049 33091 5083
rect 33241 5049 33275 5083
rect 33333 5049 33367 5083
rect 1869 4981 1903 5015
rect 2237 4981 2271 5015
rect 5917 4981 5951 5015
rect 11713 4981 11747 5015
rect 13461 4981 13495 5015
rect 16313 4981 16347 5015
rect 26985 4981 27019 5015
rect 27445 4981 27479 5015
rect 31309 4981 31343 5015
rect 5089 4777 5123 4811
rect 6193 4777 6227 4811
rect 8677 4777 8711 4811
rect 9413 4777 9447 4811
rect 10149 4777 10183 4811
rect 11713 4777 11747 4811
rect 12081 4777 12115 4811
rect 12725 4777 12759 4811
rect 13093 4777 13127 4811
rect 16497 4777 16531 4811
rect 18245 4777 18279 4811
rect 18843 4777 18877 4811
rect 21419 4777 21453 4811
rect 22385 4777 22419 4811
rect 23213 4777 23247 4811
rect 23857 4777 23891 4811
rect 25605 4777 25639 4811
rect 27031 4777 27065 4811
rect 27629 4777 27663 4811
rect 29469 4777 29503 4811
rect 31217 4777 31251 4811
rect 31953 4777 31987 4811
rect 33241 4777 33275 4811
rect 34437 4777 34471 4811
rect 2973 4709 3007 4743
rect 5917 4709 5951 4743
rect 8401 4709 8435 4743
rect 10793 4709 10827 4743
rect 12311 4709 12345 4743
rect 13369 4709 13403 4743
rect 13921 4709 13955 4743
rect 16037 4709 16071 4743
rect 17325 4709 17359 4743
rect 19947 4709 19981 4743
rect 23489 4709 23523 4743
rect 24133 4709 24167 4743
rect 25237 4709 25271 4743
rect 28089 4709 28123 4743
rect 29929 4709 29963 4743
rect 30481 4709 30515 4743
rect 32873 4709 32907 4743
rect 2513 4641 2547 4675
rect 2789 4641 2823 4675
rect 4905 4641 4939 4675
rect 6101 4641 6135 4675
rect 7297 4641 7331 4675
rect 7573 4641 7607 4675
rect 12224 4641 12258 4675
rect 15485 4641 15519 4675
rect 15853 4641 15887 4675
rect 18705 4641 18739 4675
rect 19844 4641 19878 4675
rect 21281 4641 21315 4675
rect 22109 4641 22143 4675
rect 23004 4641 23038 4675
rect 26960 4641 26994 4675
rect 32137 4641 32171 4675
rect 32597 4641 32631 4675
rect 33701 4641 33735 4675
rect 34748 4641 34782 4675
rect 7757 4573 7791 4607
rect 10701 4573 10735 4607
rect 13277 4573 13311 4607
rect 17233 4573 17267 4607
rect 17601 4573 17635 4607
rect 24041 4573 24075 4607
rect 24409 4573 24443 4607
rect 27997 4573 28031 4607
rect 28273 4573 28307 4607
rect 29837 4573 29871 4607
rect 7389 4505 7423 4539
rect 11253 4505 11287 4539
rect 7205 4437 7239 4471
rect 14197 4437 14231 4471
rect 34851 4437 34885 4471
rect 1593 4233 1627 4267
rect 2421 4233 2455 4267
rect 2789 4233 2823 4267
rect 3065 4233 3099 4267
rect 3663 4233 3697 4267
rect 4905 4233 4939 4267
rect 5273 4233 5307 4267
rect 7021 4233 7055 4267
rect 8033 4233 8067 4267
rect 12265 4233 12299 4267
rect 13461 4233 13495 4267
rect 17509 4233 17543 4267
rect 18199 4233 18233 4267
rect 19211 4233 19245 4267
rect 19809 4233 19843 4267
rect 21649 4233 21683 4267
rect 23489 4233 23523 4267
rect 23811 4233 23845 4267
rect 26433 4233 26467 4267
rect 27629 4233 27663 4267
rect 27905 4233 27939 4267
rect 28227 4233 28261 4267
rect 29009 4233 29043 4267
rect 35081 4233 35115 4267
rect 9965 4165 9999 4199
rect 15393 4165 15427 4199
rect 16589 4165 16623 4199
rect 25973 4165 26007 4199
rect 26249 4165 26283 4199
rect 29469 4165 29503 4199
rect 29561 4165 29595 4199
rect 3985 4097 4019 4131
rect 8585 4097 8619 4131
rect 11253 4097 11287 4131
rect 13001 4097 13035 4131
rect 14565 4097 14599 4131
rect 16313 4097 16347 4131
rect 17233 4097 17267 4131
rect 18889 4097 18923 4131
rect 21281 4097 21315 4131
rect 25513 4097 25547 4131
rect 1409 4029 1443 4063
rect 2580 4029 2614 4063
rect 3592 4029 3626 4063
rect 5365 4029 5399 4063
rect 5549 4029 5583 4063
rect 6193 4029 6227 4063
rect 6561 4029 6595 4063
rect 7389 4029 7423 4063
rect 9505 4029 9539 4063
rect 12725 4029 12759 4063
rect 12909 4029 12943 4063
rect 14013 4029 14047 4063
rect 14473 4029 14507 4063
rect 15577 4029 15611 4063
rect 16037 4029 16071 4063
rect 18128 4029 18162 4063
rect 19073 4029 19107 4063
rect 21465 4029 21499 4063
rect 21925 4029 21959 4063
rect 23740 4029 23774 4063
rect 24869 4029 24903 4063
rect 25237 4029 25271 4063
rect 25421 4029 25455 4063
rect 26525 4029 26559 4063
rect 26985 4029 27019 4063
rect 28124 4029 28158 4063
rect 28549 4029 28583 4063
rect 29285 4029 29319 4063
rect 5917 3961 5951 3995
rect 7205 3961 7239 3995
rect 8401 3961 8435 3995
rect 8906 3961 8940 3995
rect 10333 3961 10367 3995
rect 10885 3961 10919 3995
rect 10977 3961 11011 3995
rect 13921 3961 13955 3995
rect 15117 3961 15151 3995
rect 26249 3961 26283 3995
rect 30205 4097 30239 4131
rect 31401 4097 31435 4131
rect 31769 4097 31803 4131
rect 32137 4097 32171 4131
rect 32965 4097 32999 4131
rect 29745 4029 29779 4063
rect 30665 4029 30699 4063
rect 31217 4029 31251 4063
rect 32505 4029 32539 4063
rect 32689 4029 32723 4063
rect 29561 3961 29595 3995
rect 30573 3961 30607 3995
rect 2053 3893 2087 3927
rect 7481 3893 7515 3927
rect 10609 3893 10643 3927
rect 11897 3893 11931 3927
rect 18613 3893 18647 3927
rect 23029 3893 23063 3927
rect 24225 3893 24259 3927
rect 26617 3893 26651 3927
rect 2697 3689 2731 3723
rect 6009 3689 6043 3723
rect 6561 3689 6595 3723
rect 6929 3689 6963 3723
rect 7205 3689 7239 3723
rect 10609 3689 10643 3723
rect 11345 3689 11379 3723
rect 12173 3689 12207 3723
rect 12909 3689 12943 3723
rect 13277 3689 13311 3723
rect 13461 3689 13495 3723
rect 14013 3689 14047 3723
rect 15669 3689 15703 3723
rect 16037 3689 16071 3723
rect 16911 3689 16945 3723
rect 17923 3689 17957 3723
rect 19165 3689 19199 3723
rect 24041 3689 24075 3723
rect 24961 3689 24995 3723
rect 27997 3689 28031 3723
rect 29837 3689 29871 3723
rect 32321 3689 32355 3723
rect 32689 3689 32723 3723
rect 2283 3621 2317 3655
rect 7757 3621 7791 3655
rect 31125 3621 31159 3655
rect 2196 3553 2230 3587
rect 6377 3553 6411 3587
rect 10793 3553 10827 3587
rect 12173 3553 12207 3587
rect 12357 3553 12391 3587
rect 15485 3553 15519 3587
rect 16808 3553 16842 3587
rect 17820 3553 17854 3587
rect 30665 3553 30699 3587
rect 30941 3553 30975 3587
rect 8125 3485 8159 3519
rect 7573 3417 7607 3451
rect 8033 3417 8067 3451
rect 7895 3349 7929 3383
rect 8217 3349 8251 3383
rect 2237 3145 2271 3179
rect 6377 3145 6411 3179
rect 7297 3145 7331 3179
rect 8217 3145 8251 3179
rect 8585 3145 8619 3179
rect 9781 3145 9815 3179
rect 10517 3145 10551 3179
rect 11529 3145 11563 3179
rect 14151 3145 14185 3179
rect 15485 3145 15519 3179
rect 15853 3145 15887 3179
rect 30757 3145 30791 3179
rect 10149 3077 10183 3111
rect 16773 3077 16807 3111
rect 17785 3077 17819 3111
rect 30481 3077 30515 3111
rect 10609 3009 10643 3043
rect 13001 3009 13035 3043
rect 7389 2941 7423 2975
rect 9597 2941 9631 2975
rect 12725 2941 12759 2975
rect 12909 2941 12943 2975
rect 14048 2941 14082 2975
rect 14473 2941 14507 2975
rect 15669 2941 15703 2975
rect 16129 2941 16163 2975
rect 7849 2873 7883 2907
rect 7573 2805 7607 2839
rect 11805 2805 11839 2839
rect 12173 2805 12207 2839
rect 7757 2601 7791 2635
rect 10425 2601 10459 2635
rect 10793 2601 10827 2635
rect 13277 2601 13311 2635
rect 28825 2601 28859 2635
rect 10241 2465 10275 2499
rect 11564 2465 11598 2499
rect 11989 2465 12023 2499
rect 12633 2465 12667 2499
rect 28181 2465 28215 2499
rect 28365 2329 28399 2363
rect 11667 2261 11701 2295
rect 12817 2261 12851 2295
<< metal1 >>
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 19150 15620 19156 15632
rect 11204 15592 19156 15620
rect 11204 15580 11210 15592
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 16206 15552 16212 15564
rect 15528 15524 16212 15552
rect 15528 15512 15534 15524
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28718 15552 28724 15564
rect 28040 15524 28724 15552
rect 28040 15512 28046 15524
rect 28718 15512 28724 15524
rect 28776 15512 28782 15564
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 21212 13379 21270 13385
rect 21212 13376 21224 13379
rect 20864 13348 21224 13376
rect 20864 13336 20870 13348
rect 21212 13345 21224 13348
rect 21258 13345 21270 13379
rect 21212 13339 21270 13345
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11882 13308 11888 13320
rect 11563 13280 11888 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20438 13308 20444 13320
rect 20119 13280 20444 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 106 13132 112 13184
rect 164 13172 170 13184
rect 12342 13172 12348 13184
rect 164 13144 12348 13172
rect 164 13132 170 13144
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 16117 13175 16175 13181
rect 16117 13172 16129 13175
rect 15896 13144 16129 13172
rect 15896 13132 15902 13144
rect 16117 13141 16129 13144
rect 16163 13141 16175 13175
rect 16117 13135 16175 13141
rect 20070 13132 20076 13184
rect 20128 13172 20134 13184
rect 21315 13175 21373 13181
rect 21315 13172 21327 13175
rect 20128 13144 21327 13172
rect 20128 13132 20134 13144
rect 21315 13141 21327 13144
rect 21361 13141 21373 13175
rect 21315 13135 21373 13141
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 7055 12971 7113 12977
rect 7055 12937 7067 12971
rect 7101 12968 7113 12971
rect 7190 12968 7196 12980
rect 7101 12940 7196 12968
rect 7101 12937 7113 12940
rect 7055 12931 7113 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 10919 12971 10977 12977
rect 10919 12937 10931 12971
rect 10965 12968 10977 12971
rect 13354 12968 13360 12980
rect 10965 12940 13360 12968
rect 10965 12937 10977 12940
rect 10919 12931 10977 12937
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 22097 12971 22155 12977
rect 22097 12937 22109 12971
rect 22143 12968 22155 12971
rect 23750 12968 23756 12980
rect 22143 12940 23756 12968
rect 22143 12937 22155 12940
rect 22097 12931 22155 12937
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 25225 12971 25283 12977
rect 25225 12937 25237 12971
rect 25271 12968 25283 12971
rect 25774 12968 25780 12980
rect 25271 12940 25780 12968
rect 25271 12937 25283 12940
rect 25225 12931 25283 12937
rect 25774 12928 25780 12940
rect 25832 12928 25838 12980
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 29457 12903 29515 12909
rect 29457 12869 29469 12903
rect 29503 12900 29515 12903
rect 35894 12900 35900 12912
rect 29503 12872 35900 12900
rect 29503 12869 29515 12872
rect 29457 12863 29515 12869
rect 35894 12860 35900 12872
rect 35952 12860 35958 12912
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 13262 12832 13268 12844
rect 7515 12804 13268 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 2593 12767 2651 12773
rect 2593 12733 2605 12767
rect 2639 12764 2651 12767
rect 2774 12764 2780 12776
rect 2639 12736 2780 12764
rect 2639 12733 2651 12736
rect 2593 12727 2651 12733
rect 2774 12724 2780 12736
rect 2832 12764 2838 12776
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 2832 12736 3065 12764
rect 2832 12724 2838 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 6984 12767 7042 12773
rect 6984 12733 6996 12767
rect 7030 12764 7042 12767
rect 7484 12764 7512 12795
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 24486 12832 24492 12844
rect 19996 12804 24492 12832
rect 7030 12736 7512 12764
rect 8757 12767 8815 12773
rect 7030 12733 7042 12736
rect 6984 12727 7042 12733
rect 8757 12733 8769 12767
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12628 2835 12631
rect 3142 12628 3148 12640
rect 2823 12600 3148 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 8662 12628 8668 12640
rect 8619 12600 8668 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 8662 12588 8668 12600
rect 8720 12628 8726 12640
rect 8772 12628 8800 12727
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10848 12767 10906 12773
rect 10848 12764 10860 12767
rect 10468 12736 10860 12764
rect 10468 12724 10474 12736
rect 10848 12733 10860 12736
rect 10894 12764 10906 12767
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 10894 12736 11253 12764
rect 10894 12733 10906 12736
rect 10848 12727 10906 12733
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 19996 12773 20024 12804
rect 24486 12792 24492 12804
rect 24544 12792 24550 12844
rect 25685 12835 25743 12841
rect 25685 12801 25697 12835
rect 25731 12832 25743 12835
rect 32766 12832 32772 12844
rect 25731 12804 32772 12832
rect 25731 12801 25743 12804
rect 25685 12795 25743 12801
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 13412 12736 14933 12764
rect 13412 12724 13418 12736
rect 14921 12733 14933 12736
rect 14967 12764 14979 12767
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 14967 12736 15393 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15381 12733 15393 12736
rect 15427 12733 15439 12767
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 15381 12727 15439 12733
rect 19812 12736 19993 12764
rect 15838 12656 15844 12708
rect 15896 12696 15902 12708
rect 16209 12699 16267 12705
rect 16209 12696 16221 12699
rect 15896 12668 16221 12696
rect 15896 12656 15902 12668
rect 16209 12665 16221 12668
rect 16255 12665 16267 12699
rect 16209 12659 16267 12665
rect 16301 12699 16359 12705
rect 16301 12665 16313 12699
rect 16347 12665 16359 12699
rect 16301 12659 16359 12665
rect 8938 12628 8944 12640
rect 8720 12600 8800 12628
rect 8899 12600 8944 12628
rect 8720 12588 8726 12600
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 15105 12631 15163 12637
rect 15105 12597 15117 12631
rect 15151 12628 15163 12631
rect 15746 12628 15752 12640
rect 15151 12600 15752 12628
rect 15151 12597 15163 12600
rect 15105 12591 15163 12597
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 16316 12628 16344 12659
rect 19812 12640 19840 12736
rect 19981 12733 19993 12736
rect 20027 12733 20039 12767
rect 20438 12764 20444 12776
rect 20399 12736 20444 12764
rect 19981 12727 20039 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 21450 12724 21456 12776
rect 21508 12764 21514 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 21508 12736 21925 12764
rect 21508 12724 21514 12736
rect 21913 12733 21925 12736
rect 21959 12764 21971 12767
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 21959 12736 22477 12764
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22465 12733 22477 12736
rect 22511 12764 22523 12767
rect 22511 12736 23474 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 20714 12696 20720 12708
rect 20675 12668 20720 12696
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 23446 12696 23474 12736
rect 24394 12724 24400 12776
rect 24452 12764 24458 12776
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 24452 12736 25053 12764
rect 24452 12724 24458 12736
rect 25041 12733 25053 12736
rect 25087 12764 25099 12767
rect 25700 12764 25728 12795
rect 32766 12792 32772 12804
rect 32824 12792 32830 12844
rect 26180 12767 26238 12773
rect 26180 12764 26192 12767
rect 25087 12736 25728 12764
rect 25087 12733 25099 12736
rect 25041 12727 25099 12733
rect 26160 12733 26192 12764
rect 26226 12764 26238 12767
rect 26605 12767 26663 12773
rect 26605 12764 26617 12767
rect 26226 12736 26617 12764
rect 26226 12733 26238 12736
rect 26160 12727 26238 12733
rect 26605 12733 26617 12736
rect 26651 12764 26663 12767
rect 26651 12736 28994 12764
rect 26651 12733 26663 12736
rect 26605 12727 26663 12733
rect 26160 12696 26188 12727
rect 23446 12668 26188 12696
rect 28966 12696 28994 12736
rect 33870 12724 33876 12776
rect 33928 12764 33934 12776
rect 35437 12767 35495 12773
rect 35437 12764 35449 12767
rect 33928 12736 35449 12764
rect 33928 12724 33934 12736
rect 35437 12733 35449 12736
rect 35483 12764 35495 12767
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35483 12736 36001 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 31294 12696 31300 12708
rect 28966 12668 31300 12696
rect 31294 12656 31300 12668
rect 31352 12656 31358 12708
rect 18230 12628 18236 12640
rect 16071 12600 18236 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 19794 12628 19800 12640
rect 19755 12600 19800 12628
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 20864 12600 21189 12628
rect 20864 12588 20870 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 21177 12591 21235 12597
rect 26283 12631 26341 12637
rect 26283 12597 26295 12631
rect 26329 12628 26341 12631
rect 26418 12628 26424 12640
rect 26329 12600 26424 12628
rect 26329 12597 26341 12600
rect 26283 12591 26341 12597
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 29086 12628 29092 12640
rect 28999 12600 29092 12628
rect 29086 12588 29092 12600
rect 29144 12628 29150 12640
rect 29825 12631 29883 12637
rect 29825 12628 29837 12631
rect 29144 12600 29837 12628
rect 29144 12588 29150 12600
rect 29825 12597 29837 12600
rect 29871 12597 29883 12631
rect 29825 12591 29883 12597
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 18782 12424 18788 12436
rect 15620 12396 18788 12424
rect 15620 12384 15626 12396
rect 18782 12384 18788 12396
rect 18840 12424 18846 12436
rect 23290 12424 23296 12436
rect 18840 12396 23296 12424
rect 18840 12384 18846 12396
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 14 12316 20 12368
rect 72 12356 78 12368
rect 4203 12359 4261 12365
rect 4203 12356 4215 12359
rect 72 12328 4215 12356
rect 72 12316 78 12328
rect 4203 12325 4215 12328
rect 4249 12325 4261 12359
rect 16206 12356 16212 12368
rect 16167 12328 16212 12356
rect 4203 12319 4261 12325
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 21266 12316 21272 12368
rect 21324 12356 21330 12368
rect 26326 12356 26332 12368
rect 21324 12328 26332 12356
rect 21324 12316 21330 12328
rect 26326 12316 26332 12328
rect 26384 12356 26390 12368
rect 29086 12356 29092 12368
rect 26384 12328 29092 12356
rect 26384 12316 26390 12328
rect 29086 12316 29092 12328
rect 29144 12316 29150 12368
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2372 12260 2789 12288
rect 2372 12248 2378 12260
rect 2777 12257 2789 12260
rect 2823 12288 2835 12291
rect 3418 12288 3424 12300
rect 2823 12260 3424 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 4116 12291 4174 12297
rect 4116 12257 4128 12291
rect 4162 12288 4174 12291
rect 4982 12288 4988 12300
rect 4162 12260 4988 12288
rect 4162 12257 4174 12260
rect 4116 12251 4174 12257
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 6546 12288 6552 12300
rect 6507 12260 6552 12288
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 7596 12291 7654 12297
rect 7596 12288 7608 12291
rect 7524 12260 7608 12288
rect 7524 12248 7530 12260
rect 7596 12257 7608 12260
rect 7642 12257 7654 12291
rect 7596 12251 7654 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 10962 12288 10968 12300
rect 10923 12260 10968 12288
rect 10781 12251 10839 12257
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 10594 12112 10600 12164
rect 10652 12152 10658 12164
rect 10796 12152 10824 12251
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 12066 12288 12072 12300
rect 12027 12260 12072 12288
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 13078 12288 13084 12300
rect 13039 12260 13084 12288
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 19518 12248 19524 12300
rect 19576 12288 19582 12300
rect 19832 12291 19890 12297
rect 19832 12288 19844 12291
rect 19576 12260 19844 12288
rect 19576 12248 19582 12260
rect 19832 12257 19844 12260
rect 19878 12288 19890 12291
rect 21284 12288 21312 12316
rect 19878 12260 21312 12288
rect 22072 12291 22130 12297
rect 19878 12257 19890 12260
rect 19832 12251 19890 12257
rect 22072 12257 22084 12291
rect 22118 12288 22130 12291
rect 22278 12288 22284 12300
rect 22118 12260 22284 12288
rect 22118 12257 22130 12260
rect 22072 12251 22130 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 23014 12288 23020 12300
rect 22975 12260 23020 12288
rect 23014 12248 23020 12260
rect 23072 12248 23078 12300
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 26580 12291 26638 12297
rect 26580 12288 26592 12291
rect 25179 12260 26592 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 26580 12257 26592 12260
rect 26626 12288 26638 12291
rect 27430 12288 27436 12300
rect 26626 12260 27436 12288
rect 26626 12257 26638 12260
rect 26580 12251 26638 12257
rect 27430 12248 27436 12260
rect 27488 12248 27494 12300
rect 27985 12291 28043 12297
rect 27985 12257 27997 12291
rect 28031 12288 28043 12291
rect 28074 12288 28080 12300
rect 28031 12260 28080 12288
rect 28031 12257 28043 12260
rect 27985 12251 28043 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 33594 12248 33600 12300
rect 33652 12288 33658 12300
rect 33724 12291 33782 12297
rect 33724 12288 33736 12291
rect 33652 12260 33736 12288
rect 33652 12248 33658 12260
rect 33724 12257 33736 12260
rect 33770 12257 33782 12291
rect 33724 12251 33782 12257
rect 34768 12291 34826 12297
rect 34768 12257 34780 12291
rect 34814 12288 34826 12291
rect 35342 12288 35348 12300
rect 34814 12260 35348 12288
rect 34814 12257 34826 12260
rect 34768 12251 34826 12257
rect 35342 12248 35348 12260
rect 35400 12248 35406 12300
rect 11054 12220 11060 12232
rect 11015 12192 11060 12220
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12220 21051 12223
rect 21266 12220 21272 12232
rect 21039 12192 21272 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 16482 12152 16488 12164
rect 10652 12124 16488 12152
rect 10652 12112 10658 12124
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 16666 12152 16672 12164
rect 16627 12124 16672 12152
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 21910 12112 21916 12164
rect 21968 12152 21974 12164
rect 23155 12155 23213 12161
rect 23155 12152 23167 12155
rect 21968 12124 23167 12152
rect 21968 12112 21974 12124
rect 23155 12121 23167 12124
rect 23201 12121 23213 12155
rect 23155 12115 23213 12121
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2222 12084 2228 12096
rect 2087 12056 2228 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 3786 12084 3792 12096
rect 3747 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 6730 12084 6736 12096
rect 6691 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7699 12087 7757 12093
rect 7699 12053 7711 12087
rect 7745 12084 7757 12087
rect 8110 12084 8116 12096
rect 7745 12056 8116 12084
rect 7745 12053 7757 12056
rect 7699 12047 7757 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13446 12084 13452 12096
rect 13311 12056 13452 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13446 12044 13452 12056
rect 13504 12084 13510 12096
rect 19794 12084 19800 12096
rect 13504 12056 19800 12084
rect 13504 12044 13510 12056
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 19935 12087 19993 12093
rect 19935 12053 19947 12087
rect 19981 12084 19993 12087
rect 21726 12084 21732 12096
rect 19981 12056 21732 12084
rect 19981 12053 19993 12056
rect 19935 12047 19993 12053
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 22143 12087 22201 12093
rect 22143 12053 22155 12087
rect 22189 12084 22201 12087
rect 22922 12084 22928 12096
rect 22189 12056 22928 12084
rect 22189 12053 22201 12056
rect 22143 12047 22201 12053
rect 22922 12044 22928 12056
rect 22980 12044 22986 12096
rect 24670 12084 24676 12096
rect 24631 12056 24676 12084
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 25314 12084 25320 12096
rect 25275 12056 25320 12084
rect 25314 12044 25320 12056
rect 25372 12044 25378 12096
rect 26510 12044 26516 12096
rect 26568 12084 26574 12096
rect 26651 12087 26709 12093
rect 26651 12084 26663 12087
rect 26568 12056 26663 12084
rect 26568 12044 26574 12056
rect 26651 12053 26663 12056
rect 26697 12053 26709 12087
rect 26651 12047 26709 12053
rect 28169 12087 28227 12093
rect 28169 12053 28181 12087
rect 28215 12084 28227 12087
rect 28994 12084 29000 12096
rect 28215 12056 29000 12084
rect 28215 12053 28227 12056
rect 28169 12047 28227 12053
rect 28994 12044 29000 12056
rect 29052 12044 29058 12096
rect 33827 12087 33885 12093
rect 33827 12053 33839 12087
rect 33873 12084 33885 12087
rect 34698 12084 34704 12096
rect 33873 12056 34704 12084
rect 33873 12053 33885 12056
rect 33827 12047 33885 12053
rect 34698 12044 34704 12056
rect 34756 12044 34762 12096
rect 34839 12087 34897 12093
rect 34839 12053 34851 12087
rect 34885 12084 34897 12087
rect 36538 12084 36544 12096
rect 34885 12056 36544 12084
rect 34885 12053 34897 12056
rect 34839 12047 34897 12053
rect 36538 12044 36544 12056
rect 36596 12044 36602 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 10594 11880 10600 11892
rect 10555 11852 10600 11880
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 14231 11883 14289 11889
rect 14231 11849 14243 11883
rect 14277 11880 14289 11883
rect 15838 11880 15844 11892
rect 14277 11852 15844 11880
rect 14277 11849 14289 11852
rect 14231 11843 14289 11849
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16206 11880 16212 11892
rect 16071 11852 16212 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 21177 11883 21235 11889
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21266 11880 21272 11892
rect 21223 11852 21272 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 21266 11840 21272 11852
rect 21324 11880 21330 11892
rect 24486 11880 24492 11892
rect 21324 11852 21404 11880
rect 24447 11852 24492 11880
rect 21324 11840 21330 11852
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 2038 11812 2044 11824
rect 1719 11784 2044 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 2038 11772 2044 11784
rect 2096 11812 2102 11824
rect 2225 11815 2283 11821
rect 2225 11812 2237 11815
rect 2096 11784 2237 11812
rect 2096 11772 2102 11784
rect 2225 11781 2237 11784
rect 2271 11812 2283 11815
rect 2314 11812 2320 11824
rect 2271 11784 2320 11812
rect 2271 11781 2283 11784
rect 2225 11775 2283 11781
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 3694 11812 3700 11824
rect 2924 11784 3700 11812
rect 2924 11772 2930 11784
rect 3694 11772 3700 11784
rect 3752 11812 3758 11824
rect 3789 11815 3847 11821
rect 3789 11812 3801 11815
rect 3752 11784 3801 11812
rect 3752 11772 3758 11784
rect 3789 11781 3801 11784
rect 3835 11781 3847 11815
rect 12802 11812 12808 11824
rect 3789 11775 3847 11781
rect 11256 11784 12808 11812
rect 2774 11744 2780 11756
rect 2735 11716 2780 11744
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9214 11744 9220 11756
rect 8628 11716 9220 11744
rect 8628 11704 8634 11716
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 10410 11744 10416 11756
rect 9907 11716 10416 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 2130 11676 2136 11688
rect 2091 11648 2136 11676
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2372 11648 2421 11676
rect 2372 11636 2378 11648
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 2409 11639 2467 11645
rect 3160 11648 3709 11676
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3160 11549 3188 11648
rect 3697 11645 3709 11648
rect 3743 11676 3755 11679
rect 3786 11676 3792 11688
rect 3743 11648 3792 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4430 11676 4436 11688
rect 4019 11648 4436 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 2924 11512 3157 11540
rect 2924 11500 2930 11512
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3145 11503 3203 11509
rect 3510 11500 3516 11512
rect 3568 11540 3574 11552
rect 3988 11540 4016 11639
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 7650 11676 7656 11688
rect 7611 11648 7656 11676
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 10965 11679 11023 11685
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 6546 11608 6552 11620
rect 4672 11580 6552 11608
rect 4672 11568 4678 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 8294 11608 8300 11620
rect 8255 11580 8300 11608
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 9309 11611 9367 11617
rect 9309 11577 9321 11611
rect 9355 11577 9367 11611
rect 9309 11571 9367 11577
rect 3568 11512 4016 11540
rect 3568 11500 3574 11512
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 4120 11512 4169 11540
rect 4120 11500 4126 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 4982 11540 4988 11552
rect 4847 11512 4988 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5258 11540 5264 11552
rect 5219 11512 5264 11540
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 7466 11540 7472 11552
rect 5868 11512 7472 11540
rect 5868 11500 5874 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9324 11540 9352 11571
rect 10980 11552 11008 11639
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11256 11685 11284 11784
rect 12802 11772 12808 11784
rect 12860 11812 12866 11824
rect 13078 11812 13084 11824
rect 12860 11784 13084 11812
rect 12860 11772 12866 11784
rect 13078 11772 13084 11784
rect 13136 11812 13142 11824
rect 13449 11815 13507 11821
rect 13449 11812 13461 11815
rect 13136 11784 13461 11812
rect 13136 11772 13142 11784
rect 13449 11781 13461 11784
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 16666 11812 16672 11824
rect 13780 11784 16672 11812
rect 13780 11772 13786 11784
rect 16666 11772 16672 11784
rect 16724 11812 16730 11824
rect 16761 11815 16819 11821
rect 16761 11812 16773 11815
rect 16724 11784 16773 11812
rect 16724 11772 16730 11784
rect 16761 11781 16773 11784
rect 16807 11781 16819 11815
rect 16761 11775 16819 11781
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 12066 11744 12072 11756
rect 11931 11716 12072 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 15243 11747 15301 11753
rect 12124 11716 13216 11744
rect 12124 11704 12130 11716
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 11204 11648 11253 11676
rect 11204 11636 11210 11648
rect 11241 11645 11253 11648
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 13188 11620 13216 11716
rect 15243 11713 15255 11747
rect 15289 11744 15301 11747
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 15289 11716 16221 11744
rect 15289 11713 15301 11716
rect 15243 11707 15301 11713
rect 16209 11713 16221 11716
rect 16255 11744 16267 11747
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 16255 11716 17509 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 17497 11713 17509 11716
rect 17543 11713 17555 11747
rect 17497 11707 17555 11713
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 20438 11744 20444 11756
rect 19300 11716 20444 11744
rect 19300 11704 19306 11716
rect 14160 11679 14218 11685
rect 14160 11645 14172 11679
rect 14206 11676 14218 11679
rect 14206 11648 14688 11676
rect 14206 11645 14218 11648
rect 14160 11639 14218 11645
rect 11514 11608 11520 11620
rect 11475 11580 11520 11608
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12526 11608 12532 11620
rect 12487 11580 12532 11608
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13170 11608 13176 11620
rect 12676 11580 12721 11608
rect 13131 11580 13176 11608
rect 12676 11568 12682 11580
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 8996 11512 9352 11540
rect 10229 11543 10287 11549
rect 8996 11500 9002 11512
rect 10229 11509 10241 11543
rect 10275 11540 10287 11543
rect 10962 11540 10968 11552
rect 10275 11512 10968 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12636 11540 12664 11568
rect 14660 11549 14688 11648
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 15140 11679 15198 11685
rect 15140 11676 15152 11679
rect 14976 11648 15152 11676
rect 14976 11636 14982 11648
rect 15140 11645 15152 11648
rect 15186 11676 15198 11679
rect 15562 11676 15568 11688
rect 15186 11648 15568 11676
rect 15186 11645 15198 11648
rect 15140 11639 15198 11645
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 19518 11676 19524 11688
rect 17736 11648 19524 11676
rect 17736 11636 17742 11648
rect 19518 11636 19524 11648
rect 19576 11636 19582 11688
rect 20180 11685 20208 11716
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 21376 11753 21404 11852
rect 24486 11840 24492 11852
rect 24544 11880 24550 11892
rect 30098 11880 30104 11892
rect 24544 11852 30104 11880
rect 24544 11840 24550 11852
rect 30098 11840 30104 11852
rect 30156 11840 30162 11892
rect 31294 11880 31300 11892
rect 31255 11852 31300 11880
rect 31294 11840 31300 11852
rect 31352 11840 31358 11892
rect 33594 11880 33600 11892
rect 33555 11852 33600 11880
rect 33594 11840 33600 11852
rect 33652 11840 33658 11892
rect 35483 11883 35541 11889
rect 35483 11849 35495 11883
rect 35529 11880 35541 11883
rect 35710 11880 35716 11892
rect 35529 11852 35716 11880
rect 35529 11849 35541 11852
rect 35483 11843 35541 11849
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 25130 11772 25136 11824
rect 25188 11812 25194 11824
rect 27982 11812 27988 11824
rect 25188 11784 27988 11812
rect 25188 11772 25194 11784
rect 27982 11772 27988 11784
rect 28040 11772 28046 11824
rect 21361 11747 21419 11753
rect 21361 11713 21373 11747
rect 21407 11713 21419 11747
rect 24118 11744 24124 11756
rect 24079 11716 24124 11744
rect 21361 11707 21419 11713
rect 24118 11704 24124 11716
rect 24176 11744 24182 11756
rect 32122 11744 32128 11756
rect 24176 11716 32128 11744
rect 24176 11704 24182 11716
rect 32122 11704 32128 11716
rect 32180 11704 32186 11756
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11645 19855 11679
rect 19797 11639 19855 11645
rect 20165 11679 20223 11685
rect 20165 11645 20177 11679
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 23728 11679 23786 11685
rect 23728 11645 23740 11679
rect 23774 11676 23786 11679
rect 24136 11676 24164 11704
rect 23774 11648 24164 11676
rect 23774 11645 23786 11648
rect 23728 11639 23786 11645
rect 16298 11608 16304 11620
rect 16259 11580 16304 11608
rect 16298 11568 16304 11580
rect 16356 11568 16362 11620
rect 16482 11568 16488 11620
rect 16540 11608 16546 11620
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 16540 11580 18889 11608
rect 16540 11568 16546 11580
rect 18877 11577 18889 11580
rect 18923 11608 18935 11611
rect 18923 11580 19723 11608
rect 18923 11577 18935 11580
rect 18877 11571 18935 11577
rect 12299 11512 12664 11540
rect 14645 11543 14703 11549
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 15010 11540 15016 11552
rect 14691 11512 15016 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 17129 11543 17187 11549
rect 17129 11540 17141 11543
rect 16172 11512 17141 11540
rect 16172 11500 16178 11512
rect 17129 11509 17141 11512
rect 17175 11509 17187 11543
rect 19242 11540 19248 11552
rect 19203 11512 19248 11540
rect 17129 11503 17187 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 19695 11540 19723 11580
rect 19812 11552 19840 11639
rect 24486 11636 24492 11688
rect 24544 11676 24550 11688
rect 24673 11679 24731 11685
rect 24673 11676 24685 11679
rect 24544 11648 24685 11676
rect 24544 11636 24550 11648
rect 24673 11645 24685 11648
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 24762 11636 24768 11688
rect 24820 11676 24826 11688
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24820 11648 25145 11676
rect 24820 11636 24826 11648
rect 25133 11645 25145 11648
rect 25179 11676 25191 11679
rect 26050 11676 26056 11688
rect 25179 11648 26056 11676
rect 25179 11645 25191 11648
rect 25133 11639 25191 11645
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 26513 11679 26571 11685
rect 26513 11645 26525 11679
rect 26559 11645 26571 11679
rect 26694 11676 26700 11688
rect 26655 11648 26700 11676
rect 26513 11639 26571 11645
rect 20438 11608 20444 11620
rect 20399 11580 20444 11608
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 21453 11611 21511 11617
rect 21453 11577 21465 11611
rect 21499 11608 21511 11611
rect 21542 11608 21548 11620
rect 21499 11580 21548 11608
rect 21499 11577 21511 11580
rect 21453 11571 21511 11577
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 22002 11608 22008 11620
rect 21963 11580 22008 11608
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 22094 11568 22100 11620
rect 22152 11608 22158 11620
rect 23014 11608 23020 11620
rect 22152 11580 23020 11608
rect 22152 11568 22158 11580
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 25406 11608 25412 11620
rect 25367 11580 25412 11608
rect 25406 11568 25412 11580
rect 25464 11568 25470 11620
rect 25777 11611 25835 11617
rect 25777 11577 25789 11611
rect 25823 11608 25835 11611
rect 26528 11608 26556 11639
rect 26694 11636 26700 11648
rect 26752 11636 26758 11688
rect 30812 11679 30870 11685
rect 30812 11645 30824 11679
rect 30858 11676 30870 11679
rect 31294 11676 31300 11688
rect 30858 11648 31300 11676
rect 30858 11645 30870 11648
rect 30812 11639 30870 11645
rect 31294 11636 31300 11648
rect 31352 11636 31358 11688
rect 33848 11679 33906 11685
rect 33848 11645 33860 11679
rect 33894 11676 33906 11679
rect 33962 11676 33968 11688
rect 33894 11648 33968 11676
rect 33894 11645 33906 11648
rect 33848 11639 33906 11645
rect 33962 11636 33968 11648
rect 34020 11676 34026 11688
rect 34241 11679 34299 11685
rect 34241 11676 34253 11679
rect 34020 11648 34253 11676
rect 34020 11636 34026 11648
rect 34241 11645 34253 11648
rect 34287 11645 34299 11679
rect 34241 11639 34299 11645
rect 35158 11636 35164 11688
rect 35216 11676 35222 11688
rect 35380 11679 35438 11685
rect 35380 11676 35392 11679
rect 35216 11648 35392 11676
rect 35216 11636 35222 11648
rect 35380 11645 35392 11648
rect 35426 11676 35438 11679
rect 35805 11679 35863 11685
rect 35805 11676 35817 11679
rect 35426 11648 35817 11676
rect 35426 11645 35438 11648
rect 35380 11639 35438 11645
rect 35805 11645 35817 11648
rect 35851 11645 35863 11679
rect 35805 11639 35863 11645
rect 26602 11608 26608 11620
rect 25823 11580 26223 11608
rect 26528 11580 26608 11608
rect 25823 11577 25835 11580
rect 25777 11571 25835 11577
rect 19794 11540 19800 11552
rect 19695 11512 19800 11540
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 22278 11540 22284 11552
rect 22239 11512 22284 11540
rect 22278 11500 22284 11512
rect 22336 11500 22342 11552
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 23799 11543 23857 11549
rect 23799 11540 23811 11543
rect 23256 11512 23811 11540
rect 23256 11500 23262 11512
rect 23799 11509 23811 11512
rect 23845 11509 23857 11543
rect 26195 11540 26223 11580
rect 26602 11568 26608 11580
rect 26660 11568 26666 11620
rect 26970 11608 26976 11620
rect 26931 11580 26976 11608
rect 26970 11568 26976 11580
rect 27028 11568 27034 11620
rect 27341 11543 27399 11549
rect 27341 11540 27353 11543
rect 26195 11512 27353 11540
rect 23799 11503 23857 11509
rect 27341 11509 27353 11512
rect 27387 11540 27399 11543
rect 27430 11540 27436 11552
rect 27387 11512 27436 11540
rect 27387 11509 27399 11512
rect 27341 11503 27399 11509
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27522 11500 27528 11552
rect 27580 11540 27586 11552
rect 27801 11543 27859 11549
rect 27801 11540 27813 11543
rect 27580 11512 27813 11540
rect 27580 11500 27586 11512
rect 27801 11509 27813 11512
rect 27847 11509 27859 11543
rect 27801 11503 27859 11509
rect 28074 11500 28080 11552
rect 28132 11540 28138 11552
rect 28261 11543 28319 11549
rect 28261 11540 28273 11543
rect 28132 11512 28273 11540
rect 28132 11500 28138 11512
rect 28261 11509 28273 11512
rect 28307 11509 28319 11543
rect 28261 11503 28319 11509
rect 30883 11543 30941 11549
rect 30883 11509 30895 11543
rect 30929 11540 30941 11543
rect 31110 11540 31116 11552
rect 30929 11512 31116 11540
rect 30929 11509 30941 11512
rect 30883 11503 30941 11509
rect 31110 11500 31116 11512
rect 31168 11500 31174 11552
rect 31754 11540 31760 11552
rect 31715 11512 31760 11540
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 32766 11500 32772 11552
rect 32824 11540 32830 11552
rect 33594 11540 33600 11552
rect 32824 11512 33600 11540
rect 32824 11500 32830 11512
rect 33594 11500 33600 11512
rect 33652 11500 33658 11552
rect 33919 11543 33977 11549
rect 33919 11509 33931 11543
rect 33965 11540 33977 11543
rect 34146 11540 34152 11552
rect 33965 11512 34152 11540
rect 33965 11509 33977 11512
rect 33919 11503 33977 11509
rect 34146 11500 34152 11512
rect 34204 11500 34210 11552
rect 35161 11543 35219 11549
rect 35161 11509 35173 11543
rect 35207 11540 35219 11543
rect 35342 11540 35348 11552
rect 35207 11512 35348 11540
rect 35207 11509 35219 11512
rect 35161 11503 35219 11509
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 3694 11336 3700 11348
rect 3655 11308 3700 11336
rect 3694 11296 3700 11308
rect 3752 11336 3758 11348
rect 4246 11336 4252 11348
rect 3752 11308 4252 11336
rect 3752 11296 3758 11308
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 7650 11336 7656 11348
rect 7611 11308 7656 11336
rect 7650 11296 7656 11308
rect 7708 11336 7714 11348
rect 9214 11336 9220 11348
rect 7708 11308 8248 11336
rect 9175 11308 9220 11336
rect 7708 11296 7714 11308
rect 8110 11268 8116 11280
rect 8071 11240 8116 11268
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8220 11277 8248 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 18690 11336 18696 11348
rect 12584 11308 18696 11336
rect 12584 11296 12590 11308
rect 8205 11271 8263 11277
rect 8205 11237 8217 11271
rect 8251 11268 8263 11271
rect 8938 11268 8944 11280
rect 8251 11240 8944 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 11974 11268 11980 11280
rect 11935 11240 11980 11268
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 13538 11268 13544 11280
rect 13499 11240 13544 11268
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 17236 11277 17264 11308
rect 18690 11296 18696 11308
rect 18748 11336 18754 11348
rect 18748 11308 18828 11336
rect 18748 11296 18754 11308
rect 16669 11271 16727 11277
rect 16669 11268 16681 11271
rect 16264 11240 16681 11268
rect 16264 11228 16270 11240
rect 16669 11237 16681 11240
rect 16715 11237 16727 11271
rect 16669 11231 16727 11237
rect 17221 11271 17279 11277
rect 17221 11237 17233 11271
rect 17267 11237 17279 11271
rect 18230 11268 18236 11280
rect 18191 11240 18236 11268
rect 17221 11231 17279 11237
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18800 11277 18828 11308
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 19935 11339 19993 11345
rect 19935 11336 19947 11339
rect 19208 11308 19947 11336
rect 19208 11296 19214 11308
rect 19935 11305 19947 11308
rect 19981 11305 19993 11339
rect 19935 11299 19993 11305
rect 20530 11296 20536 11348
rect 20588 11336 20594 11348
rect 23707 11339 23765 11345
rect 20588 11308 22667 11336
rect 20588 11296 20594 11308
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11237 18843 11271
rect 18785 11231 18843 11237
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 21913 11271 21971 11277
rect 21913 11268 21925 11271
rect 21692 11240 21925 11268
rect 21692 11228 21698 11240
rect 21913 11237 21925 11240
rect 21959 11237 21971 11271
rect 21913 11231 21971 11237
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1820 11172 1961 11200
rect 1820 11160 1826 11172
rect 1949 11169 1961 11172
rect 1995 11169 2007 11203
rect 1949 11163 2007 11169
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 2222 11200 2228 11212
rect 2096 11172 2141 11200
rect 2183 11172 2228 11200
rect 2096 11160 2102 11172
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4430 11200 4436 11212
rect 4387 11172 4436 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15508 11203 15566 11209
rect 15508 11200 15520 11203
rect 15344 11172 15520 11200
rect 15344 11160 15350 11172
rect 15508 11169 15520 11172
rect 15554 11169 15566 11203
rect 16298 11200 16304 11212
rect 16259 11172 16304 11200
rect 15508 11163 15566 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 19864 11203 19922 11209
rect 19864 11169 19876 11203
rect 19910 11169 19922 11203
rect 22639 11200 22667 11308
rect 23707 11305 23719 11339
rect 23753 11336 23765 11339
rect 27982 11336 27988 11348
rect 23753 11308 27988 11336
rect 23753 11305 23765 11308
rect 23707 11299 23765 11305
rect 27982 11296 27988 11308
rect 28040 11296 28046 11348
rect 30374 11336 30380 11348
rect 30335 11308 30380 11336
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 32309 11339 32367 11345
rect 32309 11305 32321 11339
rect 32355 11336 32367 11339
rect 33318 11336 33324 11348
rect 32355 11308 33324 11336
rect 32355 11305 32367 11308
rect 32309 11299 32367 11305
rect 33318 11296 33324 11308
rect 33376 11296 33382 11348
rect 26234 11268 26240 11280
rect 26195 11240 26240 11268
rect 26234 11228 26240 11240
rect 26292 11228 26298 11280
rect 26418 11228 26424 11280
rect 26476 11268 26482 11280
rect 26605 11271 26663 11277
rect 26605 11268 26617 11271
rect 26476 11240 26617 11268
rect 26476 11228 26482 11240
rect 26605 11237 26617 11240
rect 26651 11237 26663 11271
rect 26605 11231 26663 11237
rect 26694 11228 26700 11280
rect 26752 11268 26758 11280
rect 28307 11271 28365 11277
rect 26752 11240 26797 11268
rect 26752 11228 26758 11240
rect 28307 11237 28319 11271
rect 28353 11268 28365 11271
rect 30834 11268 30840 11280
rect 28353 11240 30840 11268
rect 28353 11237 28365 11240
rect 28307 11231 28365 11237
rect 30834 11228 30840 11240
rect 30892 11228 30898 11280
rect 34146 11228 34152 11280
rect 34204 11268 34210 11280
rect 34425 11271 34483 11277
rect 34425 11268 34437 11271
rect 34204 11240 34437 11268
rect 34204 11228 34210 11240
rect 34425 11237 34437 11240
rect 34471 11237 34483 11271
rect 34425 11231 34483 11237
rect 34517 11271 34575 11277
rect 34517 11237 34529 11271
rect 34563 11268 34575 11271
rect 34606 11268 34612 11280
rect 34563 11240 34612 11268
rect 34563 11237 34575 11240
rect 34517 11231 34575 11237
rect 34606 11228 34612 11240
rect 34664 11228 34670 11280
rect 22639 11172 23152 11200
rect 19864 11163 19922 11169
rect 1394 11092 1400 11144
rect 1452 11132 1458 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 1452 11104 2421 11132
rect 1452 11092 1458 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 2556 11104 4537 11132
rect 2556 11092 2562 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 8478 11132 8484 11144
rect 7239 11104 8484 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 8803 11104 9781 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9769 11101 9781 11104
rect 9815 11132 9827 11135
rect 10134 11132 10140 11144
rect 9815 11104 10140 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13630 11132 13636 11144
rect 13495 11104 13636 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 15611 11135 15669 11141
rect 15611 11101 15623 11135
rect 15657 11132 15669 11135
rect 16574 11132 16580 11144
rect 15657 11104 16580 11132
rect 15657 11101 15669 11104
rect 15611 11095 15669 11101
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4246 11064 4252 11076
rect 4203 11036 4252 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 12437 11067 12495 11073
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 13170 11064 13176 11076
rect 12483 11036 13176 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 13170 11024 13176 11036
rect 13228 11064 13234 11076
rect 13740 11064 13768 11095
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 19058 11132 19064 11144
rect 18187 11104 19064 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 13228 11036 13768 11064
rect 13228 11024 13234 11036
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 19879 11064 19907 11163
rect 21818 11132 21824 11144
rect 21779 11104 21824 11132
rect 21818 11092 21824 11104
rect 21876 11092 21882 11144
rect 22002 11092 22008 11144
rect 22060 11132 22066 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22060 11104 22477 11132
rect 22060 11092 22066 11104
rect 22465 11101 22477 11104
rect 22511 11132 22523 11135
rect 23014 11132 23020 11144
rect 22511 11104 23020 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 22020 11064 22048 11092
rect 19576 11036 22048 11064
rect 19576 11024 19582 11036
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 2866 10956 2872 11008
rect 2924 10996 2930 11008
rect 2961 10999 3019 11005
rect 2961 10996 2973 10999
rect 2924 10968 2973 10996
rect 2924 10956 2930 10968
rect 2961 10965 2973 10968
rect 3007 10965 3019 10999
rect 2961 10959 3019 10965
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 5077 10999 5135 11005
rect 5077 10996 5089 10999
rect 4948 10968 5089 10996
rect 4948 10956 4954 10968
rect 5077 10965 5089 10968
rect 5123 10965 5135 10999
rect 5077 10959 5135 10965
rect 10873 10999 10931 11005
rect 10873 10965 10885 10999
rect 10919 10996 10931 10999
rect 10962 10996 10968 11008
rect 10919 10968 10968 10996
rect 10919 10965 10931 10968
rect 10873 10959 10931 10965
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11146 10996 11152 11008
rect 11107 10968 11152 10996
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 15933 10999 15991 11005
rect 15933 10996 15945 10999
rect 15896 10968 15945 10996
rect 15896 10956 15902 10968
rect 15933 10965 15945 10968
rect 15979 10965 15991 10999
rect 15933 10959 15991 10965
rect 21361 10999 21419 11005
rect 21361 10965 21373 10999
rect 21407 10996 21419 10999
rect 21542 10996 21548 11008
rect 21407 10968 21548 10996
rect 21407 10965 21419 10968
rect 21361 10959 21419 10965
rect 21542 10956 21548 10968
rect 21600 10956 21606 11008
rect 23124 10996 23152 11172
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 23636 11203 23694 11209
rect 23636 11200 23648 11203
rect 23348 11172 23648 11200
rect 23348 11160 23354 11172
rect 23636 11169 23648 11172
rect 23682 11200 23694 11203
rect 23934 11200 23940 11212
rect 23682 11172 23940 11200
rect 23682 11169 23694 11172
rect 23636 11163 23694 11169
rect 23934 11160 23940 11172
rect 23992 11160 23998 11212
rect 24762 11200 24768 11212
rect 24723 11172 24768 11200
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 25041 11203 25099 11209
rect 25041 11169 25053 11203
rect 25087 11169 25099 11203
rect 25041 11163 25099 11169
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11200 28135 11203
rect 28166 11200 28172 11212
rect 28123 11172 28172 11200
rect 28123 11169 28135 11172
rect 28077 11163 28135 11169
rect 25056 11132 25084 11163
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 30098 11200 30104 11212
rect 30059 11172 30104 11200
rect 30098 11160 30104 11172
rect 30156 11160 30162 11212
rect 30561 11203 30619 11209
rect 30561 11169 30573 11203
rect 30607 11169 30619 11203
rect 32122 11200 32128 11212
rect 32083 11172 32128 11200
rect 30561 11163 30619 11169
rect 24136 11104 25084 11132
rect 25317 11135 25375 11141
rect 24136 11073 24164 11104
rect 25317 11101 25329 11135
rect 25363 11132 25375 11135
rect 26602 11132 26608 11144
rect 25363 11104 26608 11132
rect 25363 11101 25375 11104
rect 25317 11095 25375 11101
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 26878 11132 26884 11144
rect 26839 11104 26884 11132
rect 26878 11092 26884 11104
rect 26936 11092 26942 11144
rect 28994 11092 29000 11144
rect 29052 11132 29058 11144
rect 30576 11132 30604 11163
rect 32122 11160 32128 11172
rect 32180 11200 32186 11212
rect 33356 11203 33414 11209
rect 33356 11200 33368 11203
rect 32180 11172 33368 11200
rect 32180 11160 32186 11172
rect 33356 11169 33368 11172
rect 33402 11169 33414 11203
rect 33356 11163 33414 11169
rect 35897 11203 35955 11209
rect 35897 11169 35909 11203
rect 35943 11200 35955 11203
rect 35986 11200 35992 11212
rect 35943 11172 35992 11200
rect 35943 11169 35955 11172
rect 35897 11163 35955 11169
rect 35986 11160 35992 11172
rect 36044 11160 36050 11212
rect 31018 11132 31024 11144
rect 29052 11104 31024 11132
rect 29052 11092 29058 11104
rect 31018 11092 31024 11104
rect 31076 11092 31082 11144
rect 24121 11067 24179 11073
rect 24121 11064 24133 11067
rect 23584 11036 24133 11064
rect 23584 11008 23612 11036
rect 24121 11033 24133 11036
rect 24167 11033 24179 11067
rect 24121 11027 24179 11033
rect 26234 11024 26240 11076
rect 26292 11064 26298 11076
rect 31386 11064 31392 11076
rect 26292 11036 31392 11064
rect 26292 11024 26298 11036
rect 31386 11024 31392 11036
rect 31444 11024 31450 11076
rect 34974 11064 34980 11076
rect 34935 11036 34980 11064
rect 34974 11024 34980 11036
rect 35032 11064 35038 11076
rect 35713 11067 35771 11073
rect 35713 11064 35725 11067
rect 35032 11036 35725 11064
rect 35032 11024 35038 11036
rect 35713 11033 35725 11036
rect 35759 11033 35771 11067
rect 35713 11027 35771 11033
rect 23566 10996 23572 11008
rect 23124 10968 23572 10996
rect 23566 10956 23572 10968
rect 23624 10956 23630 11008
rect 25774 10996 25780 11008
rect 25735 10968 25780 10996
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 29822 10996 29828 11008
rect 29783 10968 29828 10996
rect 29822 10956 29828 10968
rect 29880 10956 29886 11008
rect 32950 10956 32956 11008
rect 33008 10996 33014 11008
rect 33459 10999 33517 11005
rect 33459 10996 33471 10999
rect 33008 10968 33471 10996
rect 33008 10956 33014 10968
rect 33459 10965 33471 10968
rect 33505 10965 33517 10999
rect 33459 10959 33517 10965
rect 35066 10956 35072 11008
rect 35124 10996 35130 11008
rect 35345 10999 35403 11005
rect 35345 10996 35357 10999
rect 35124 10968 35357 10996
rect 35124 10956 35130 10968
rect 35345 10965 35357 10968
rect 35391 10965 35403 10999
rect 35345 10959 35403 10965
rect 35802 10956 35808 11008
rect 35860 10996 35866 11008
rect 36035 10999 36093 11005
rect 36035 10996 36047 10999
rect 35860 10968 36047 10996
rect 35860 10956 35866 10968
rect 36035 10965 36047 10968
rect 36081 10965 36093 10999
rect 36035 10959 36093 10965
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2096 10764 2329 10792
rect 2096 10752 2102 10764
rect 2317 10761 2329 10764
rect 2363 10792 2375 10795
rect 4430 10792 4436 10804
rect 2363 10764 3004 10792
rect 4391 10764 4436 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2976 10736 3004 10764
rect 4430 10752 4436 10764
rect 4488 10752 4494 10804
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 6914 10792 6920 10804
rect 6595 10764 6920 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8352 10764 9321 10792
rect 8352 10752 8358 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 1578 10684 1584 10736
rect 1636 10724 1642 10736
rect 2685 10727 2743 10733
rect 2685 10724 2697 10727
rect 1636 10696 2697 10724
rect 1636 10684 1642 10696
rect 2685 10693 2697 10696
rect 2731 10693 2743 10727
rect 2958 10724 2964 10736
rect 2871 10696 2964 10724
rect 2685 10687 2743 10693
rect 2700 10656 2728 10687
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4982 10724 4988 10736
rect 4028 10696 4988 10724
rect 4028 10684 4034 10696
rect 4982 10684 4988 10696
rect 5040 10724 5046 10736
rect 5353 10727 5411 10733
rect 5353 10724 5365 10727
rect 5040 10696 5365 10724
rect 5040 10684 5046 10696
rect 5353 10693 5365 10696
rect 5399 10693 5411 10727
rect 5353 10687 5411 10693
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 7101 10727 7159 10733
rect 7101 10724 7113 10727
rect 6788 10696 7113 10724
rect 6788 10684 6794 10696
rect 7101 10693 7113 10696
rect 7147 10724 7159 10727
rect 8018 10724 8024 10736
rect 7147 10696 8024 10724
rect 7147 10693 7159 10696
rect 7101 10687 7159 10693
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 8938 10724 8944 10736
rect 8899 10696 8944 10724
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 3510 10656 3516 10668
rect 2700 10628 3516 10656
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1670 10588 1676 10600
rect 1443 10560 1676 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2866 10588 2872 10600
rect 2188 10560 2872 10588
rect 2188 10548 2194 10560
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3160 10597 3188 10628
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 4614 10656 4620 10668
rect 3651 10628 4620 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 4798 10656 4804 10668
rect 4711 10628 4804 10656
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 5258 10656 5264 10668
rect 4856 10628 5264 10656
rect 4856 10616 4862 10628
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10557 3203 10591
rect 7742 10588 7748 10600
rect 7703 10560 7748 10588
rect 3145 10551 3203 10557
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 4890 10480 4896 10532
rect 4948 10520 4954 10532
rect 7926 10520 7932 10532
rect 4948 10492 4993 10520
rect 7576 10492 7932 10520
rect 4948 10480 4954 10492
rect 106 10412 112 10464
rect 164 10452 170 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 164 10424 1593 10452
rect 164 10412 170 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1820 10424 1961 10452
rect 1820 10412 1826 10424
rect 1949 10421 1961 10424
rect 1995 10452 2007 10455
rect 4062 10452 4068 10464
rect 1995 10424 4068 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7576 10461 7604 10492
rect 7926 10480 7932 10492
rect 7984 10520 7990 10532
rect 8066 10523 8124 10529
rect 8066 10520 8078 10523
rect 7984 10492 8078 10520
rect 7984 10480 7990 10492
rect 8066 10489 8078 10492
rect 8112 10489 8124 10523
rect 9324 10520 9352 10755
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 9916 10764 10517 10792
rect 9916 10752 9922 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13538 10792 13544 10804
rect 13403 10764 13544 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13538 10752 13544 10764
rect 13596 10792 13602 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 13596 10764 13645 10792
rect 13596 10752 13602 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 14507 10795 14565 10801
rect 14507 10761 14519 10795
rect 14553 10792 14565 10795
rect 16114 10792 16120 10804
rect 14553 10764 16120 10792
rect 14553 10761 14565 10764
rect 14507 10755 14565 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16206 10752 16212 10804
rect 16264 10792 16270 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 16264 10764 16313 10792
rect 16264 10752 16270 10764
rect 16301 10761 16313 10764
rect 16347 10792 16359 10795
rect 16577 10795 16635 10801
rect 16577 10792 16589 10795
rect 16347 10764 16589 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16577 10761 16589 10764
rect 16623 10761 16635 10795
rect 16577 10755 16635 10761
rect 17865 10795 17923 10801
rect 17865 10761 17877 10795
rect 17911 10792 17923 10795
rect 18230 10792 18236 10804
rect 17911 10764 18236 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18230 10752 18236 10764
rect 18288 10752 18294 10804
rect 19058 10792 19064 10804
rect 19019 10764 19064 10792
rect 19058 10752 19064 10764
rect 19116 10792 19122 10804
rect 19751 10795 19809 10801
rect 19751 10792 19763 10795
rect 19116 10764 19763 10792
rect 19116 10752 19122 10764
rect 19751 10761 19763 10764
rect 19797 10761 19809 10795
rect 21542 10792 21548 10804
rect 21503 10764 21548 10792
rect 19751 10755 19809 10761
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 21818 10752 21824 10804
rect 21876 10792 21882 10804
rect 22189 10795 22247 10801
rect 22189 10792 22201 10795
rect 21876 10764 22201 10792
rect 21876 10752 21882 10764
rect 22189 10761 22201 10764
rect 22235 10792 22247 10795
rect 25222 10792 25228 10804
rect 22235 10764 25228 10792
rect 22235 10761 22247 10764
rect 22189 10755 22247 10761
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 26878 10752 26884 10804
rect 26936 10792 26942 10804
rect 31018 10792 31024 10804
rect 26936 10764 27470 10792
rect 30979 10764 31024 10792
rect 26936 10752 26942 10764
rect 10134 10724 10140 10736
rect 10095 10696 10140 10724
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 14001 10727 14059 10733
rect 14001 10724 14013 10727
rect 13780 10696 14013 10724
rect 13780 10684 13786 10696
rect 14001 10693 14013 10696
rect 14047 10693 14059 10727
rect 15286 10724 15292 10736
rect 15199 10696 15292 10724
rect 14001 10687 14059 10693
rect 15286 10684 15292 10696
rect 15344 10724 15350 10736
rect 18690 10724 18696 10736
rect 15344 10696 18552 10724
rect 18651 10696 18696 10724
rect 15344 10684 15350 10696
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 10594 10656 10600 10668
rect 9631 10628 10600 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 11572 10628 12449 10656
rect 11572 10616 11578 10628
rect 12437 10625 12449 10628
rect 12483 10656 12495 10659
rect 12526 10656 12532 10668
rect 12483 10628 12532 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14240 10628 15393 10656
rect 14240 10616 14246 10628
rect 15381 10625 15393 10628
rect 15427 10656 15439 10659
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 15427 10628 16957 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 18524 10656 18552 10696
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 19518 10724 19524 10736
rect 19479 10696 19524 10724
rect 19518 10684 19524 10696
rect 19576 10684 19582 10736
rect 22695 10727 22753 10733
rect 19771 10696 22416 10724
rect 19771 10656 19799 10696
rect 18524 10628 19799 10656
rect 16945 10619 17003 10625
rect 20438 10616 20444 10668
rect 20496 10656 20502 10668
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 20496 10628 20637 10656
rect 20496 10616 20502 10628
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 22388 10600 22416 10696
rect 22695 10693 22707 10727
rect 22741 10724 22753 10727
rect 22741 10696 27384 10724
rect 22741 10693 22753 10696
rect 22695 10687 22753 10693
rect 27356 10668 27384 10696
rect 23566 10616 23572 10668
rect 23624 10656 23630 10668
rect 23624 10628 24624 10656
rect 23624 10616 23630 10628
rect 24596 10600 24624 10628
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 26053 10659 26111 10665
rect 26053 10656 26065 10659
rect 25280 10628 26065 10656
rect 25280 10616 25286 10628
rect 26053 10625 26065 10628
rect 26099 10625 26111 10659
rect 27338 10656 27344 10668
rect 27251 10628 27344 10656
rect 26053 10619 26111 10625
rect 27338 10616 27344 10628
rect 27396 10616 27402 10668
rect 27442 10656 27470 10764
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 32858 10792 32864 10804
rect 31168 10764 32864 10792
rect 31168 10752 31174 10764
rect 32858 10752 32864 10764
rect 32916 10792 32922 10804
rect 32953 10795 33011 10801
rect 32953 10792 32965 10795
rect 32916 10764 32965 10792
rect 32916 10752 32922 10764
rect 32953 10761 32965 10764
rect 32999 10761 33011 10795
rect 32953 10755 33011 10761
rect 33962 10752 33968 10804
rect 34020 10792 34026 10804
rect 36909 10795 36967 10801
rect 36909 10792 36921 10795
rect 34020 10764 36921 10792
rect 34020 10752 34026 10764
rect 32122 10684 32128 10736
rect 32180 10724 32186 10736
rect 32585 10727 32643 10733
rect 32585 10724 32597 10727
rect 32180 10696 32597 10724
rect 32180 10684 32186 10696
rect 32585 10693 32597 10696
rect 32631 10724 32643 10727
rect 33502 10724 33508 10736
rect 32631 10696 33508 10724
rect 32631 10693 32643 10696
rect 32585 10687 32643 10693
rect 33502 10684 33508 10696
rect 33560 10684 33566 10736
rect 35158 10724 35164 10736
rect 34854 10696 35164 10724
rect 27617 10659 27675 10665
rect 27617 10656 27629 10659
rect 27442 10628 27629 10656
rect 27617 10625 27629 10628
rect 27663 10656 27675 10659
rect 28442 10656 28448 10668
rect 27663 10628 28448 10656
rect 27663 10625 27675 10628
rect 27617 10619 27675 10625
rect 28442 10616 28448 10628
rect 28500 10616 28506 10668
rect 29822 10656 29828 10668
rect 29783 10628 29828 10656
rect 29822 10616 29828 10628
rect 29880 10616 29886 10668
rect 31481 10659 31539 10665
rect 31481 10625 31493 10659
rect 31527 10656 31539 10659
rect 31665 10659 31723 10665
rect 31665 10656 31677 10659
rect 31527 10628 31677 10656
rect 31527 10625 31539 10628
rect 31481 10619 31539 10625
rect 31665 10625 31677 10628
rect 31711 10656 31723 10659
rect 31754 10656 31760 10668
rect 31711 10628 31760 10656
rect 31711 10625 31723 10628
rect 31665 10619 31723 10625
rect 31754 10616 31760 10628
rect 31812 10616 31818 10668
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10656 32367 10659
rect 34854 10656 34882 10696
rect 35158 10684 35164 10696
rect 35216 10724 35222 10736
rect 35216 10696 35296 10724
rect 35216 10684 35222 10696
rect 34974 10656 34980 10668
rect 32355 10628 34882 10656
rect 34935 10628 34980 10656
rect 32355 10625 32367 10628
rect 32309 10619 32367 10625
rect 34974 10616 34980 10628
rect 35032 10616 35038 10668
rect 35268 10665 35296 10696
rect 35253 10659 35311 10665
rect 35253 10625 35265 10659
rect 35299 10625 35311 10659
rect 35253 10619 35311 10625
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 11124 10591 11182 10597
rect 11124 10588 11136 10591
rect 10284 10560 11136 10588
rect 10284 10548 10290 10560
rect 11124 10557 11136 10560
rect 11170 10588 11182 10591
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 11170 10560 11621 10588
rect 11170 10557 11182 10560
rect 11124 10551 11182 10557
rect 11609 10557 11621 10560
rect 11655 10588 11667 10591
rect 13630 10588 13636 10600
rect 11655 10560 13636 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 14436 10591 14494 10597
rect 14436 10557 14448 10591
rect 14482 10588 14494 10591
rect 14482 10560 14780 10588
rect 14482 10557 14494 10560
rect 14436 10551 14494 10557
rect 9677 10523 9735 10529
rect 9677 10520 9689 10523
rect 9324 10492 9689 10520
rect 8066 10483 8124 10489
rect 9677 10489 9689 10492
rect 9723 10489 9735 10523
rect 9677 10483 9735 10489
rect 10965 10523 11023 10529
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 11974 10520 11980 10532
rect 11011 10492 11980 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 11974 10480 11980 10492
rect 12032 10480 12038 10532
rect 12758 10523 12816 10529
rect 12758 10489 12770 10523
rect 12804 10489 12816 10523
rect 12758 10483 12816 10489
rect 7561 10455 7619 10461
rect 7561 10452 7573 10455
rect 7064 10424 7573 10452
rect 7064 10412 7070 10424
rect 7561 10421 7573 10424
rect 7607 10421 7619 10455
rect 8662 10452 8668 10464
rect 8575 10424 8668 10452
rect 7561 10415 7619 10421
rect 8662 10412 8668 10424
rect 8720 10452 8726 10464
rect 9858 10452 9864 10464
rect 8720 10424 9864 10452
rect 8720 10412 8726 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 11195 10455 11253 10461
rect 11195 10452 11207 10455
rect 10652 10424 11207 10452
rect 10652 10412 10658 10424
rect 11195 10421 11207 10424
rect 11241 10421 11253 10455
rect 11195 10415 11253 10421
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11388 10424 12173 10452
rect 11388 10412 11394 10424
rect 12161 10421 12173 10424
rect 12207 10452 12219 10455
rect 12773 10452 12801 10483
rect 14752 10464 14780 10560
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 16356 10560 17417 10588
rect 16356 10548 16362 10560
rect 17405 10557 17417 10560
rect 17451 10588 17463 10591
rect 19680 10591 19738 10597
rect 17451 10560 18000 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 15743 10523 15801 10529
rect 15743 10489 15755 10523
rect 15789 10520 15801 10523
rect 15838 10520 15844 10532
rect 15789 10492 15844 10520
rect 15789 10489 15801 10492
rect 15743 10483 15801 10489
rect 15838 10480 15844 10492
rect 15896 10480 15902 10532
rect 12207 10424 12801 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14792 10424 14841 10452
rect 14792 10412 14798 10424
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 17972 10452 18000 10560
rect 19680 10557 19692 10591
rect 19726 10588 19738 10591
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 19726 10560 20085 10588
rect 19726 10557 19738 10560
rect 19680 10551 19738 10557
rect 20073 10557 20085 10560
rect 20119 10588 20131 10591
rect 21450 10588 21456 10600
rect 20119 10560 21456 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22592 10591 22650 10597
rect 22592 10588 22604 10591
rect 22428 10560 22604 10588
rect 22428 10548 22434 10560
rect 22592 10557 22604 10560
rect 22638 10588 22650 10591
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22638 10560 23029 10588
rect 22638 10557 22650 10560
rect 22592 10551 22650 10557
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23934 10588 23940 10600
rect 23895 10560 23940 10588
rect 23017 10551 23075 10557
rect 23934 10548 23940 10560
rect 23992 10548 23998 10600
rect 24118 10588 24124 10600
rect 24079 10560 24124 10588
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24578 10588 24584 10600
rect 24491 10560 24584 10588
rect 24578 10548 24584 10560
rect 24636 10548 24642 10600
rect 30745 10591 30803 10597
rect 30745 10557 30757 10591
rect 30791 10588 30803 10591
rect 30791 10560 31385 10588
rect 30791 10557 30803 10560
rect 30745 10551 30803 10557
rect 18138 10520 18144 10532
rect 18099 10492 18144 10520
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10489 18291 10523
rect 18233 10483 18291 10489
rect 20533 10523 20591 10529
rect 20533 10489 20545 10523
rect 20579 10520 20591 10523
rect 20987 10523 21045 10529
rect 20987 10520 20999 10523
rect 20579 10492 20999 10520
rect 20579 10489 20591 10492
rect 20533 10483 20591 10489
rect 20987 10489 20999 10492
rect 21033 10520 21045 10523
rect 21266 10520 21272 10532
rect 21033 10492 21272 10520
rect 21033 10489 21045 10492
rect 20987 10483 21045 10489
rect 18248 10452 18276 10483
rect 21266 10480 21272 10492
rect 21324 10480 21330 10532
rect 24854 10520 24860 10532
rect 24815 10492 24860 10520
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 24946 10480 24952 10532
rect 25004 10520 25010 10532
rect 25774 10520 25780 10532
rect 25004 10492 25780 10520
rect 25004 10480 25010 10492
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 25869 10523 25927 10529
rect 25869 10489 25881 10523
rect 25915 10520 25927 10523
rect 27065 10523 27123 10529
rect 27065 10520 27077 10523
rect 25915 10492 27077 10520
rect 25915 10489 25927 10492
rect 25869 10483 25927 10489
rect 27065 10489 27077 10492
rect 27111 10489 27123 10523
rect 27065 10483 27123 10489
rect 27433 10523 27491 10529
rect 27433 10489 27445 10523
rect 27479 10489 27491 10523
rect 27433 10483 27491 10489
rect 30146 10523 30204 10529
rect 30146 10489 30158 10523
rect 30192 10489 30204 10523
rect 31357 10520 31385 10560
rect 32398 10548 32404 10600
rect 32456 10588 32462 10600
rect 36531 10597 36559 10764
rect 36909 10761 36921 10764
rect 36955 10792 36967 10795
rect 39574 10792 39580 10804
rect 36955 10764 39580 10792
rect 36955 10761 36967 10764
rect 36909 10755 36967 10761
rect 39574 10752 39580 10764
rect 39632 10752 39638 10804
rect 37918 10656 37924 10668
rect 37879 10628 37924 10656
rect 37918 10616 37924 10628
rect 37976 10616 37982 10668
rect 33204 10591 33262 10597
rect 33204 10588 33216 10591
rect 32456 10560 33216 10588
rect 32456 10548 32462 10560
rect 33204 10557 33216 10560
rect 33250 10588 33262 10591
rect 33965 10591 34023 10597
rect 33965 10588 33977 10591
rect 33250 10560 33977 10588
rect 33250 10557 33262 10560
rect 33204 10551 33262 10557
rect 33965 10557 33977 10560
rect 34011 10557 34023 10591
rect 33965 10551 34023 10557
rect 36516 10591 36574 10597
rect 36516 10557 36528 10591
rect 36562 10557 36574 10591
rect 36516 10551 36574 10557
rect 37512 10591 37570 10597
rect 37512 10557 37524 10591
rect 37558 10588 37570 10591
rect 37936 10588 37964 10616
rect 37558 10560 37964 10588
rect 37558 10557 37570 10560
rect 37512 10551 37570 10557
rect 31662 10520 31668 10532
rect 31357 10492 31668 10520
rect 30146 10483 30204 10489
rect 17972 10424 18276 10452
rect 14829 10415 14887 10421
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 21692 10424 21833 10452
rect 21692 10412 21698 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 25225 10455 25283 10461
rect 25225 10452 25237 10455
rect 24820 10424 25237 10452
rect 24820 10412 24826 10424
rect 25225 10421 25237 10424
rect 25271 10452 25283 10455
rect 25314 10452 25320 10464
rect 25271 10424 25320 10452
rect 25271 10421 25283 10424
rect 25225 10415 25283 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 25590 10412 25596 10424
rect 25648 10452 25654 10464
rect 25884 10452 25912 10483
rect 26694 10452 26700 10464
rect 25648 10424 25912 10452
rect 26655 10424 26700 10452
rect 25648 10412 25654 10424
rect 26694 10412 26700 10424
rect 26752 10412 26758 10464
rect 27080 10452 27108 10483
rect 27448 10452 27476 10483
rect 27080 10424 27476 10452
rect 28166 10412 28172 10464
rect 28224 10452 28230 10464
rect 28261 10455 28319 10461
rect 28261 10452 28273 10455
rect 28224 10424 28273 10452
rect 28224 10412 28230 10424
rect 28261 10421 28273 10424
rect 28307 10421 28319 10455
rect 28261 10415 28319 10421
rect 29733 10455 29791 10461
rect 29733 10421 29745 10455
rect 29779 10452 29791 10455
rect 30161 10452 30189 10483
rect 31662 10480 31668 10492
rect 31720 10520 31726 10532
rect 31757 10523 31815 10529
rect 31757 10520 31769 10523
rect 31720 10492 31769 10520
rect 31720 10480 31726 10492
rect 31757 10489 31769 10492
rect 31803 10489 31815 10523
rect 31757 10483 31815 10489
rect 32490 10480 32496 10532
rect 32548 10520 32554 10532
rect 33410 10520 33416 10532
rect 32548 10492 33416 10520
rect 32548 10480 32554 10492
rect 33410 10480 33416 10492
rect 33468 10520 33474 10532
rect 34333 10523 34391 10529
rect 34333 10520 34345 10523
rect 33468 10492 34345 10520
rect 33468 10480 33474 10492
rect 34333 10489 34345 10492
rect 34379 10520 34391 10523
rect 34606 10520 34612 10532
rect 34379 10492 34612 10520
rect 34379 10489 34391 10492
rect 34333 10483 34391 10489
rect 34606 10480 34612 10492
rect 34664 10480 34670 10532
rect 35066 10520 35072 10532
rect 35027 10492 35072 10520
rect 35066 10480 35072 10492
rect 35124 10480 35130 10532
rect 35986 10520 35992 10532
rect 35947 10492 35992 10520
rect 35986 10480 35992 10492
rect 36044 10480 36050 10532
rect 36078 10480 36084 10532
rect 36136 10520 36142 10532
rect 37599 10523 37657 10529
rect 37599 10520 37611 10523
rect 36136 10492 37611 10520
rect 36136 10480 36142 10492
rect 37599 10489 37611 10492
rect 37645 10489 37657 10523
rect 37599 10483 37657 10489
rect 30650 10452 30656 10464
rect 29779 10424 30656 10452
rect 29779 10421 29791 10424
rect 29733 10415 29791 10421
rect 30650 10412 30656 10424
rect 30708 10412 30714 10464
rect 33134 10412 33140 10464
rect 33192 10452 33198 10464
rect 33275 10455 33333 10461
rect 33275 10452 33287 10455
rect 33192 10424 33287 10452
rect 33192 10412 33198 10424
rect 33275 10421 33287 10424
rect 33321 10421 33333 10455
rect 33275 10415 33333 10421
rect 33502 10412 33508 10464
rect 33560 10452 33566 10464
rect 33597 10455 33655 10461
rect 33597 10452 33609 10455
rect 33560 10424 33609 10452
rect 33560 10412 33566 10424
rect 33597 10421 33609 10424
rect 33643 10421 33655 10455
rect 33597 10415 33655 10421
rect 35250 10412 35256 10464
rect 35308 10452 35314 10464
rect 36587 10455 36645 10461
rect 36587 10452 36599 10455
rect 35308 10424 36599 10452
rect 35308 10412 35314 10424
rect 36587 10421 36599 10424
rect 36633 10421 36645 10455
rect 36587 10415 36645 10421
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 2958 10248 2964 10260
rect 2919 10220 2964 10248
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4798 10248 4804 10260
rect 4759 10220 4804 10248
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 4948 10220 5825 10248
rect 4948 10208 4954 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 5813 10211 5871 10217
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7098 10248 7104 10260
rect 6963 10220 7104 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7098 10208 7104 10220
rect 7156 10248 7162 10260
rect 7742 10248 7748 10260
rect 7156 10220 7748 10248
rect 7156 10208 7162 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8168 10220 8769 10248
rect 8168 10208 8174 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 10134 10248 10140 10260
rect 9539 10220 10140 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10229 10251 10287 10257
rect 10229 10217 10241 10251
rect 10275 10248 10287 10251
rect 10594 10248 10600 10260
rect 10275 10220 10600 10248
rect 10275 10217 10287 10220
rect 10229 10211 10287 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11054 10248 11060 10260
rect 10919 10220 11060 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 2317 10183 2375 10189
rect 2317 10180 2329 10183
rect 2280 10152 2329 10180
rect 2280 10140 2286 10152
rect 2317 10149 2329 10152
rect 2363 10180 2375 10183
rect 3237 10183 3295 10189
rect 3237 10180 3249 10183
rect 2363 10152 3249 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 3237 10149 3249 10152
rect 3283 10149 3295 10183
rect 5214 10183 5272 10189
rect 5214 10180 5226 10183
rect 3237 10143 3295 10149
rect 4724 10152 5226 10180
rect 4724 10124 4752 10152
rect 5214 10149 5226 10152
rect 5260 10149 5272 10183
rect 5214 10143 5272 10149
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 4706 10072 4712 10124
rect 4764 10072 4770 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8938 10112 8944 10124
rect 8527 10084 8944 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 10980 10121 11008 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 11974 10248 11980 10260
rect 11931 10220 11980 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 12676 10220 13645 10248
rect 12676 10208 12682 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 15838 10248 15844 10260
rect 15799 10220 15844 10248
rect 13633 10211 13691 10217
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 16298 10208 16304 10260
rect 16356 10248 16362 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 16356 10220 16405 10248
rect 16356 10208 16362 10220
rect 16393 10217 16405 10220
rect 16439 10217 16451 10251
rect 16393 10211 16451 10217
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16632 10220 17049 10248
rect 16632 10208 16638 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17586 10248 17592 10260
rect 17547 10220 17592 10248
rect 17037 10211 17095 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18782 10248 18788 10260
rect 18196 10220 18788 10248
rect 18196 10208 18202 10220
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20496 10220 20637 10248
rect 20496 10208 20502 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 20625 10211 20683 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21821 10251 21879 10257
rect 21821 10217 21833 10251
rect 21867 10248 21879 10251
rect 24118 10248 24124 10260
rect 21867 10220 22876 10248
rect 24079 10220 24124 10248
rect 21867 10217 21879 10220
rect 21821 10211 21879 10217
rect 22848 10192 22876 10220
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 26329 10251 26387 10257
rect 26329 10217 26341 10251
rect 26375 10248 26387 10251
rect 26418 10248 26424 10260
rect 26375 10220 26424 10248
rect 26375 10217 26387 10220
rect 26329 10211 26387 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 26568 10220 26648 10248
rect 26568 10208 26574 10220
rect 12986 10180 12992 10192
rect 12947 10152 12992 10180
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 22830 10180 22836 10192
rect 22743 10152 22836 10180
rect 22830 10140 22836 10152
rect 22888 10140 22894 10192
rect 25038 10180 25044 10192
rect 24999 10152 25044 10180
rect 25038 10140 25044 10152
rect 25096 10140 25102 10192
rect 26620 10189 26648 10220
rect 27338 10208 27344 10260
rect 27396 10248 27402 10260
rect 27525 10251 27583 10257
rect 27525 10248 27537 10251
rect 27396 10220 27537 10248
rect 27396 10208 27402 10220
rect 27525 10217 27537 10220
rect 27571 10217 27583 10251
rect 30098 10248 30104 10260
rect 30059 10220 30104 10248
rect 27525 10211 27583 10217
rect 30098 10208 30104 10220
rect 30156 10208 30162 10260
rect 30650 10248 30656 10260
rect 30611 10220 30656 10248
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 31662 10248 31668 10260
rect 31623 10220 31668 10248
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 34146 10208 34152 10260
rect 34204 10248 34210 10260
rect 34241 10251 34299 10257
rect 34241 10248 34253 10251
rect 34204 10220 34253 10248
rect 34204 10208 34210 10220
rect 34241 10217 34253 10220
rect 34287 10217 34299 10251
rect 34241 10211 34299 10217
rect 34698 10208 34704 10260
rect 34756 10248 34762 10260
rect 35437 10251 35495 10257
rect 35437 10248 35449 10251
rect 34756 10220 35449 10248
rect 34756 10208 34762 10220
rect 35437 10217 35449 10220
rect 35483 10217 35495 10251
rect 35437 10211 35495 10217
rect 25961 10183 26019 10189
rect 25961 10149 25973 10183
rect 26007 10180 26019 10183
rect 26605 10183 26663 10189
rect 26605 10180 26617 10183
rect 26007 10152 26617 10180
rect 26007 10149 26019 10152
rect 25961 10143 26019 10149
rect 26605 10149 26617 10152
rect 26651 10149 26663 10183
rect 26605 10143 26663 10149
rect 26694 10140 26700 10192
rect 26752 10180 26758 10192
rect 28258 10180 28264 10192
rect 26752 10152 26797 10180
rect 28219 10152 28264 10180
rect 26752 10140 26758 10152
rect 28258 10140 28264 10152
rect 28316 10140 28322 10192
rect 33054 10183 33112 10189
rect 33054 10149 33066 10183
rect 33100 10180 33112 10183
rect 33410 10180 33416 10192
rect 33100 10152 33416 10180
rect 33100 10149 33112 10152
rect 33054 10143 33112 10149
rect 33410 10140 33416 10152
rect 33468 10140 33474 10192
rect 34606 10180 34612 10192
rect 34567 10152 34612 10180
rect 34606 10140 34612 10152
rect 34664 10140 34670 10192
rect 35158 10180 35164 10192
rect 35119 10152 35164 10180
rect 35158 10140 35164 10152
rect 35216 10140 35222 10192
rect 35897 10183 35955 10189
rect 35897 10149 35909 10183
rect 35943 10180 35955 10183
rect 36078 10180 36084 10192
rect 35943 10152 36084 10180
rect 35943 10149 35955 10152
rect 35897 10143 35955 10149
rect 36078 10140 36084 10152
rect 36136 10140 36142 10192
rect 36170 10140 36176 10192
rect 36228 10180 36234 10192
rect 36228 10152 36273 10180
rect 36228 10140 36234 10152
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9088 10084 9689 10112
rect 9088 10072 9094 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11882 10072 11888 10124
rect 11940 10112 11946 10124
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 11940 10084 12173 10112
rect 11940 10072 11946 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 18230 10112 18236 10124
rect 18187 10084 18236 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19705 10115 19763 10121
rect 19705 10081 19717 10115
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 4890 10044 4896 10056
rect 4851 10016 4896 10044
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7524 10016 7573 10044
rect 7524 10004 7530 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 11572 10016 12725 10044
rect 11572 10004 11578 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 15252 10016 15485 10044
rect 15252 10004 15258 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 17218 10044 17224 10056
rect 17179 10016 17224 10044
rect 15473 10007 15531 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 19058 10004 19064 10056
rect 19116 10044 19122 10056
rect 19242 10044 19248 10056
rect 19116 10016 19248 10044
rect 19116 10004 19122 10016
rect 19242 10004 19248 10016
rect 19300 10044 19306 10056
rect 19720 10044 19748 10075
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20772 10084 20913 10112
rect 20772 10072 20778 10084
rect 20901 10081 20913 10084
rect 20947 10112 20959 10115
rect 21910 10112 21916 10124
rect 20947 10084 21916 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21910 10072 21916 10084
rect 21968 10072 21974 10124
rect 30285 10115 30343 10121
rect 30285 10081 30297 10115
rect 30331 10112 30343 10115
rect 30374 10112 30380 10124
rect 30331 10084 30380 10112
rect 30331 10081 30343 10084
rect 30285 10075 30343 10081
rect 30374 10072 30380 10084
rect 30432 10072 30438 10124
rect 19978 10044 19984 10056
rect 19300 10016 19748 10044
rect 19939 10016 19984 10044
rect 19300 10004 19306 10016
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 22738 10044 22744 10056
rect 22699 10016 22744 10044
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 23014 10044 23020 10056
rect 22975 10016 23020 10044
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10013 25007 10047
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 24949 10007 25007 10013
rect 24762 9936 24768 9988
rect 24820 9976 24826 9988
rect 24964 9976 24992 10007
rect 25222 10004 25228 10016
rect 25280 10044 25286 10056
rect 26881 10047 26939 10053
rect 26881 10044 26893 10047
rect 25280 10016 26893 10044
rect 25280 10004 25286 10016
rect 26881 10013 26893 10016
rect 26927 10013 26939 10047
rect 26881 10007 26939 10013
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28169 10047 28227 10053
rect 28169 10044 28181 10047
rect 28040 10016 28181 10044
rect 28040 10004 28046 10016
rect 28169 10013 28181 10016
rect 28215 10013 28227 10047
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 28169 10007 28227 10013
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 32950 10044 32956 10056
rect 32815 10016 32956 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 32950 10004 32956 10016
rect 33008 10004 33014 10056
rect 33597 10047 33655 10053
rect 33597 10013 33609 10047
rect 33643 10044 33655 10047
rect 33965 10047 34023 10053
rect 33965 10044 33977 10047
rect 33643 10016 33977 10044
rect 33643 10013 33655 10016
rect 33597 10007 33655 10013
rect 33965 10013 33977 10016
rect 34011 10044 34023 10047
rect 34517 10047 34575 10053
rect 34517 10044 34529 10047
rect 34011 10016 34529 10044
rect 34011 10013 34023 10016
rect 33965 10007 34023 10013
rect 34517 10013 34529 10016
rect 34563 10044 34575 10047
rect 34882 10044 34888 10056
rect 34563 10016 34888 10044
rect 34563 10013 34575 10016
rect 34517 10007 34575 10013
rect 34882 10004 34888 10016
rect 34940 10004 34946 10056
rect 34974 10004 34980 10056
rect 35032 10044 35038 10056
rect 36357 10047 36415 10053
rect 36357 10044 36369 10047
rect 35032 10016 36369 10044
rect 35032 10004 35038 10016
rect 36357 10013 36369 10016
rect 36403 10013 36415 10047
rect 36357 10007 36415 10013
rect 25866 9976 25872 9988
rect 24820 9948 25872 9976
rect 24820 9936 24826 9948
rect 25866 9936 25872 9948
rect 25924 9936 25930 9988
rect 7190 9908 7196 9920
rect 7151 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 9861 9911 9919 9917
rect 9861 9877 9873 9911
rect 9907 9908 9919 9911
rect 10962 9908 10968 9920
rect 9907 9880 10968 9908
rect 9907 9877 9919 9880
rect 9861 9871 9919 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 13780 9880 14381 9908
rect 13780 9868 13786 9880
rect 14369 9877 14381 9880
rect 14415 9877 14427 9911
rect 16666 9908 16672 9920
rect 16627 9880 16672 9908
rect 14369 9871 14427 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 24118 9908 24124 9920
rect 23440 9880 24124 9908
rect 23440 9868 23446 9880
rect 24118 9868 24124 9880
rect 24176 9868 24182 9920
rect 31202 9908 31208 9920
rect 31163 9880 31208 9908
rect 31202 9868 31208 9880
rect 31260 9868 31266 9920
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 2958 9704 2964 9716
rect 1964 9676 2964 9704
rect 1964 9645 1992 9676
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 9140 9676 9781 9704
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9605 2007 9639
rect 1949 9599 2007 9605
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 2188 9608 7639 9636
rect 2188 9596 2194 9608
rect 1670 9528 1676 9580
rect 1728 9568 1734 9580
rect 1728 9540 2176 9568
rect 1728 9528 1734 9540
rect 2148 9509 2176 9540
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 4948 9540 5549 9568
rect 4948 9528 4954 9540
rect 5537 9537 5549 9540
rect 5583 9568 5595 9571
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 5583 9540 5825 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5813 9537 5825 9540
rect 5859 9537 5871 9571
rect 7611 9568 7639 9608
rect 7611 9540 8064 9568
rect 5813 9531 5871 9537
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1780 9472 1869 9500
rect 1780 9376 1808 9472
rect 1857 9469 1869 9472
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9469 2191 9503
rect 2133 9463 2191 9469
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 2639 9472 3433 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 3421 9469 3433 9472
rect 3467 9500 3479 9503
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3467 9472 3893 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5166 9500 5172 9512
rect 5123 9472 5172 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 6914 9500 6920 9512
rect 5399 9472 6920 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 3510 9392 3516 9444
rect 3568 9432 3574 9444
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 3568 9404 4353 9432
rect 3568 9392 3574 9404
rect 4341 9401 4353 9404
rect 4387 9432 4399 9435
rect 5368 9432 5396 9463
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7190 9500 7196 9512
rect 7151 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 8036 9509 8064 9540
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 9140 9568 9168 9676
rect 9769 9673 9781 9676
rect 9815 9704 9827 9707
rect 10226 9704 10232 9716
rect 9815 9676 10232 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 12986 9704 12992 9716
rect 12636 9676 12992 9704
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9950 9636 9956 9648
rect 9355 9608 9956 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 8260 9540 9168 9568
rect 8260 9528 8266 9540
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8570 9500 8576 9512
rect 8067 9472 8576 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 4387 9404 5396 9432
rect 6641 9435 6699 9441
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 6641 9401 6653 9435
rect 6687 9432 6699 9435
rect 7374 9432 7380 9444
rect 6687 9404 7380 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7374 9392 7380 9404
rect 7432 9432 7438 9444
rect 7668 9432 7696 9463
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9140 9509 9168 9540
rect 11330 9528 11336 9580
rect 11388 9568 11394 9580
rect 12636 9577 12664 9676
rect 12986 9664 12992 9676
rect 13044 9704 13050 9716
rect 15381 9707 15439 9713
rect 15381 9704 15393 9707
rect 13044 9676 15393 9704
rect 13044 9664 13050 9676
rect 15381 9673 15393 9676
rect 15427 9704 15439 9707
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15427 9676 15761 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15749 9673 15761 9676
rect 15795 9704 15807 9707
rect 15838 9704 15844 9716
rect 15795 9676 15844 9704
rect 15795 9673 15807 9676
rect 15749 9667 15807 9673
rect 15838 9664 15844 9676
rect 15896 9704 15902 9716
rect 17221 9707 17279 9713
rect 17221 9704 17233 9707
rect 15896 9676 17233 9704
rect 15896 9664 15902 9676
rect 17221 9673 17233 9676
rect 17267 9704 17279 9707
rect 17586 9704 17592 9716
rect 17267 9676 17592 9704
rect 17267 9673 17279 9676
rect 17221 9667 17279 9673
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 18782 9664 18788 9716
rect 18840 9704 18846 9716
rect 19843 9707 19901 9713
rect 19843 9704 19855 9707
rect 18840 9676 19855 9704
rect 18840 9664 18846 9676
rect 19843 9673 19855 9676
rect 19889 9673 19901 9707
rect 21634 9704 21640 9716
rect 21595 9676 21640 9704
rect 19843 9667 19901 9673
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21910 9704 21916 9716
rect 21871 9676 21916 9704
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22465 9707 22523 9713
rect 22465 9673 22477 9707
rect 22511 9704 22523 9707
rect 22738 9704 22744 9716
rect 22511 9676 22744 9704
rect 22511 9673 22523 9676
rect 22465 9667 22523 9673
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 22830 9664 22836 9716
rect 22888 9704 22894 9716
rect 23385 9707 23443 9713
rect 23385 9704 23397 9707
rect 22888 9676 23397 9704
rect 22888 9664 22894 9676
rect 23385 9673 23397 9676
rect 23431 9673 23443 9707
rect 23385 9667 23443 9673
rect 23983 9707 24041 9713
rect 23983 9673 23995 9707
rect 24029 9704 24041 9707
rect 24946 9704 24952 9716
rect 24029 9676 24952 9704
rect 24029 9673 24041 9676
rect 23983 9667 24041 9673
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 25038 9664 25044 9716
rect 25096 9704 25102 9716
rect 25777 9707 25835 9713
rect 25777 9704 25789 9707
rect 25096 9676 25789 9704
rect 25096 9664 25102 9676
rect 25777 9673 25789 9676
rect 25823 9704 25835 9707
rect 26145 9707 26203 9713
rect 26145 9704 26157 9707
rect 25823 9676 26157 9704
rect 25823 9673 25835 9676
rect 25777 9667 25835 9673
rect 26145 9673 26157 9676
rect 26191 9704 26203 9707
rect 28169 9707 28227 9713
rect 28169 9704 28181 9707
rect 26191 9676 28181 9704
rect 26191 9673 26203 9676
rect 26145 9667 26203 9673
rect 28169 9673 28181 9676
rect 28215 9704 28227 9707
rect 28258 9704 28264 9716
rect 28215 9676 28264 9704
rect 28215 9673 28227 9676
rect 28169 9667 28227 9673
rect 28258 9664 28264 9676
rect 28316 9664 28322 9716
rect 28994 9704 29000 9716
rect 28955 9676 29000 9704
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 31202 9664 31208 9716
rect 31260 9704 31266 9716
rect 34333 9707 34391 9713
rect 34333 9704 34345 9707
rect 31260 9676 34345 9704
rect 31260 9664 31266 9676
rect 34333 9673 34345 9676
rect 34379 9704 34391 9707
rect 34606 9704 34612 9716
rect 34379 9676 34612 9704
rect 34379 9673 34391 9676
rect 34333 9667 34391 9673
rect 34606 9664 34612 9676
rect 34664 9664 34670 9716
rect 36081 9707 36139 9713
rect 36081 9673 36093 9707
rect 36127 9704 36139 9707
rect 36170 9704 36176 9716
rect 36127 9676 36176 9704
rect 36127 9673 36139 9676
rect 36081 9667 36139 9673
rect 36170 9664 36176 9676
rect 36228 9664 36234 9716
rect 13722 9636 13728 9648
rect 13188 9608 13728 9636
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 11388 9540 12633 9568
rect 11388 9528 11394 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 9125 9463 9183 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 10888 9432 10916 9463
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11020 9472 12265 9500
rect 11020 9460 11026 9472
rect 12253 9469 12265 9472
rect 12299 9500 12311 9503
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12299 9472 13093 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 13081 9469 13093 9472
rect 13127 9500 13139 9503
rect 13188 9500 13216 9608
rect 13722 9596 13728 9608
rect 13780 9636 13786 9648
rect 16853 9639 16911 9645
rect 13780 9608 14412 9636
rect 13780 9596 13786 9608
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 14182 9568 14188 9580
rect 13587 9540 14188 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 13354 9500 13360 9512
rect 13127 9472 13216 9500
rect 13267 9472 13360 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13354 9460 13360 9472
rect 13412 9500 13418 9512
rect 14384 9509 14412 9608
rect 16853 9605 16865 9639
rect 16899 9636 16911 9639
rect 18414 9636 18420 9648
rect 16899 9608 18420 9636
rect 16899 9605 16911 9608
rect 16853 9599 16911 9605
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 19334 9636 19340 9648
rect 19247 9608 19340 9636
rect 19334 9596 19340 9608
rect 19392 9636 19398 9648
rect 22756 9636 22784 9664
rect 23658 9636 23664 9648
rect 19392 9608 21588 9636
rect 22756 9608 23664 9636
rect 19392 9596 19398 9608
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 17218 9568 17224 9580
rect 15151 9540 17224 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 17218 9528 17224 9540
rect 17276 9568 17282 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 17276 9540 17601 9568
rect 17276 9528 17282 9540
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 18506 9568 18512 9580
rect 18467 9540 18512 9568
rect 17589 9531 17647 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20036 9540 20729 9568
rect 20036 9528 20042 9540
rect 20717 9537 20729 9540
rect 20763 9568 20775 9571
rect 21450 9568 21456 9580
rect 20763 9540 21456 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 21560 9568 21588 9608
rect 23658 9596 23664 9608
rect 23716 9596 23722 9648
rect 24394 9636 24400 9648
rect 24355 9608 24400 9636
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 26694 9596 26700 9648
rect 26752 9636 26758 9648
rect 27525 9639 27583 9645
rect 27525 9636 27537 9639
rect 26752 9608 27537 9636
rect 26752 9596 26758 9608
rect 27525 9605 27537 9608
rect 27571 9605 27583 9639
rect 27525 9599 27583 9605
rect 27982 9596 27988 9648
rect 28040 9636 28046 9648
rect 28445 9639 28503 9645
rect 28445 9636 28457 9639
rect 28040 9608 28457 9636
rect 28040 9596 28046 9608
rect 28445 9605 28457 9608
rect 28491 9605 28503 9639
rect 28445 9599 28503 9605
rect 24578 9568 24584 9580
rect 21560 9540 24584 9568
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 24854 9568 24860 9580
rect 24815 9540 24860 9568
rect 24854 9528 24860 9540
rect 24912 9528 24918 9580
rect 26602 9568 26608 9580
rect 26563 9540 26608 9568
rect 26602 9528 26608 9540
rect 26660 9528 26666 9580
rect 29012 9568 29040 9664
rect 31941 9639 31999 9645
rect 31941 9605 31953 9639
rect 31987 9636 31999 9639
rect 35066 9636 35072 9648
rect 31987 9608 35072 9636
rect 31987 9605 31999 9608
rect 31941 9599 31999 9605
rect 35066 9596 35072 9608
rect 35124 9596 35130 9648
rect 29822 9568 29828 9580
rect 29012 9540 29684 9568
rect 29783 9540 29828 9568
rect 14369 9503 14427 9509
rect 13412 9472 13814 9500
rect 13412 9460 13418 9472
rect 12158 9432 12164 9444
rect 7432 9404 7696 9432
rect 10244 9404 12164 9432
rect 7432 9392 7438 9404
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3605 9367 3663 9373
rect 3605 9364 3617 9367
rect 2648 9336 3617 9364
rect 2648 9324 2654 9336
rect 3605 9333 3617 9336
rect 3651 9333 3663 9367
rect 4706 9364 4712 9376
rect 4667 9336 4712 9364
rect 3605 9327 3663 9333
rect 4706 9324 4712 9336
rect 4764 9364 4770 9376
rect 7006 9364 7012 9376
rect 4764 9336 7012 9364
rect 4764 9324 4770 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 7156 9336 7297 9364
rect 7156 9324 7162 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 7285 9327 7343 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10244 9373 10272 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 9824 9336 10241 9364
rect 9824 9324 9830 9336
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 10229 9327 10287 9333
rect 10689 9367 10747 9373
rect 10689 9333 10701 9367
rect 10735 9364 10747 9367
rect 10870 9364 10876 9376
rect 10735 9336 10876 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11330 9364 11336 9376
rect 11020 9336 11336 9364
rect 11020 9324 11026 9336
rect 11330 9324 11336 9336
rect 11388 9364 11394 9376
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11388 9336 11437 9364
rect 11388 9324 11394 9336
rect 11425 9333 11437 9336
rect 11471 9333 11483 9367
rect 11425 9327 11483 9333
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11572 9336 11805 9364
rect 11572 9324 11578 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 13786 9364 13814 9472
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 14090 9392 14096 9444
rect 14148 9432 14154 9444
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 14148 9404 14289 9432
rect 14148 9392 14154 9404
rect 14277 9401 14289 9404
rect 14323 9432 14335 9435
rect 14844 9432 14872 9463
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15436 9472 15945 9500
rect 15436 9460 15442 9472
rect 15933 9469 15945 9472
rect 15979 9500 15991 9503
rect 16666 9500 16672 9512
rect 15979 9472 16672 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 19772 9503 19830 9509
rect 19772 9469 19784 9503
rect 19818 9500 19830 9503
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19818 9472 20269 9500
rect 19818 9469 19830 9472
rect 19772 9463 19830 9469
rect 20257 9469 20269 9472
rect 20303 9500 20315 9503
rect 22608 9503 22666 9509
rect 22608 9500 22620 9503
rect 20303 9472 22620 9500
rect 20303 9469 20315 9472
rect 20257 9463 20315 9469
rect 22608 9469 22620 9472
rect 22654 9500 22666 9503
rect 23912 9503 23970 9509
rect 22654 9469 22667 9500
rect 22608 9463 22667 9469
rect 23912 9469 23924 9503
rect 23958 9500 23970 9503
rect 24394 9500 24400 9512
rect 23958 9472 24400 9500
rect 23958 9469 23970 9472
rect 23912 9463 23970 9469
rect 14323 9404 14872 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 16022 9392 16028 9444
rect 16080 9432 16086 9444
rect 16254 9435 16312 9441
rect 16254 9432 16266 9435
rect 16080 9404 16266 9432
rect 16080 9392 16086 9404
rect 16254 9401 16266 9404
rect 16300 9401 16312 9435
rect 18138 9432 18144 9444
rect 18099 9404 18144 9432
rect 16254 9395 16312 9401
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9432 18291 9435
rect 18414 9432 18420 9444
rect 18279 9404 18420 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18414 9392 18420 9404
rect 18472 9392 18478 9444
rect 20625 9435 20683 9441
rect 20625 9401 20637 9435
rect 20671 9432 20683 9435
rect 21079 9435 21137 9441
rect 21079 9432 21091 9435
rect 20671 9404 21091 9432
rect 20671 9401 20683 9404
rect 20625 9395 20683 9401
rect 21079 9401 21091 9404
rect 21125 9432 21137 9435
rect 21266 9432 21272 9444
rect 21125 9404 21272 9432
rect 21125 9401 21137 9404
rect 21079 9395 21137 9401
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 13909 9367 13967 9373
rect 13909 9364 13921 9367
rect 13786 9336 13921 9364
rect 11793 9327 11851 9333
rect 13909 9333 13921 9336
rect 13955 9364 13967 9367
rect 13998 9364 14004 9376
rect 13955 9336 14004 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 19334 9364 19340 9376
rect 14700 9336 19340 9364
rect 14700 9324 14706 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 22639 9364 22667 9463
rect 24394 9460 24400 9472
rect 24452 9500 24458 9512
rect 27338 9500 27344 9512
rect 24452 9472 27344 9500
rect 24452 9460 24458 9472
rect 27338 9460 27344 9472
rect 27396 9460 27402 9512
rect 29270 9500 29276 9512
rect 29231 9472 29276 9500
rect 29270 9460 29276 9472
rect 29328 9460 29334 9512
rect 29656 9500 29684 9540
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 32858 9528 32864 9580
rect 32916 9568 32922 9580
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32916 9540 33057 9568
rect 32916 9528 32922 9540
rect 33045 9537 33057 9540
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 34974 9528 34980 9580
rect 35032 9568 35038 9580
rect 35253 9571 35311 9577
rect 35253 9568 35265 9571
rect 35032 9540 35265 9568
rect 35032 9528 35038 9540
rect 35253 9537 35265 9540
rect 35299 9537 35311 9571
rect 36538 9568 36544 9580
rect 36499 9540 36544 9568
rect 35253 9531 35311 9537
rect 36538 9528 36544 9540
rect 36596 9568 36602 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 36596 9540 37473 9568
rect 36596 9528 36602 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29656 9472 29745 9500
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 31021 9503 31079 9509
rect 31021 9469 31033 9503
rect 31067 9500 31079 9503
rect 31478 9500 31484 9512
rect 31067 9472 31484 9500
rect 31067 9469 31079 9472
rect 31021 9463 31079 9469
rect 31478 9460 31484 9472
rect 31536 9460 31542 9512
rect 22695 9435 22753 9441
rect 22695 9401 22707 9435
rect 22741 9432 22753 9435
rect 24762 9432 24768 9444
rect 22741 9404 24768 9432
rect 22741 9401 22753 9404
rect 22695 9395 22753 9401
rect 24762 9392 24768 9404
rect 24820 9392 24826 9444
rect 25178 9435 25236 9441
rect 25178 9432 25190 9435
rect 25056 9404 25190 9432
rect 25056 9376 25084 9404
rect 25178 9401 25190 9404
rect 25224 9401 25236 9435
rect 25178 9395 25236 9401
rect 26926 9435 26984 9441
rect 26926 9401 26938 9435
rect 26972 9401 26984 9435
rect 26926 9395 26984 9401
rect 30377 9435 30435 9441
rect 30377 9401 30389 9435
rect 30423 9432 30435 9435
rect 30650 9432 30656 9444
rect 30423 9404 30656 9432
rect 30423 9401 30435 9404
rect 30377 9395 30435 9401
rect 23106 9364 23112 9376
rect 22639 9336 23112 9364
rect 23106 9324 23112 9336
rect 23164 9324 23170 9376
rect 24673 9367 24731 9373
rect 24673 9333 24685 9367
rect 24719 9364 24731 9367
rect 25038 9364 25044 9376
rect 24719 9336 25044 9364
rect 24719 9333 24731 9336
rect 24673 9327 24731 9333
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 26510 9364 26516 9376
rect 26471 9336 26516 9364
rect 26510 9324 26516 9336
rect 26568 9364 26574 9376
rect 26941 9364 26969 9395
rect 30650 9392 30656 9404
rect 30708 9432 30714 9444
rect 30929 9435 30987 9441
rect 30929 9432 30941 9435
rect 30708 9404 30941 9432
rect 30708 9392 30714 9404
rect 30929 9401 30941 9404
rect 30975 9432 30987 9435
rect 31383 9435 31441 9441
rect 31383 9432 31395 9435
rect 30975 9404 31395 9432
rect 30975 9401 30987 9404
rect 30929 9395 30987 9401
rect 31383 9401 31395 9404
rect 31429 9432 31441 9435
rect 31570 9432 31576 9444
rect 31429 9404 31576 9432
rect 31429 9401 31441 9404
rect 31383 9395 31441 9401
rect 31570 9392 31576 9404
rect 31628 9392 31634 9444
rect 33137 9435 33195 9441
rect 32416 9404 32996 9432
rect 26568 9336 26969 9364
rect 26568 9324 26574 9336
rect 32306 9324 32312 9376
rect 32364 9364 32370 9376
rect 32416 9373 32444 9404
rect 32401 9367 32459 9373
rect 32401 9364 32413 9367
rect 32364 9336 32413 9364
rect 32364 9324 32370 9336
rect 32401 9333 32413 9336
rect 32447 9333 32459 9367
rect 32401 9327 32459 9333
rect 32490 9324 32496 9376
rect 32548 9364 32554 9376
rect 32769 9367 32827 9373
rect 32769 9364 32781 9367
rect 32548 9336 32781 9364
rect 32548 9324 32554 9336
rect 32769 9333 32781 9336
rect 32815 9333 32827 9367
rect 32968 9364 32996 9404
rect 33137 9401 33149 9435
rect 33183 9401 33195 9435
rect 33686 9432 33692 9444
rect 33647 9404 33692 9432
rect 33137 9395 33195 9401
rect 33152 9364 33180 9395
rect 33686 9392 33692 9404
rect 33744 9392 33750 9444
rect 34790 9392 34796 9444
rect 34848 9432 34854 9444
rect 34977 9435 35035 9441
rect 34977 9432 34989 9435
rect 34848 9404 34989 9432
rect 34848 9392 34854 9404
rect 34977 9401 34989 9404
rect 35023 9401 35035 9435
rect 34977 9395 35035 9401
rect 35069 9435 35127 9441
rect 35069 9401 35081 9435
rect 35115 9401 35127 9435
rect 35069 9395 35127 9401
rect 35728 9404 36124 9432
rect 34422 9364 34428 9376
rect 32968 9336 34428 9364
rect 32769 9327 32827 9333
rect 34422 9324 34428 9336
rect 34480 9324 34486 9376
rect 34514 9324 34520 9376
rect 34572 9364 34578 9376
rect 34701 9367 34759 9373
rect 34701 9364 34713 9367
rect 34572 9336 34713 9364
rect 34572 9324 34578 9336
rect 34701 9333 34713 9336
rect 34747 9364 34759 9367
rect 35084 9364 35112 9395
rect 35728 9364 35756 9404
rect 34747 9336 35756 9364
rect 36096 9364 36124 9404
rect 36630 9392 36636 9444
rect 36688 9432 36694 9444
rect 37182 9432 37188 9444
rect 36688 9404 36733 9432
rect 37143 9404 37188 9432
rect 36688 9392 36694 9404
rect 37182 9392 37188 9404
rect 37240 9392 37246 9444
rect 36648 9364 36676 9392
rect 36096 9336 36676 9364
rect 34747 9333 34759 9336
rect 34701 9327 34759 9333
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1728 9132 1869 9160
rect 1728 9120 1734 9132
rect 1857 9129 1869 9132
rect 1903 9160 1915 9163
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 1903 9132 2237 9160
rect 1903 9129 1915 9132
rect 1857 9123 1915 9129
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 7009 9163 7067 9169
rect 4028 9132 4844 9160
rect 4028 9120 4034 9132
rect 4816 9104 4844 9132
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 7055 9132 7205 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7193 9129 7205 9132
rect 7239 9160 7251 9163
rect 7466 9160 7472 9172
rect 7239 9132 7472 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8478 9160 8484 9172
rect 8439 9132 8484 9160
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10686 9160 10692 9172
rect 10551 9132 10692 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 13412 9132 14381 9160
rect 13412 9120 13418 9132
rect 14369 9129 14381 9132
rect 14415 9160 14427 9163
rect 14642 9160 14648 9172
rect 14415 9132 14648 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9160 16267 9163
rect 21450 9160 21456 9172
rect 16255 9132 17540 9160
rect 21411 9132 21456 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 17512 9104 17540 9132
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 23845 9163 23903 9169
rect 23845 9129 23857 9163
rect 23891 9160 23903 9163
rect 24210 9160 24216 9172
rect 23891 9132 24216 9160
rect 23891 9129 23903 9132
rect 23845 9123 23903 9129
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 24581 9163 24639 9169
rect 24581 9129 24593 9163
rect 24627 9160 24639 9163
rect 24854 9160 24860 9172
rect 24627 9132 24860 9160
rect 24627 9129 24639 9132
rect 24581 9123 24639 9129
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25038 9160 25044 9172
rect 24999 9132 25044 9160
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 25590 9160 25596 9172
rect 25551 9132 25596 9160
rect 25590 9120 25596 9132
rect 25648 9120 25654 9172
rect 25866 9160 25872 9172
rect 25827 9132 25872 9160
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 26329 9163 26387 9169
rect 26329 9129 26341 9163
rect 26375 9160 26387 9163
rect 26694 9160 26700 9172
rect 26375 9132 26700 9160
rect 26375 9129 26387 9132
rect 26329 9123 26387 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 26970 9120 26976 9172
rect 27028 9160 27034 9172
rect 27065 9163 27123 9169
rect 27065 9160 27077 9163
rect 27028 9132 27077 9160
rect 27028 9120 27034 9132
rect 27065 9129 27077 9132
rect 27111 9129 27123 9163
rect 29270 9160 29276 9172
rect 27065 9123 27123 9129
rect 27172 9132 29276 9160
rect 1946 9092 1952 9104
rect 1412 9064 1952 9092
rect 1412 9033 1440 9064
rect 1946 9052 1952 9064
rect 2004 9092 2010 9104
rect 3786 9092 3792 9104
rect 2004 9064 3792 9092
rect 2004 9052 2010 9064
rect 3786 9052 3792 9064
rect 3844 9052 3850 9104
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4249 9095 4307 9101
rect 4249 9092 4261 9095
rect 3936 9064 4261 9092
rect 3936 9052 3942 9064
rect 4249 9061 4261 9064
rect 4295 9061 4307 9095
rect 4798 9092 4804 9104
rect 4711 9064 4804 9092
rect 4249 9055 4307 9061
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11194 9095 11252 9101
rect 11194 9092 11206 9095
rect 11020 9064 11206 9092
rect 11020 9052 11026 9064
rect 11194 9061 11206 9064
rect 11240 9061 11252 9095
rect 12805 9095 12863 9101
rect 12805 9092 12817 9095
rect 11194 9055 11252 9061
rect 11808 9064 12817 9092
rect 11808 9036 11836 9064
rect 12805 9061 12817 9064
rect 12851 9061 12863 9095
rect 12805 9055 12863 9061
rect 15651 9095 15709 9101
rect 15651 9061 15663 9095
rect 15697 9092 15709 9095
rect 15930 9092 15936 9104
rect 15697 9064 15936 9092
rect 15697 9061 15709 9064
rect 15651 9055 15709 9061
rect 15930 9052 15936 9064
rect 15988 9052 15994 9104
rect 17494 9092 17500 9104
rect 17407 9064 17500 9092
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 19426 9092 19432 9104
rect 19387 9064 19432 9092
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 21910 9092 21916 9104
rect 21871 9064 21916 9092
rect 21910 9052 21916 9064
rect 21968 9052 21974 9104
rect 27172 9092 27200 9132
rect 29270 9120 29276 9132
rect 29328 9120 29334 9172
rect 30374 9120 30380 9172
rect 30432 9160 30438 9172
rect 31113 9163 31171 9169
rect 31113 9160 31125 9163
rect 30432 9132 31125 9160
rect 30432 9120 30438 9132
rect 31113 9129 31125 9132
rect 31159 9129 31171 9163
rect 34514 9160 34520 9172
rect 34475 9132 34520 9160
rect 31113 9123 31171 9129
rect 34514 9120 34520 9132
rect 34572 9120 34578 9172
rect 34974 9160 34980 9172
rect 34887 9132 34980 9160
rect 34974 9120 34980 9132
rect 35032 9160 35038 9172
rect 35802 9160 35808 9172
rect 35032 9132 35808 9160
rect 35032 9120 35038 9132
rect 35802 9120 35808 9132
rect 35860 9120 35866 9172
rect 36170 9120 36176 9172
rect 36228 9160 36234 9172
rect 36265 9163 36323 9169
rect 36265 9160 36277 9163
rect 36228 9132 36277 9160
rect 36228 9120 36234 9132
rect 36265 9129 36277 9132
rect 36311 9129 36323 9163
rect 36630 9160 36636 9172
rect 36591 9132 36636 9160
rect 36265 9123 36323 9129
rect 36630 9120 36636 9132
rect 36688 9120 36694 9172
rect 25792 9064 27200 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2372 8996 2421 9024
rect 2372 8984 2378 8996
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3510 9024 3516 9036
rect 3007 8996 3516 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 5718 9024 5724 9036
rect 5679 8996 5724 9024
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6178 9024 6184 9036
rect 5951 8996 6184 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7524 8996 7573 9024
rect 7524 8984 7530 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 11790 9024 11796 9036
rect 11703 8996 11796 9024
rect 7929 8987 7987 8993
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4212 8928 4257 8956
rect 4212 8916 4218 8928
rect 7282 8916 7288 8968
rect 7340 8956 7346 8968
rect 7944 8956 7972 8987
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 14182 9024 14188 9036
rect 14143 8996 14188 9024
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 23474 8984 23480 9036
rect 23532 9024 23538 9036
rect 23661 9027 23719 9033
rect 23661 9024 23673 9027
rect 23532 8996 23673 9024
rect 23532 8984 23538 8996
rect 23661 8993 23673 8996
rect 23707 9024 23719 9027
rect 25792 9024 25820 9064
rect 27522 9052 27528 9104
rect 27580 9092 27586 9104
rect 27801 9095 27859 9101
rect 27801 9092 27813 9095
rect 27580 9064 27813 9092
rect 27580 9052 27586 9064
rect 27801 9061 27813 9064
rect 27847 9061 27859 9095
rect 27801 9055 27859 9061
rect 27893 9095 27951 9101
rect 27893 9061 27905 9095
rect 27939 9092 27951 9095
rect 27982 9092 27988 9104
rect 27939 9064 27988 9092
rect 27939 9061 27951 9064
rect 27893 9055 27951 9061
rect 27982 9052 27988 9064
rect 28040 9052 28046 9104
rect 30279 9095 30337 9101
rect 30279 9061 30291 9095
rect 30325 9092 30337 9095
rect 30650 9092 30656 9104
rect 30325 9064 30656 9092
rect 30325 9061 30337 9064
rect 30279 9055 30337 9061
rect 30650 9052 30656 9064
rect 30708 9052 30714 9104
rect 33959 9095 34017 9101
rect 33959 9061 33971 9095
rect 34005 9092 34017 9095
rect 34606 9092 34612 9104
rect 34005 9064 34612 9092
rect 34005 9061 34017 9064
rect 33959 9055 34017 9061
rect 34606 9052 34612 9064
rect 34664 9092 34670 9104
rect 35707 9095 35765 9101
rect 35707 9092 35719 9095
rect 34664 9064 35719 9092
rect 34664 9052 34670 9064
rect 35707 9061 35719 9064
rect 35753 9092 35765 9095
rect 35894 9092 35900 9104
rect 35753 9064 35900 9092
rect 35753 9061 35765 9064
rect 35707 9055 35765 9061
rect 35894 9052 35900 9064
rect 35952 9052 35958 9104
rect 23707 8996 25820 9024
rect 23707 8993 23719 8996
rect 23661 8987 23719 8993
rect 26326 8984 26332 9036
rect 26384 9024 26390 9036
rect 26548 9027 26606 9033
rect 26548 9024 26560 9027
rect 26384 8996 26560 9024
rect 26384 8984 26390 8996
rect 26548 8993 26560 8996
rect 26594 8993 26606 9027
rect 26548 8987 26606 8993
rect 26694 8984 26700 9036
rect 26752 9024 26758 9036
rect 27433 9027 27491 9033
rect 27433 9024 27445 9027
rect 26752 8996 27445 9024
rect 26752 8984 26758 8996
rect 27433 8993 27445 8996
rect 27479 8993 27491 9027
rect 27433 8987 27491 8993
rect 30837 9027 30895 9033
rect 30837 8993 30849 9027
rect 30883 9024 30895 9027
rect 32490 9024 32496 9036
rect 30883 8996 32496 9024
rect 30883 8993 30895 8996
rect 30837 8987 30895 8993
rect 32490 8984 32496 8996
rect 32548 8984 32554 9036
rect 34422 8984 34428 9036
rect 34480 9024 34486 9036
rect 36630 9024 36636 9036
rect 34480 8996 36636 9024
rect 34480 8984 34486 8996
rect 36630 8984 36636 8996
rect 36688 9024 36694 9036
rect 36909 9027 36967 9033
rect 36909 9024 36921 9027
rect 36688 8996 36921 9024
rect 36688 8984 36694 8996
rect 36909 8993 36921 8996
rect 36955 8993 36967 9027
rect 36909 8987 36967 8993
rect 7340 8928 7972 8956
rect 9861 8959 9919 8965
rect 7340 8916 7346 8928
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10870 8956 10876 8968
rect 9907 8928 10272 8956
rect 10831 8928 10876 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 10244 8888 10272 8928
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 12713 8919 12771 8925
rect 12618 8888 12624 8900
rect 1627 8860 4108 8888
rect 10244 8860 12624 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 3970 8820 3976 8832
rect 3927 8792 3976 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4080 8820 4108 8860
rect 12618 8848 12624 8860
rect 12676 8888 12682 8900
rect 12728 8888 12756 8919
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8956 17463 8959
rect 17586 8956 17592 8968
rect 17451 8928 17592 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 17586 8916 17592 8928
rect 17644 8916 17650 8968
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8956 17739 8959
rect 18506 8956 18512 8968
rect 17727 8928 18512 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 13262 8888 13268 8900
rect 12676 8860 12756 8888
rect 13175 8860 13268 8888
rect 12676 8848 12682 8860
rect 13262 8848 13268 8860
rect 13320 8888 13326 8900
rect 17696 8888 17724 8919
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8956 19395 8959
rect 20070 8956 20076 8968
rect 19383 8928 20076 8956
rect 19383 8925 19395 8928
rect 19337 8919 19395 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 21818 8956 21824 8968
rect 21779 8928 21824 8956
rect 21818 8916 21824 8928
rect 21876 8916 21882 8968
rect 24026 8956 24032 8968
rect 21928 8928 24032 8956
rect 13320 8860 17724 8888
rect 13320 8848 13326 8860
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 18196 8860 19901 8888
rect 18196 8848 18202 8860
rect 19889 8857 19901 8860
rect 19935 8888 19947 8891
rect 21928 8888 21956 8928
rect 24026 8916 24032 8928
rect 24084 8916 24090 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24136 8928 24685 8956
rect 19935 8860 21956 8888
rect 22373 8891 22431 8897
rect 19935 8857 19947 8860
rect 19889 8851 19947 8857
rect 22373 8857 22385 8891
rect 22419 8857 22431 8891
rect 22373 8851 22431 8857
rect 5166 8820 5172 8832
rect 4080 8792 5172 8820
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5408 8792 6009 8820
rect 5408 8780 5414 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15194 8820 15200 8832
rect 15151 8792 15200 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17221 8823 17279 8829
rect 17221 8789 17233 8823
rect 17267 8820 17279 8823
rect 18156 8820 18184 8848
rect 18598 8820 18604 8832
rect 17267 8792 18184 8820
rect 18559 8792 18604 8820
rect 17267 8789 17279 8792
rect 17221 8783 17279 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19058 8820 19064 8832
rect 19019 8792 19064 8820
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 21177 8823 21235 8829
rect 21177 8789 21189 8823
rect 21223 8820 21235 8823
rect 21266 8820 21272 8832
rect 21223 8792 21272 8820
rect 21223 8789 21235 8792
rect 21177 8783 21235 8789
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 22388 8820 22416 8851
rect 24136 8832 24164 8928
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 27246 8916 27252 8968
rect 27304 8956 27310 8968
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 27304 8928 28089 8956
rect 27304 8916 27310 8928
rect 28077 8925 28089 8928
rect 28123 8956 28135 8959
rect 28166 8956 28172 8968
rect 28123 8928 28172 8956
rect 28123 8925 28135 8928
rect 28077 8919 28135 8925
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 29914 8956 29920 8968
rect 29875 8928 29920 8956
rect 29914 8916 29920 8928
rect 29972 8916 29978 8968
rect 33042 8916 33048 8968
rect 33100 8956 33106 8968
rect 33597 8959 33655 8965
rect 33597 8956 33609 8959
rect 33100 8928 33609 8956
rect 33100 8916 33106 8928
rect 33597 8925 33609 8928
rect 33643 8925 33655 8959
rect 33597 8919 33655 8925
rect 33870 8916 33876 8968
rect 33928 8956 33934 8968
rect 35345 8959 35403 8965
rect 35345 8956 35357 8959
rect 33928 8928 35357 8956
rect 33928 8916 33934 8928
rect 35345 8925 35357 8928
rect 35391 8956 35403 8959
rect 36262 8956 36268 8968
rect 35391 8928 36268 8956
rect 35391 8925 35403 8928
rect 35345 8919 35403 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 22554 8820 22560 8832
rect 21416 8792 22560 8820
rect 21416 8780 21422 8792
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 24118 8820 24124 8832
rect 24079 8792 24124 8820
rect 24118 8780 24124 8792
rect 24176 8780 24182 8832
rect 26651 8823 26709 8829
rect 26651 8789 26663 8823
rect 26697 8820 26709 8823
rect 26970 8820 26976 8832
rect 26697 8792 26976 8820
rect 26697 8789 26709 8792
rect 26651 8783 26709 8789
rect 26970 8780 26976 8792
rect 27028 8780 27034 8832
rect 31478 8820 31484 8832
rect 31439 8792 31484 8820
rect 31478 8780 31484 8792
rect 31536 8780 31542 8832
rect 32490 8820 32496 8832
rect 32451 8792 32496 8820
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 32723 8823 32781 8829
rect 32723 8789 32735 8823
rect 32769 8820 32781 8823
rect 33134 8820 33140 8832
rect 32769 8792 33140 8820
rect 32769 8789 32781 8792
rect 32723 8783 32781 8789
rect 33134 8780 33140 8792
rect 33192 8780 33198 8832
rect 33321 8823 33379 8829
rect 33321 8789 33333 8823
rect 33367 8820 33379 8823
rect 33410 8820 33416 8832
rect 33367 8792 33416 8820
rect 33367 8789 33379 8792
rect 33321 8783 33379 8789
rect 33410 8780 33416 8792
rect 33468 8780 33474 8832
rect 33594 8780 33600 8832
rect 33652 8820 33658 8832
rect 35342 8820 35348 8832
rect 33652 8792 35348 8820
rect 33652 8780 33658 8792
rect 35342 8780 35348 8792
rect 35400 8780 35406 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 3510 8576 3516 8628
rect 3568 8616 3574 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3568 8588 3985 8616
rect 3568 8576 3574 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 3973 8579 4031 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9180 8588 10824 8616
rect 9180 8576 9186 8588
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 3936 8520 5365 8548
rect 3936 8508 3942 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 5353 8511 5411 8517
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 10796 8548 10824 8588
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 10928 8588 11253 8616
rect 10928 8576 10934 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11241 8579 11299 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12158 8616 12164 8628
rect 12119 8588 12164 8616
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 13504 8588 14473 8616
rect 13504 8576 13510 8588
rect 14461 8585 14473 8588
rect 14507 8585 14519 8619
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 14461 8579 14519 8585
rect 10962 8548 10968 8560
rect 5592 8520 10272 8548
rect 10796 8520 10968 8548
rect 5592 8508 5598 8520
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3200 8452 4154 8480
rect 3200 8440 3206 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2682 8412 2688 8424
rect 1443 8384 2084 8412
rect 2643 8384 2688 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2056 8285 2084 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 4126 8412 4154 8452
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8478 8480 8484 8492
rect 8159 8452 8484 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 10244 8489 10272 8520
rect 10962 8508 10968 8520
rect 11020 8548 11026 8560
rect 12066 8548 12072 8560
rect 11020 8520 12072 8548
rect 11020 8508 11026 8520
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9631 8452 9965 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 12176 8480 12204 8576
rect 14182 8548 14188 8560
rect 13786 8520 14188 8548
rect 13786 8480 13814 8520
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 12176 8452 13584 8480
rect 10229 8443 10287 8449
rect 4430 8412 4436 8424
rect 4126 8384 4436 8412
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6687 8384 6837 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 7668 8412 7696 8440
rect 13556 8424 13584 8452
rect 13648 8452 13814 8480
rect 6871 8384 7696 8412
rect 9033 8415 9091 8421
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 12989 8415 13047 8421
rect 9079 8384 9812 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 3047 8347 3105 8353
rect 3047 8344 3059 8347
rect 2639 8316 3059 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 3047 8313 3059 8316
rect 3093 8344 3105 8347
rect 4706 8344 4712 8356
rect 3093 8316 4154 8344
rect 4664 8316 4712 8344
rect 3093 8313 3105 8316
rect 3047 8307 3105 8313
rect 2041 8279 2099 8285
rect 2041 8245 2053 8279
rect 2087 8276 2099 8279
rect 2406 8276 2412 8288
rect 2087 8248 2412 8276
rect 2087 8245 2099 8248
rect 2041 8239 2099 8245
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 3602 8276 3608 8288
rect 3563 8248 3608 8276
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 4126 8276 4154 8316
rect 4706 8304 4712 8316
rect 4764 8353 4770 8356
rect 4764 8347 4812 8353
rect 4764 8313 4766 8347
rect 4800 8313 4812 8347
rect 4764 8307 4812 8313
rect 4764 8304 4797 8307
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5776 8316 5825 8344
rect 5776 8304 5782 8316
rect 5813 8313 5825 8316
rect 5859 8344 5871 8347
rect 7190 8344 7196 8356
rect 5859 8316 7196 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 8018 8304 8024 8356
rect 8076 8344 8082 8356
rect 8434 8347 8492 8353
rect 8434 8344 8446 8347
rect 8076 8316 8446 8344
rect 8076 8304 8082 8316
rect 8434 8313 8446 8316
rect 8480 8344 8492 8347
rect 9122 8344 9128 8356
rect 8480 8316 9128 8344
rect 8480 8313 8492 8316
rect 8434 8307 8492 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 4338 8276 4344 8288
rect 4126 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8276 4402 8288
rect 4769 8276 4797 8304
rect 6178 8276 6184 8288
rect 4396 8248 4797 8276
rect 6139 8248 6184 8276
rect 4396 8236 4402 8248
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7282 8276 7288 8288
rect 6696 8248 7288 8276
rect 6696 8236 6702 8248
rect 7282 8236 7288 8248
rect 7340 8276 7346 8288
rect 7377 8279 7435 8285
rect 7377 8276 7389 8279
rect 7340 8248 7389 8276
rect 7340 8236 7346 8248
rect 7377 8245 7389 8248
rect 7423 8245 7435 8279
rect 7377 8239 7435 8245
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9784 8285 9812 8384
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13354 8412 13360 8424
rect 13035 8384 13360 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 13538 8412 13544 8424
rect 13451 8384 13544 8412
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 10100 8316 10145 8344
rect 10100 8304 10106 8316
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 12710 8344 12716 8356
rect 11204 8316 12716 8344
rect 11204 8304 11210 8316
rect 12710 8304 12716 8316
rect 12768 8344 12774 8356
rect 13648 8344 13676 8452
rect 14476 8412 14504 8579
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17644 8588 17785 8616
rect 17644 8576 17650 8588
rect 17773 8585 17785 8588
rect 17819 8616 17831 8619
rect 21358 8616 21364 8628
rect 17819 8588 21364 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 21453 8619 21511 8625
rect 21453 8585 21465 8619
rect 21499 8616 21511 8619
rect 21818 8616 21824 8628
rect 21499 8588 21824 8616
rect 21499 8585 21511 8588
rect 21453 8579 21511 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22922 8576 22928 8628
rect 22980 8616 22986 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22980 8588 23029 8616
rect 22980 8576 22986 8588
rect 23017 8585 23029 8588
rect 23063 8616 23075 8619
rect 23063 8588 23796 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 17129 8551 17187 8557
rect 17129 8517 17141 8551
rect 17175 8548 17187 8551
rect 19521 8551 19579 8557
rect 17175 8520 19057 8548
rect 17175 8517 17187 8520
rect 17129 8511 17187 8517
rect 15378 8480 15384 8492
rect 15339 8452 15384 8480
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8480 16267 8483
rect 16482 8480 16488 8492
rect 16255 8452 16488 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 19029 8480 19057 8520
rect 19521 8517 19533 8551
rect 19567 8548 19579 8551
rect 21729 8551 21787 8557
rect 21729 8548 21741 8551
rect 19567 8520 21741 8548
rect 19567 8517 19579 8520
rect 19521 8511 19579 8517
rect 21729 8517 21741 8520
rect 21775 8548 21787 8551
rect 21910 8548 21916 8560
rect 21775 8520 21916 8548
rect 21775 8517 21787 8520
rect 21729 8511 21787 8517
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 22554 8548 22560 8560
rect 22515 8520 22560 8548
rect 22554 8508 22560 8520
rect 22612 8508 22618 8560
rect 23474 8508 23480 8560
rect 23532 8548 23538 8560
rect 23532 8520 23577 8548
rect 23532 8508 23538 8520
rect 19426 8480 19432 8492
rect 19029 8452 19432 8480
rect 19426 8440 19432 8452
rect 19484 8480 19490 8492
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 19484 8452 19809 8480
rect 19484 8440 19490 8452
rect 19797 8449 19809 8452
rect 19843 8480 19855 8483
rect 21928 8480 21956 8508
rect 23768 8489 23796 8588
rect 26326 8576 26332 8628
rect 26384 8616 26390 8628
rect 26513 8619 26571 8625
rect 26513 8616 26525 8619
rect 26384 8588 26525 8616
rect 26384 8576 26390 8588
rect 26513 8585 26525 8588
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 27522 8576 27528 8628
rect 27580 8616 27586 8628
rect 28261 8619 28319 8625
rect 28261 8616 28273 8619
rect 27580 8588 28273 8616
rect 27580 8576 27586 8588
rect 28261 8585 28273 8588
rect 28307 8585 28319 8619
rect 28994 8616 29000 8628
rect 28955 8588 29000 8616
rect 28261 8579 28319 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 32306 8616 32312 8628
rect 32267 8588 32312 8616
rect 32306 8576 32312 8588
rect 32364 8576 32370 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32677 8619 32735 8625
rect 32677 8616 32689 8619
rect 32548 8588 32689 8616
rect 32548 8576 32554 8588
rect 32677 8585 32689 8588
rect 32723 8616 32735 8619
rect 33594 8616 33600 8628
rect 32723 8588 33600 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 33594 8576 33600 8588
rect 33652 8576 33658 8628
rect 35250 8616 35256 8628
rect 34164 8588 35256 8616
rect 23753 8483 23811 8489
rect 19843 8452 21220 8480
rect 21928 8452 23612 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14476 8384 14657 8412
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 15102 8412 15108 8424
rect 15063 8384 15108 8412
rect 14645 8375 14703 8381
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 18598 8412 18604 8424
rect 17184 8384 18604 8412
rect 17184 8372 17190 8384
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 12768 8316 13676 8344
rect 13817 8347 13875 8353
rect 12768 8304 12774 8316
rect 13817 8313 13829 8347
rect 13863 8344 13875 8347
rect 15286 8344 15292 8356
rect 13863 8316 15292 8344
rect 13863 8313 13875 8316
rect 13817 8307 13875 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 15930 8344 15936 8356
rect 15795 8316 15936 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 15930 8304 15936 8316
rect 15988 8344 15994 8356
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15988 8316 16129 8344
rect 15988 8304 15994 8316
rect 16117 8313 16129 8316
rect 16163 8344 16175 8347
rect 16571 8347 16629 8353
rect 16571 8344 16583 8347
rect 16163 8316 16583 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 16571 8313 16583 8316
rect 16617 8344 16629 8347
rect 18922 8347 18980 8353
rect 18922 8344 18934 8347
rect 16617 8316 18934 8344
rect 16617 8313 16629 8316
rect 16571 8307 16629 8313
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 8628 8248 9321 8276
rect 8628 8236 8634 8248
rect 9309 8245 9321 8248
rect 9355 8276 9367 8279
rect 9585 8279 9643 8285
rect 9585 8276 9597 8279
rect 9355 8248 9597 8276
rect 9355 8245 9367 8248
rect 9309 8239 9367 8245
rect 9585 8245 9597 8248
rect 9631 8245 9643 8279
rect 9585 8239 9643 8245
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8276 9827 8279
rect 10060 8276 10088 8304
rect 18616 8288 18644 8316
rect 18922 8313 18934 8316
rect 18968 8313 18980 8347
rect 20438 8344 20444 8356
rect 20399 8316 20444 8344
rect 18922 8307 18980 8313
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 20588 8316 20633 8344
rect 20588 8304 20594 8316
rect 9815 8248 10088 8276
rect 18509 8279 18567 8285
rect 9815 8245 9827 8248
rect 9769 8239 9827 8245
rect 18509 8245 18521 8279
rect 18555 8276 18567 8279
rect 18598 8276 18604 8288
rect 18555 8248 18604 8276
rect 18555 8245 18567 8248
rect 18509 8239 18567 8245
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 20254 8276 20260 8288
rect 20215 8248 20260 8276
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 21192 8276 21220 8452
rect 21269 8347 21327 8353
rect 21269 8313 21281 8347
rect 21315 8344 21327 8347
rect 21358 8344 21364 8356
rect 21315 8316 21364 8344
rect 21315 8313 21327 8316
rect 21269 8307 21327 8313
rect 21358 8304 21364 8316
rect 21416 8304 21422 8356
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 22005 8347 22063 8353
rect 22005 8344 22017 8347
rect 21784 8316 22017 8344
rect 21784 8304 21790 8316
rect 22005 8313 22017 8316
rect 22051 8313 22063 8347
rect 22005 8307 22063 8313
rect 22097 8347 22155 8353
rect 22097 8313 22109 8347
rect 22143 8313 22155 8347
rect 22097 8307 22155 8313
rect 21910 8276 21916 8288
rect 21192 8248 21916 8276
rect 21910 8236 21916 8248
rect 21968 8276 21974 8288
rect 22112 8276 22140 8307
rect 21968 8248 22140 8276
rect 23584 8276 23612 8452
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 24026 8480 24032 8492
rect 23987 8452 24032 8480
rect 23753 8443 23811 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 25317 8483 25375 8489
rect 25317 8449 25329 8483
rect 25363 8480 25375 8483
rect 25406 8480 25412 8492
rect 25363 8452 25412 8480
rect 25363 8449 25375 8452
rect 25317 8443 25375 8449
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 27062 8480 27068 8492
rect 27023 8452 27068 8480
rect 27062 8440 27068 8452
rect 27120 8440 27126 8492
rect 29012 8480 29040 8576
rect 30561 8483 30619 8489
rect 29012 8452 30328 8480
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 26418 8412 26424 8424
rect 24636 8384 26424 8412
rect 24636 8372 24642 8384
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 29086 8412 29092 8424
rect 26476 8384 29092 8412
rect 26476 8372 26482 8384
rect 29086 8372 29092 8384
rect 29144 8412 29150 8424
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 29144 8384 29837 8412
rect 29144 8372 29150 8384
rect 29825 8381 29837 8384
rect 29871 8412 29883 8415
rect 30006 8412 30012 8424
rect 29871 8384 30012 8412
rect 29871 8381 29883 8384
rect 29825 8375 29883 8381
rect 30006 8372 30012 8384
rect 30064 8372 30070 8424
rect 30300 8421 30328 8452
rect 30561 8449 30573 8483
rect 30607 8480 30619 8483
rect 31478 8480 31484 8492
rect 30607 8452 31484 8480
rect 30607 8449 30619 8452
rect 30561 8443 30619 8449
rect 31478 8440 31484 8452
rect 31536 8440 31542 8492
rect 32950 8440 32956 8492
rect 33008 8480 33014 8492
rect 33321 8483 33379 8489
rect 33321 8480 33333 8483
rect 33008 8452 33333 8480
rect 33008 8440 33014 8452
rect 33321 8449 33333 8452
rect 33367 8480 33379 8483
rect 34164 8480 34192 8588
rect 35250 8576 35256 8588
rect 35308 8576 35314 8628
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 34333 8551 34391 8557
rect 34333 8517 34345 8551
rect 34379 8548 34391 8551
rect 34606 8548 34612 8560
rect 34379 8520 34612 8548
rect 34379 8517 34391 8520
rect 34333 8511 34391 8517
rect 34606 8508 34612 8520
rect 34664 8508 34670 8560
rect 34882 8508 34888 8560
rect 34940 8548 34946 8560
rect 35529 8551 35587 8557
rect 35529 8548 35541 8551
rect 34940 8520 35541 8548
rect 34940 8508 34946 8520
rect 35529 8517 35541 8520
rect 35575 8548 35587 8551
rect 37182 8548 37188 8560
rect 35575 8520 37188 8548
rect 35575 8517 35587 8520
rect 35529 8511 35587 8517
rect 37182 8508 37188 8520
rect 37240 8508 37246 8560
rect 34974 8480 34980 8492
rect 33367 8452 34192 8480
rect 34935 8452 34980 8480
rect 33367 8449 33379 8452
rect 33321 8443 33379 8449
rect 34974 8440 34980 8452
rect 35032 8440 35038 8492
rect 35710 8440 35716 8492
rect 35768 8480 35774 8492
rect 36817 8483 36875 8489
rect 36817 8480 36829 8483
rect 35768 8452 36829 8480
rect 35768 8440 35774 8452
rect 36817 8449 36829 8452
rect 36863 8449 36875 8483
rect 36817 8443 36875 8449
rect 30285 8415 30343 8421
rect 30285 8381 30297 8415
rect 30331 8412 30343 8415
rect 30834 8412 30840 8424
rect 30331 8384 30840 8412
rect 30331 8381 30343 8384
rect 30285 8375 30343 8381
rect 30834 8372 30840 8384
rect 30892 8372 30898 8424
rect 30929 8415 30987 8421
rect 30929 8381 30941 8415
rect 30975 8412 30987 8415
rect 31294 8412 31300 8424
rect 30975 8384 31300 8412
rect 30975 8381 30987 8384
rect 30929 8375 30987 8381
rect 31294 8372 31300 8384
rect 31352 8412 31358 8424
rect 31389 8415 31447 8421
rect 31389 8412 31401 8415
rect 31352 8384 31401 8412
rect 31352 8372 31358 8384
rect 31389 8381 31401 8384
rect 31435 8381 31447 8415
rect 31389 8375 31447 8381
rect 23750 8304 23756 8356
rect 23808 8344 23814 8356
rect 23845 8347 23903 8353
rect 23845 8344 23857 8347
rect 23808 8316 23857 8344
rect 23808 8304 23814 8316
rect 23845 8313 23857 8316
rect 23891 8313 23903 8347
rect 23845 8307 23903 8313
rect 24765 8347 24823 8353
rect 24765 8313 24777 8347
rect 24811 8344 24823 8347
rect 25038 8344 25044 8356
rect 24811 8316 25044 8344
rect 24811 8313 24823 8316
rect 24765 8307 24823 8313
rect 25038 8304 25044 8316
rect 25096 8344 25102 8356
rect 25225 8347 25283 8353
rect 25225 8344 25237 8347
rect 25096 8316 25237 8344
rect 25096 8304 25102 8316
rect 25225 8313 25237 8316
rect 25271 8344 25283 8347
rect 25679 8347 25737 8353
rect 25679 8344 25691 8347
rect 25271 8316 25691 8344
rect 25271 8313 25283 8316
rect 25225 8307 25283 8313
rect 25679 8313 25691 8316
rect 25725 8344 25737 8347
rect 26510 8344 26516 8356
rect 25725 8316 26516 8344
rect 25725 8313 25737 8316
rect 25679 8307 25737 8313
rect 26510 8304 26516 8316
rect 26568 8344 26574 8356
rect 27386 8347 27444 8353
rect 27386 8344 27398 8347
rect 26568 8316 27398 8344
rect 26568 8304 26574 8316
rect 24394 8276 24400 8288
rect 23584 8248 24400 8276
rect 21968 8236 21974 8248
rect 24394 8236 24400 8248
rect 24452 8236 24458 8288
rect 26234 8276 26240 8288
rect 26195 8248 26240 8276
rect 26234 8236 26240 8248
rect 26292 8236 26298 8288
rect 26988 8285 27016 8316
rect 27386 8313 27398 8316
rect 27432 8344 27444 8347
rect 31570 8344 31576 8356
rect 27432 8316 28994 8344
rect 27432 8313 27444 8316
rect 27386 8307 27444 8313
rect 26973 8279 27031 8285
rect 26973 8245 26985 8279
rect 27019 8276 27031 8279
rect 27062 8276 27068 8288
rect 27019 8248 27068 8276
rect 27019 8245 27031 8248
rect 26973 8239 27031 8245
rect 27062 8236 27068 8248
rect 27120 8236 27126 8288
rect 27982 8276 27988 8288
rect 27943 8248 27988 8276
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 28966 8276 28994 8316
rect 31312 8316 31576 8344
rect 31312 8285 31340 8316
rect 31570 8304 31576 8316
rect 31628 8344 31634 8356
rect 31751 8347 31809 8353
rect 31751 8344 31763 8347
rect 31628 8316 31763 8344
rect 31628 8304 31634 8316
rect 31751 8313 31763 8316
rect 31797 8344 31809 8347
rect 33318 8344 33324 8356
rect 31797 8316 33324 8344
rect 31797 8313 31809 8316
rect 31751 8307 31809 8313
rect 33318 8304 33324 8316
rect 33376 8304 33382 8356
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 33962 8344 33968 8356
rect 33468 8316 33513 8344
rect 33923 8316 33968 8344
rect 33468 8304 33474 8316
rect 33962 8304 33968 8316
rect 34020 8304 34026 8356
rect 34701 8347 34759 8353
rect 34701 8313 34713 8347
rect 34747 8344 34759 8347
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34747 8316 35081 8344
rect 34747 8313 34759 8316
rect 34701 8307 34759 8313
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 36170 8344 36176 8356
rect 35069 8307 35127 8313
rect 35728 8316 36176 8344
rect 29733 8279 29791 8285
rect 29733 8276 29745 8279
rect 28966 8248 29745 8276
rect 29733 8245 29745 8248
rect 29779 8276 29791 8279
rect 31297 8279 31355 8285
rect 31297 8276 31309 8279
rect 29779 8248 31309 8276
rect 29779 8245 29791 8248
rect 29733 8239 29791 8245
rect 31297 8245 31309 8248
rect 31343 8245 31355 8279
rect 33042 8276 33048 8288
rect 33003 8248 33048 8276
rect 31297 8239 31355 8245
rect 33042 8236 33048 8248
rect 33100 8236 33106 8288
rect 35084 8276 35112 8307
rect 35728 8276 35756 8316
rect 36170 8304 36176 8316
rect 36228 8304 36234 8356
rect 36538 8344 36544 8356
rect 36499 8316 36544 8344
rect 36538 8304 36544 8316
rect 36596 8304 36602 8356
rect 36630 8304 36636 8356
rect 36688 8344 36694 8356
rect 36688 8316 36733 8344
rect 36688 8304 36694 8316
rect 35894 8276 35900 8288
rect 35084 8248 35756 8276
rect 35855 8248 35900 8276
rect 35894 8236 35900 8248
rect 35952 8236 35958 8288
rect 36556 8276 36584 8304
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 36556 8248 37473 8276
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8072 2746 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2740 8044 3433 8072
rect 2740 8032 2746 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3421 8035 3479 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4488 8044 5089 8072
rect 4488 8032 4494 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 7190 8072 7196 8084
rect 6880 8044 7196 8072
rect 6880 8032 6886 8044
rect 7190 8032 7196 8044
rect 7248 8072 7254 8084
rect 12618 8072 12624 8084
rect 7248 8044 11560 8072
rect 12579 8044 12624 8072
rect 7248 8032 7254 8044
rect 1854 8004 1860 8016
rect 1412 7976 1860 8004
rect 1412 7945 1440 7976
rect 1854 7964 1860 7976
rect 1912 8004 1918 8016
rect 2498 8004 2504 8016
rect 1912 7976 2504 8004
rect 1912 7964 1918 7976
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 3050 8004 3056 8016
rect 2700 7976 3056 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 1397 7899 1455 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2700 7945 2728 7976
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 3602 7964 3608 8016
rect 3660 8004 3666 8016
rect 4246 8004 4252 8016
rect 3660 7976 4252 8004
rect 3660 7964 3666 7976
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 4798 8004 4804 8016
rect 4759 7976 4804 8004
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10137 8007 10195 8013
rect 10137 8004 10149 8007
rect 10100 7976 10149 8004
rect 10100 7964 10106 7976
rect 10137 7973 10149 7976
rect 10183 8004 10195 8007
rect 11333 8007 11391 8013
rect 11333 8004 11345 8007
rect 10183 7976 11345 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 11333 7973 11345 7976
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7905 2743 7939
rect 2958 7936 2964 7948
rect 2871 7908 2964 7936
rect 2685 7899 2743 7905
rect 2958 7896 2964 7908
rect 3016 7936 3022 7948
rect 3510 7936 3516 7948
rect 3016 7908 3516 7936
rect 3016 7896 3022 7908
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6144 7908 6193 7936
rect 6144 7896 6150 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 11532 7945 11560 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15344 8044 15485 8072
rect 15344 8032 15350 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 22462 8072 22468 8084
rect 19659 8044 22468 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 22462 8032 22468 8044
rect 22520 8072 22526 8084
rect 22520 8044 22692 8072
rect 22520 8032 22526 8044
rect 12066 7964 12072 8016
rect 12124 8004 12130 8016
rect 13218 8007 13276 8013
rect 13218 8004 13230 8007
rect 12124 7976 13230 8004
rect 12124 7964 12130 7976
rect 13218 7973 13230 7976
rect 13264 7973 13276 8007
rect 13218 7967 13276 7973
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 14645 8007 14703 8013
rect 14645 8004 14657 8007
rect 13596 7976 14657 8004
rect 13596 7964 13602 7976
rect 14645 7973 14657 7976
rect 14691 8004 14703 8007
rect 15102 8004 15108 8016
rect 14691 7976 15108 8004
rect 14691 7973 14703 7976
rect 14645 7967 14703 7973
rect 15102 7964 15108 7976
rect 15160 8004 15166 8016
rect 15160 7976 16344 8004
rect 15160 7964 15166 7976
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 7524 7908 7665 7936
rect 7524 7896 7530 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7936 11575 7939
rect 11606 7936 11612 7948
rect 11563 7908 11612 7936
rect 11563 7905 11575 7908
rect 11517 7899 11575 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 11790 7936 11796 7948
rect 11747 7908 11796 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16316 7945 16344 7976
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 16577 8007 16635 8013
rect 16577 8004 16589 8007
rect 16540 7976 16589 8004
rect 16540 7964 16546 7976
rect 16577 7973 16589 7976
rect 16623 7973 16635 8007
rect 16577 7967 16635 7973
rect 18598 7964 18604 8016
rect 18656 8004 18662 8016
rect 19014 8007 19072 8013
rect 19014 8004 19026 8007
rect 18656 7976 19026 8004
rect 18656 7964 18662 7976
rect 19014 7973 19026 7976
rect 19060 7973 19072 8007
rect 19014 7967 19072 7973
rect 19981 8007 20039 8013
rect 19981 7973 19993 8007
rect 20027 8004 20039 8007
rect 20070 8004 20076 8016
rect 20027 7976 20076 8004
rect 20027 7973 20039 7976
rect 19981 7967 20039 7973
rect 20070 7964 20076 7976
rect 20128 7964 20134 8016
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 20530 8004 20536 8016
rect 20312 7976 20536 8004
rect 20312 7964 20318 7976
rect 20530 7964 20536 7976
rect 20588 8004 20594 8016
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 20588 7976 21097 8004
rect 20588 7964 20594 7976
rect 21085 7973 21097 7976
rect 21131 7973 21143 8007
rect 21910 8004 21916 8016
rect 21871 7976 21916 8004
rect 21085 7967 21143 7973
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 22664 8013 22692 8044
rect 23198 8032 23204 8084
rect 23256 8072 23262 8084
rect 25406 8072 25412 8084
rect 23256 8044 24164 8072
rect 25367 8044 25412 8072
rect 23256 8032 23262 8044
rect 22649 8007 22707 8013
rect 22649 7973 22661 8007
rect 22695 8004 22707 8007
rect 23750 8004 23756 8016
rect 22695 7976 23756 8004
rect 22695 7973 22707 7976
rect 22649 7967 22707 7973
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 24136 8013 24164 8044
rect 25406 8032 25412 8044
rect 25464 8032 25470 8084
rect 27801 8075 27859 8081
rect 27801 8041 27813 8075
rect 27847 8072 27859 8075
rect 27982 8072 27988 8084
rect 27847 8044 27988 8072
rect 27847 8041 27859 8044
rect 27801 8035 27859 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 28813 8075 28871 8081
rect 28813 8041 28825 8075
rect 28859 8072 28871 8075
rect 28994 8072 29000 8084
rect 28859 8044 29000 8072
rect 28859 8041 28871 8044
rect 28813 8035 28871 8041
rect 28994 8032 29000 8044
rect 29052 8032 29058 8084
rect 30006 8072 30012 8084
rect 29967 8044 30012 8072
rect 30006 8032 30012 8044
rect 30064 8032 30070 8084
rect 32950 8072 32956 8084
rect 32911 8044 32956 8072
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 33318 8032 33324 8084
rect 33376 8072 33382 8084
rect 33413 8075 33471 8081
rect 33413 8072 33425 8075
rect 33376 8044 33425 8072
rect 33376 8032 33382 8044
rect 33413 8041 33425 8044
rect 33459 8041 33471 8075
rect 33413 8035 33471 8041
rect 36633 8075 36691 8081
rect 36633 8041 36645 8075
rect 36679 8072 36691 8075
rect 37734 8072 37740 8084
rect 36679 8044 37740 8072
rect 36679 8041 36691 8044
rect 36633 8035 36691 8041
rect 37734 8032 37740 8044
rect 37792 8032 37798 8084
rect 24121 8007 24179 8013
rect 24121 7973 24133 8007
rect 24167 7973 24179 8007
rect 24121 7967 24179 7973
rect 24213 8007 24271 8013
rect 24213 7973 24225 8007
rect 24259 8004 24271 8007
rect 24394 8004 24400 8016
rect 24259 7976 24400 8004
rect 24259 7973 24271 7976
rect 24213 7967 24271 7973
rect 24394 7964 24400 7976
rect 24452 7964 24458 8016
rect 26234 7964 26240 8016
rect 26292 8004 26298 8016
rect 26697 8007 26755 8013
rect 26697 8004 26709 8007
rect 26292 7976 26709 8004
rect 26292 7964 26298 7976
rect 26697 7973 26709 7976
rect 26743 8004 26755 8007
rect 26786 8004 26792 8016
rect 26743 7976 26792 8004
rect 26743 7973 26755 7976
rect 26697 7967 26755 7973
rect 26786 7964 26792 7976
rect 26844 7964 26850 8016
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15804 7908 15853 7936
rect 15804 7896 15810 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7936 16359 7939
rect 16850 7936 16856 7948
rect 16347 7908 16856 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17368 7908 17417 7936
rect 17368 7896 17374 7908
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 21726 7896 21732 7948
rect 21784 7936 21790 7948
rect 22281 7939 22339 7945
rect 22281 7936 22293 7939
rect 21784 7908 22293 7936
rect 21784 7896 21790 7908
rect 22281 7905 22293 7908
rect 22327 7905 22339 7939
rect 28902 7936 28908 7948
rect 28863 7908 28908 7936
rect 22281 7899 22339 7905
rect 28902 7896 28908 7908
rect 28960 7896 28966 7948
rect 29012 7936 29040 8032
rect 29641 8007 29699 8013
rect 29641 7973 29653 8007
rect 29687 8004 29699 8007
rect 29914 8004 29920 8016
rect 29687 7976 29920 8004
rect 29687 7973 29699 7976
rect 29641 7967 29699 7973
rect 29914 7964 29920 7976
rect 29972 8004 29978 8016
rect 30285 8007 30343 8013
rect 30285 8004 30297 8007
rect 29972 7976 30297 8004
rect 29972 7964 29978 7976
rect 30285 7973 30297 7976
rect 30331 7973 30343 8007
rect 30285 7967 30343 7973
rect 31205 8007 31263 8013
rect 31205 7973 31217 8007
rect 31251 8004 31263 8007
rect 33042 8004 33048 8016
rect 31251 7976 33048 8004
rect 31251 7973 31263 7976
rect 31205 7967 31263 7973
rect 33042 7964 33048 7976
rect 33100 7964 33106 8016
rect 35066 8004 35072 8016
rect 35027 7976 35072 8004
rect 35066 7964 35072 7976
rect 35124 7964 35130 8016
rect 29365 7939 29423 7945
rect 29365 7936 29377 7939
rect 29012 7908 29377 7936
rect 29365 7905 29377 7908
rect 29411 7905 29423 7939
rect 30466 7936 30472 7948
rect 30427 7908 30472 7936
rect 29365 7899 29423 7905
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 30834 7896 30840 7948
rect 30892 7936 30898 7948
rect 30929 7939 30987 7945
rect 30929 7936 30941 7939
rect 30892 7908 30941 7936
rect 30892 7896 30898 7908
rect 30929 7905 30941 7908
rect 30975 7905 30987 7939
rect 30929 7899 30987 7905
rect 36262 7896 36268 7948
rect 36320 7936 36326 7948
rect 36449 7939 36507 7945
rect 36449 7936 36461 7939
rect 36320 7908 36461 7936
rect 36320 7896 36326 7908
rect 36449 7905 36461 7908
rect 36495 7905 36507 7939
rect 36449 7899 36507 7905
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5534 7868 5540 7880
rect 4212 7840 5540 7868
rect 4212 7828 4218 7840
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 6914 7868 6920 7880
rect 6871 7840 6920 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8110 7868 8116 7880
rect 8067 7840 8116 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8846 7868 8852 7880
rect 8803 7840 8852 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10134 7868 10140 7880
rect 10091 7840 10140 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 12894 7868 12900 7880
rect 12855 7840 12900 7868
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20404 7840 21005 7868
rect 20404 7828 20410 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 21818 7868 21824 7880
rect 21683 7840 21824 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22060 7840 22569 7868
rect 22060 7828 22066 7840
rect 22557 7837 22569 7840
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 22646 7828 22652 7880
rect 22704 7868 22710 7880
rect 22833 7871 22891 7877
rect 22833 7868 22845 7871
rect 22704 7840 22845 7868
rect 22704 7828 22710 7840
rect 22833 7837 22845 7840
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 24397 7871 24455 7877
rect 24397 7837 24409 7871
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2314 7800 2320 7812
rect 1627 7772 2320 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2314 7760 2320 7772
rect 2372 7760 2378 7812
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7791 7803 7849 7809
rect 7791 7800 7803 7803
rect 7248 7772 7803 7800
rect 7248 7760 7254 7772
rect 7791 7769 7803 7772
rect 7837 7769 7849 7803
rect 7791 7763 7849 7769
rect 18874 7760 18880 7812
rect 18932 7800 18938 7812
rect 20438 7800 20444 7812
rect 18932 7772 20444 7800
rect 18932 7760 18938 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 24026 7760 24032 7812
rect 24084 7800 24090 7812
rect 24412 7800 24440 7831
rect 26326 7828 26332 7880
rect 26384 7868 26390 7880
rect 26605 7871 26663 7877
rect 26605 7868 26617 7871
rect 26384 7840 26617 7868
rect 26384 7828 26390 7840
rect 26605 7837 26617 7840
rect 26651 7837 26663 7871
rect 27246 7868 27252 7880
rect 27207 7840 27252 7868
rect 26605 7831 26663 7837
rect 27246 7828 27252 7840
rect 27304 7828 27310 7880
rect 33042 7868 33048 7880
rect 33003 7840 33048 7868
rect 33042 7828 33048 7840
rect 33100 7828 33106 7880
rect 33962 7828 33968 7880
rect 34020 7868 34026 7880
rect 34425 7871 34483 7877
rect 34425 7868 34437 7871
rect 34020 7840 34437 7868
rect 34020 7828 34026 7840
rect 34425 7837 34437 7840
rect 34471 7868 34483 7871
rect 34977 7871 35035 7877
rect 34977 7868 34989 7871
rect 34471 7840 34989 7868
rect 34471 7837 34483 7840
rect 34425 7831 34483 7837
rect 34977 7837 34989 7840
rect 35023 7868 35035 7871
rect 35710 7868 35716 7880
rect 35023 7840 35716 7868
rect 35023 7837 35035 7840
rect 34977 7831 35035 7837
rect 35710 7828 35716 7840
rect 35768 7828 35774 7880
rect 35526 7800 35532 7812
rect 24084 7772 24440 7800
rect 35487 7772 35532 7800
rect 24084 7760 24090 7772
rect 35526 7760 35532 7772
rect 35584 7760 35590 7812
rect 7466 7732 7472 7744
rect 7427 7704 7472 7732
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8018 7732 8024 7744
rect 7975 7704 8024 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 8812 7704 9229 7732
rect 8812 7692 8818 7704
rect 9217 7701 9229 7704
rect 9263 7732 9275 7735
rect 9306 7732 9312 7744
rect 9263 7704 9312 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11112 7704 11805 7732
rect 11112 7692 11118 7704
rect 11793 7701 11805 7704
rect 11839 7701 11851 7735
rect 11793 7695 11851 7701
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 17589 7735 17647 7741
rect 13872 7704 13917 7732
rect 13872 7692 13878 7704
rect 17589 7701 17601 7735
rect 17635 7732 17647 7735
rect 18506 7732 18512 7744
rect 17635 7704 18512 7732
rect 17635 7701 17647 7704
rect 17589 7695 17647 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 33965 7735 34023 7741
rect 33965 7701 33977 7735
rect 34011 7732 34023 7735
rect 34146 7732 34152 7744
rect 34011 7704 34152 7732
rect 34011 7701 34023 7704
rect 33965 7695 34023 7701
rect 34146 7692 34152 7704
rect 34204 7692 34210 7744
rect 34793 7735 34851 7741
rect 34793 7701 34805 7735
rect 34839 7732 34851 7735
rect 35250 7732 35256 7744
rect 34839 7704 35256 7732
rect 34839 7701 34851 7704
rect 34793 7695 34851 7701
rect 35250 7692 35256 7704
rect 35308 7692 35314 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 2958 7528 2964 7540
rect 1811 7500 2964 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3421 7531 3479 7537
rect 3421 7528 3433 7531
rect 3108 7500 3433 7528
rect 3108 7488 3114 7500
rect 3421 7497 3433 7500
rect 3467 7497 3479 7531
rect 3421 7491 3479 7497
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 4304 7500 5549 7528
rect 4304 7488 4310 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 5859 7531 5917 7537
rect 5859 7497 5871 7531
rect 5905 7528 5917 7531
rect 8570 7528 8576 7540
rect 5905 7500 8576 7528
rect 5905 7497 5917 7500
rect 5859 7491 5917 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 9088 7500 9689 7528
rect 9088 7488 9094 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 15470 7528 15476 7540
rect 11296 7500 15476 7528
rect 11296 7488 11302 7500
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15804 7500 15853 7528
rect 15804 7488 15810 7500
rect 15841 7497 15853 7500
rect 15887 7528 15899 7531
rect 18046 7528 18052 7540
rect 15887 7500 18052 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7528 18291 7531
rect 19058 7528 19064 7540
rect 18279 7500 19064 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 20254 7528 20260 7540
rect 20027 7500 20260 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20254 7488 20260 7500
rect 20312 7528 20318 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20312 7500 20913 7528
rect 20312 7488 20318 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 22462 7528 22468 7540
rect 22423 7500 22468 7528
rect 20901 7491 20959 7497
rect 22462 7488 22468 7500
rect 22520 7488 22526 7540
rect 23109 7531 23167 7537
rect 23109 7497 23121 7531
rect 23155 7528 23167 7531
rect 23198 7528 23204 7540
rect 23155 7500 23204 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 26786 7528 26792 7540
rect 26747 7500 26792 7528
rect 26786 7488 26792 7500
rect 26844 7488 26850 7540
rect 29086 7528 29092 7540
rect 29047 7500 29092 7528
rect 29086 7488 29092 7500
rect 29144 7488 29150 7540
rect 30466 7528 30472 7540
rect 30427 7500 30472 7528
rect 30466 7488 30472 7500
rect 30524 7488 30530 7540
rect 34146 7488 34152 7540
rect 34204 7528 34210 7540
rect 34517 7531 34575 7537
rect 34517 7528 34529 7531
rect 34204 7500 34529 7528
rect 34204 7488 34210 7500
rect 34517 7497 34529 7500
rect 34563 7528 34575 7531
rect 34609 7531 34667 7537
rect 34609 7528 34621 7531
rect 34563 7500 34621 7528
rect 34563 7497 34575 7500
rect 34517 7491 34575 7497
rect 34609 7497 34621 7500
rect 34655 7497 34667 7531
rect 34609 7491 34667 7497
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 6144 7432 6193 7460
rect 6144 7420 6150 7432
rect 6181 7429 6193 7432
rect 6227 7460 6239 7463
rect 6454 7460 6460 7472
rect 6227 7432 6460 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 6454 7420 6460 7432
rect 6512 7460 6518 7472
rect 7926 7460 7932 7472
rect 6512 7432 7932 7460
rect 6512 7420 6518 7432
rect 7926 7420 7932 7432
rect 7984 7460 7990 7472
rect 8665 7463 8723 7469
rect 8665 7460 8677 7463
rect 7984 7432 8677 7460
rect 7984 7420 7990 7432
rect 8665 7429 8677 7432
rect 8711 7460 8723 7463
rect 9125 7463 9183 7469
rect 9125 7460 9137 7463
rect 8711 7432 9137 7460
rect 8711 7429 8723 7432
rect 8665 7423 8723 7429
rect 9125 7429 9137 7432
rect 9171 7429 9183 7463
rect 9125 7423 9183 7429
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9364 7432 9505 7460
rect 9364 7420 9370 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 13722 7460 13728 7472
rect 9493 7423 9551 7429
rect 11256 7432 13728 7460
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 8021 7395 8079 7401
rect 6687 7364 7925 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3016 7296 3985 7324
rect 3016 7284 3022 7296
rect 3973 7293 3985 7296
rect 4019 7324 4031 7327
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4019 7296 5181 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 5788 7327 5846 7333
rect 5788 7293 5800 7327
rect 5834 7324 5846 7327
rect 6656 7324 6684 7355
rect 7800 7327 7858 7333
rect 7800 7324 7812 7327
rect 5834 7296 6684 7324
rect 7484 7296 7812 7324
rect 5834 7293 5846 7296
rect 5788 7287 5846 7293
rect 4338 7265 4344 7268
rect 2133 7259 2191 7265
rect 2133 7225 2145 7259
rect 2179 7256 2191 7259
rect 2546 7259 2604 7265
rect 2546 7256 2558 7259
rect 2179 7228 2558 7256
rect 2179 7225 2191 7228
rect 2133 7219 2191 7225
rect 2546 7225 2558 7228
rect 2592 7256 2604 7259
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 2592 7228 3801 7256
rect 2592 7225 2604 7228
rect 2546 7219 2604 7225
rect 3789 7225 3801 7228
rect 3835 7256 3847 7259
rect 4335 7256 4344 7265
rect 3835 7228 4344 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4335 7219 4344 7228
rect 4338 7216 4344 7219
rect 4396 7216 4402 7268
rect 3142 7188 3148 7200
rect 3103 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 4890 7188 4896 7200
rect 4851 7160 4896 7188
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7188 7254 7200
rect 7484 7197 7512 7296
rect 7800 7293 7812 7296
rect 7846 7293 7858 7327
rect 7897 7324 7925 7364
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8110 7392 8116 7404
rect 8067 7364 8116 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 9214 7392 9220 7404
rect 8435 7364 9220 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9582 7392 9588 7404
rect 9543 7364 9588 7392
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 11256 7392 11284 7432
rect 13722 7420 13728 7432
rect 13780 7460 13786 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 13780 7432 14473 7460
rect 13780 7420 13786 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 17770 7460 17776 7472
rect 17731 7432 17776 7460
rect 14461 7423 14519 7429
rect 11514 7392 11520 7404
rect 11072 7364 11284 7392
rect 11475 7364 11520 7392
rect 8202 7324 8208 7336
rect 7897 7296 8208 7324
rect 7800 7287 7858 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9364 7327 9422 7333
rect 9364 7324 9376 7327
rect 8720 7296 9376 7324
rect 8720 7284 8726 7296
rect 9364 7293 9376 7296
rect 9410 7293 9422 7327
rect 9364 7287 9422 7293
rect 7650 7256 7656 7268
rect 7563 7228 7656 7256
rect 7650 7216 7656 7228
rect 7708 7256 7714 7268
rect 8846 7256 8852 7268
rect 7708 7228 8852 7256
rect 7708 7216 7714 7228
rect 8846 7216 8852 7228
rect 8904 7256 8910 7268
rect 9217 7259 9275 7265
rect 9217 7256 9229 7259
rect 8904 7228 9229 7256
rect 8904 7216 8910 7228
rect 9217 7225 9229 7228
rect 9263 7225 9275 7259
rect 9379 7256 9407 7287
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11072 7333 11100 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11790 7392 11796 7404
rect 11751 7364 11796 7392
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10928 7296 11069 7324
rect 10928 7284 10934 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 11204 7296 11253 7324
rect 11204 7284 11210 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12216 7296 12449 7324
rect 12216 7284 12222 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 12437 7287 12495 7293
rect 12773 7296 13645 7324
rect 12773 7265 12801 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 14476 7324 14504 7423
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 19076 7460 19104 7488
rect 23385 7463 23443 7469
rect 23385 7460 23397 7463
rect 19076 7432 23397 7460
rect 23385 7429 23397 7432
rect 23431 7460 23443 7463
rect 23431 7432 24532 7460
rect 23431 7429 23443 7432
rect 23385 7423 23443 7429
rect 15194 7392 15200 7404
rect 15155 7364 15200 7392
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 17126 7392 17132 7404
rect 17087 7364 17132 7392
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14476 7296 14657 7324
rect 13633 7287 13691 7293
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 15102 7324 15108 7336
rect 15063 7296 15108 7324
rect 14645 7287 14703 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16666 7324 16672 7336
rect 16347 7296 16672 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16850 7324 16856 7336
rect 16811 7296 16856 7324
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17788 7324 17816 7420
rect 18598 7392 18604 7404
rect 18511 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7392 18662 7404
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18656 7364 18981 7392
rect 18656 7352 18662 7364
rect 18969 7361 18981 7364
rect 19015 7392 19027 7395
rect 21266 7392 21272 7404
rect 19015 7364 21272 7392
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17788 7296 18061 7324
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 18782 7284 18788 7336
rect 18840 7324 18846 7336
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18840 7296 19073 7324
rect 18840 7284 18846 7296
rect 19061 7293 19073 7296
rect 19107 7293 19119 7327
rect 19061 7287 19119 7293
rect 10229 7259 10287 7265
rect 10229 7256 10241 7259
rect 9379 7228 10241 7256
rect 9217 7219 9275 7225
rect 10229 7225 10241 7228
rect 10275 7225 10287 7259
rect 10229 7219 10287 7225
rect 12758 7259 12816 7265
rect 12758 7225 12770 7259
rect 12804 7225 12816 7259
rect 12758 7219 12816 7225
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 7248 7160 7481 7188
rect 7248 7148 7254 7160
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 9232 7188 9260 7219
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 9232 7160 10701 7188
rect 7469 7151 7527 7157
rect 10689 7157 10701 7160
rect 10735 7188 10747 7191
rect 11698 7188 11704 7200
rect 10735 7160 11704 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 12161 7191 12219 7197
rect 12161 7188 12173 7191
rect 12124 7160 12173 7188
rect 12124 7148 12130 7160
rect 12161 7157 12173 7160
rect 12207 7188 12219 7191
rect 12773 7188 12801 7219
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 19438 7265 19466 7364
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 24504 7333 24532 7432
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 32033 7463 32091 7469
rect 26384 7432 27752 7460
rect 26384 7420 26390 7432
rect 26970 7352 26976 7404
rect 27028 7392 27034 7404
rect 27433 7395 27491 7401
rect 27433 7392 27445 7395
rect 27028 7364 27445 7392
rect 27028 7352 27034 7364
rect 27433 7361 27445 7364
rect 27479 7392 27491 7395
rect 27522 7392 27528 7404
rect 27479 7364 27528 7392
rect 27479 7361 27491 7364
rect 27433 7355 27491 7361
rect 27522 7352 27528 7364
rect 27580 7352 27586 7404
rect 27724 7401 27752 7432
rect 32033 7429 32045 7463
rect 32079 7460 32091 7463
rect 33410 7460 33416 7472
rect 32079 7432 33416 7460
rect 32079 7429 32091 7432
rect 32033 7423 32091 7429
rect 33410 7420 33416 7432
rect 33468 7420 33474 7472
rect 33965 7463 34023 7469
rect 33965 7429 33977 7463
rect 34011 7460 34023 7463
rect 35897 7463 35955 7469
rect 35897 7460 35909 7463
rect 34011 7432 35909 7460
rect 34011 7429 34023 7432
rect 33965 7423 34023 7429
rect 35897 7429 35909 7432
rect 35943 7460 35955 7463
rect 36630 7460 36636 7472
rect 35943 7432 36636 7460
rect 35943 7429 35955 7432
rect 35897 7423 35955 7429
rect 36630 7420 36636 7432
rect 36688 7420 36694 7472
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 30650 7352 30656 7404
rect 30708 7392 30714 7404
rect 33778 7392 33784 7404
rect 30708 7364 33784 7392
rect 30708 7352 30714 7364
rect 33778 7352 33784 7364
rect 33836 7352 33842 7404
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7392 35035 7395
rect 35250 7392 35256 7404
rect 35023 7364 35256 7392
rect 35023 7361 35035 7364
rect 34977 7355 35035 7361
rect 35250 7352 35256 7364
rect 35308 7352 35314 7404
rect 35618 7352 35624 7404
rect 35676 7392 35682 7404
rect 36817 7395 36875 7401
rect 36817 7392 36829 7395
rect 35676 7364 36829 7392
rect 35676 7352 35682 7364
rect 36817 7361 36829 7364
rect 36863 7361 36875 7395
rect 36817 7355 36875 7361
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23952 7296 24041 7324
rect 14001 7259 14059 7265
rect 14001 7256 14013 7259
rect 12952 7228 14013 7256
rect 12952 7216 12958 7228
rect 14001 7225 14013 7228
rect 14047 7225 14059 7259
rect 14001 7219 14059 7225
rect 19423 7259 19481 7265
rect 19423 7225 19435 7259
rect 19469 7225 19481 7259
rect 19423 7219 19481 7225
rect 20806 7216 20812 7268
rect 20864 7256 20870 7268
rect 21177 7259 21235 7265
rect 21177 7256 21189 7259
rect 20864 7228 21189 7256
rect 20864 7216 20870 7228
rect 21177 7225 21189 7228
rect 21223 7225 21235 7259
rect 21177 7219 21235 7225
rect 21269 7259 21327 7265
rect 21269 7225 21281 7259
rect 21315 7225 21327 7259
rect 21818 7256 21824 7268
rect 21779 7228 21824 7256
rect 21269 7219 21327 7225
rect 13354 7188 13360 7200
rect 12207 7160 12801 7188
rect 13315 7160 13360 7188
rect 12207 7157 12219 7160
rect 12161 7151 12219 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 17368 7160 17417 7188
rect 17368 7148 17374 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 20625 7191 20683 7197
rect 20625 7157 20637 7191
rect 20671 7188 20683 7191
rect 21284 7188 21312 7219
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 23952 7200 23980 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 24489 7327 24547 7333
rect 24489 7293 24501 7327
rect 24535 7293 24547 7327
rect 24489 7287 24547 7293
rect 25133 7327 25191 7333
rect 25133 7293 25145 7327
rect 25179 7324 25191 7327
rect 25593 7327 25651 7333
rect 25593 7324 25605 7327
rect 25179 7296 25605 7324
rect 25179 7293 25191 7296
rect 25133 7287 25191 7293
rect 25593 7293 25605 7296
rect 25639 7324 25651 7327
rect 26602 7324 26608 7336
rect 25639 7296 26608 7324
rect 25639 7293 25651 7296
rect 25593 7287 25651 7293
rect 26602 7284 26608 7296
rect 26660 7284 26666 7336
rect 29086 7284 29092 7336
rect 29144 7324 29150 7336
rect 29273 7327 29331 7333
rect 29273 7324 29285 7327
rect 29144 7296 29285 7324
rect 29144 7284 29150 7296
rect 29273 7293 29285 7296
rect 29319 7293 29331 7327
rect 29730 7324 29736 7336
rect 29691 7296 29736 7324
rect 29273 7287 29331 7293
rect 29730 7284 29736 7296
rect 29788 7284 29794 7336
rect 31110 7324 31116 7336
rect 31071 7296 31116 7324
rect 31110 7284 31116 7296
rect 31168 7284 31174 7336
rect 32858 7284 32864 7336
rect 32916 7324 32922 7336
rect 33045 7327 33103 7333
rect 33045 7324 33057 7327
rect 32916 7296 33057 7324
rect 32916 7284 32922 7296
rect 33045 7293 33057 7296
rect 33091 7324 33103 7327
rect 34241 7327 34299 7333
rect 34241 7324 34253 7327
rect 33091 7296 34253 7324
rect 33091 7293 33103 7296
rect 33045 7287 33103 7293
rect 34241 7293 34253 7296
rect 34287 7293 34299 7327
rect 34241 7287 34299 7293
rect 25914 7259 25972 7265
rect 25914 7256 25926 7259
rect 25608 7228 25926 7256
rect 25608 7200 25636 7228
rect 25914 7225 25926 7228
rect 25960 7225 25972 7259
rect 27525 7259 27583 7265
rect 27525 7256 27537 7259
rect 25914 7219 25972 7225
rect 27172 7228 27537 7256
rect 27172 7200 27200 7228
rect 27525 7225 27537 7228
rect 27571 7225 27583 7259
rect 27525 7219 27583 7225
rect 31021 7259 31079 7265
rect 31021 7225 31033 7259
rect 31067 7256 31079 7259
rect 31475 7259 31533 7265
rect 31475 7256 31487 7259
rect 31067 7228 31487 7256
rect 31067 7225 31079 7228
rect 31021 7219 31079 7225
rect 31475 7225 31487 7228
rect 31521 7256 31533 7259
rect 35069 7259 35127 7265
rect 31521 7228 32628 7256
rect 31521 7225 31533 7228
rect 31475 7219 31533 7225
rect 21726 7188 21732 7200
rect 20671 7160 21732 7188
rect 20671 7157 20683 7160
rect 20625 7151 20683 7157
rect 21726 7148 21732 7160
rect 21784 7148 21790 7200
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22097 7191 22155 7197
rect 22097 7188 22109 7191
rect 22060 7160 22109 7188
rect 22060 7148 22066 7160
rect 22097 7157 22109 7160
rect 22143 7157 22155 7191
rect 23934 7188 23940 7200
rect 23895 7160 23940 7188
rect 22097 7151 22155 7157
rect 23934 7148 23940 7160
rect 23992 7148 23998 7200
rect 24118 7188 24124 7200
rect 24079 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 25501 7191 25559 7197
rect 25501 7157 25513 7191
rect 25547 7188 25559 7191
rect 25590 7188 25596 7200
rect 25547 7160 25596 7188
rect 25547 7157 25559 7160
rect 25501 7151 25559 7157
rect 25590 7148 25596 7160
rect 25648 7148 25654 7200
rect 26513 7191 26571 7197
rect 26513 7157 26525 7191
rect 26559 7188 26571 7191
rect 26694 7188 26700 7200
rect 26559 7160 26700 7188
rect 26559 7157 26571 7160
rect 26513 7151 26571 7157
rect 26694 7148 26700 7160
rect 26752 7148 26758 7200
rect 27154 7188 27160 7200
rect 27115 7160 27160 7188
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 27430 7148 27436 7200
rect 27488 7188 27494 7200
rect 28629 7191 28687 7197
rect 28629 7188 28641 7191
rect 27488 7160 28641 7188
rect 27488 7148 27494 7160
rect 28629 7157 28641 7160
rect 28675 7188 28687 7191
rect 28902 7188 28908 7200
rect 28675 7160 28908 7188
rect 28675 7157 28687 7160
rect 28629 7151 28687 7157
rect 28902 7148 28908 7160
rect 28960 7148 28966 7200
rect 29546 7188 29552 7200
rect 29507 7160 29552 7188
rect 29546 7148 29552 7160
rect 29604 7148 29610 7200
rect 32600 7197 32628 7228
rect 35069 7225 35081 7259
rect 35115 7225 35127 7259
rect 35069 7219 35127 7225
rect 35621 7259 35679 7265
rect 35621 7225 35633 7259
rect 35667 7256 35679 7259
rect 35710 7256 35716 7268
rect 35667 7228 35716 7256
rect 35667 7225 35679 7228
rect 35621 7219 35679 7225
rect 32585 7191 32643 7197
rect 32585 7157 32597 7191
rect 32631 7188 32643 7191
rect 32953 7191 33011 7197
rect 32953 7188 32965 7191
rect 32631 7160 32965 7188
rect 32631 7157 32643 7160
rect 32585 7151 32643 7157
rect 32953 7157 32965 7160
rect 32999 7188 33011 7191
rect 33318 7188 33324 7200
rect 32999 7160 33324 7188
rect 32999 7157 33011 7160
rect 32953 7151 33011 7157
rect 33318 7148 33324 7160
rect 33376 7188 33382 7200
rect 33413 7191 33471 7197
rect 33413 7188 33425 7191
rect 33376 7160 33425 7188
rect 33376 7148 33382 7160
rect 33413 7157 33425 7160
rect 33459 7188 33471 7191
rect 34054 7188 34060 7200
rect 33459 7160 34060 7188
rect 33459 7157 33471 7160
rect 33413 7151 33471 7157
rect 34054 7148 34060 7160
rect 34112 7148 34118 7200
rect 34517 7191 34575 7197
rect 34517 7157 34529 7191
rect 34563 7188 34575 7191
rect 34606 7188 34612 7200
rect 34563 7160 34612 7188
rect 34563 7157 34575 7160
rect 34517 7151 34575 7157
rect 34606 7148 34612 7160
rect 34664 7188 34670 7200
rect 35084 7188 35112 7219
rect 35710 7216 35716 7228
rect 35768 7216 35774 7268
rect 36354 7216 36360 7268
rect 36412 7256 36418 7268
rect 36541 7259 36599 7265
rect 36541 7256 36553 7259
rect 36412 7228 36553 7256
rect 36412 7216 36418 7228
rect 36541 7225 36553 7228
rect 36587 7225 36599 7259
rect 36541 7219 36599 7225
rect 36630 7216 36636 7268
rect 36688 7256 36694 7268
rect 36688 7228 36733 7256
rect 36688 7216 36694 7228
rect 36262 7188 36268 7200
rect 34664 7160 35112 7188
rect 36223 7160 36268 7188
rect 34664 7148 34670 7160
rect 36262 7148 36268 7160
rect 36320 7148 36326 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1854 6984 1860 6996
rect 1815 6956 1860 6984
rect 1854 6944 1860 6956
rect 1912 6944 1918 6996
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 4154 6984 4160 6996
rect 3844 6956 4160 6984
rect 3844 6944 3850 6956
rect 4154 6944 4160 6956
rect 4212 6984 4218 6996
rect 4430 6984 4436 6996
rect 4212 6956 4436 6984
rect 4212 6944 4218 6956
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 7650 6984 7656 6996
rect 6236 6956 7656 6984
rect 6236 6944 6242 6956
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 9490 6944 9496 6996
rect 9548 6984 9554 6996
rect 10134 6984 10140 6996
rect 9548 6956 10140 6984
rect 9548 6944 9554 6956
rect 10134 6944 10140 6956
rect 10192 6984 10198 6996
rect 14231 6987 14289 6993
rect 14231 6984 14243 6987
rect 10192 6956 14243 6984
rect 10192 6944 10198 6956
rect 14231 6953 14243 6956
rect 14277 6953 14289 6987
rect 14231 6947 14289 6953
rect 15933 6987 15991 6993
rect 15933 6953 15945 6987
rect 15979 6984 15991 6987
rect 16850 6984 16856 6996
rect 15979 6956 16856 6984
rect 15979 6953 15991 6956
rect 15933 6947 15991 6953
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 19935 6987 19993 6993
rect 19935 6953 19947 6987
rect 19981 6984 19993 6987
rect 20346 6984 20352 6996
rect 19981 6956 20352 6984
rect 19981 6953 19993 6956
rect 19935 6947 19993 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 21266 6984 21272 6996
rect 21227 6956 21272 6984
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 21726 6944 21732 6996
rect 21784 6984 21790 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 21784 6956 21833 6984
rect 21784 6944 21790 6956
rect 21821 6953 21833 6956
rect 21867 6953 21879 6987
rect 22738 6984 22744 6996
rect 22699 6956 22744 6984
rect 21821 6947 21879 6953
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 24394 6984 24400 6996
rect 24355 6956 24400 6984
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 26237 6987 26295 6993
rect 26237 6984 26249 6987
rect 24872 6956 26249 6984
rect 2498 6876 2504 6928
rect 2556 6916 2562 6928
rect 2593 6919 2651 6925
rect 2593 6916 2605 6919
rect 2556 6888 2605 6916
rect 2556 6876 2562 6888
rect 2593 6885 2605 6888
rect 2639 6916 2651 6919
rect 4246 6916 4252 6928
rect 2639 6888 4252 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 4246 6876 4252 6888
rect 4304 6916 4310 6928
rect 4890 6916 4896 6928
rect 4304 6888 4896 6916
rect 4304 6876 4310 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 6914 6876 6920 6928
rect 6972 6916 6978 6928
rect 7377 6919 7435 6925
rect 7377 6916 7389 6919
rect 6972 6888 7389 6916
rect 6972 6876 6978 6888
rect 7377 6885 7389 6888
rect 7423 6916 7435 6919
rect 8754 6916 8760 6928
rect 7423 6888 8760 6916
rect 7423 6885 7435 6888
rect 7377 6879 7435 6885
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 10870 6916 10876 6928
rect 10831 6888 10876 6916
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 11701 6919 11759 6925
rect 11701 6916 11713 6919
rect 11664 6888 11713 6916
rect 11664 6876 11670 6888
rect 11701 6885 11713 6888
rect 11747 6885 11759 6919
rect 11701 6879 11759 6885
rect 12066 6876 12072 6928
rect 12124 6916 12130 6928
rect 12666 6919 12724 6925
rect 12666 6916 12678 6919
rect 12124 6888 12678 6916
rect 12124 6876 12130 6888
rect 12666 6885 12678 6888
rect 12712 6885 12724 6919
rect 12666 6879 12724 6885
rect 16022 6876 16028 6928
rect 16080 6916 16086 6928
rect 16438 6919 16496 6925
rect 16438 6916 16450 6919
rect 16080 6888 16450 6916
rect 16080 6876 16086 6888
rect 16438 6885 16450 6888
rect 16484 6885 16496 6919
rect 16868 6916 16896 6944
rect 18601 6919 18659 6925
rect 16868 6888 18368 6916
rect 16438 6879 16496 6885
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 6144 6820 6193 6848
rect 6144 6808 6150 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 6181 6811 6239 6817
rect 7116 6820 7757 6848
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 3602 6780 3608 6792
rect 2547 6752 3608 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4430 6780 4436 6792
rect 4212 6752 4257 6780
rect 4391 6752 4436 6780
rect 4212 6740 4218 6752
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6362 6780 6368 6792
rect 6043 6752 6368 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 7116 6780 7144 6820
rect 7745 6817 7757 6820
rect 7791 6848 7803 6851
rect 8018 6848 8024 6860
rect 7791 6820 8024 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 8018 6808 8024 6820
rect 8076 6848 8082 6860
rect 9950 6848 9956 6860
rect 8076 6820 9628 6848
rect 9911 6820 9956 6848
rect 8076 6808 8082 6820
rect 8110 6780 8116 6792
rect 6420 6752 7144 6780
rect 7208 6752 8116 6780
rect 6420 6740 6426 6752
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3970 6712 3976 6724
rect 3099 6684 3976 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3970 6672 3976 6684
rect 4028 6712 4034 6724
rect 4798 6712 4804 6724
rect 4028 6684 4804 6712
rect 4028 6672 4034 6684
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1762 6644 1768 6656
rect 1627 6616 1768 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1762 6604 1768 6616
rect 1820 6604 1826 6656
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2740 6616 3433 6644
rect 2740 6604 2746 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3421 6607 3479 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7006 6644 7012 6656
rect 6963 6616 7012 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7006 6604 7012 6616
rect 7064 6644 7070 6656
rect 7208 6653 7236 6752
rect 8110 6740 8116 6752
rect 8168 6780 8174 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8168 6752 9229 6780
rect 8168 6740 8174 6752
rect 9217 6749 9229 6752
rect 9263 6780 9275 6783
rect 9398 6780 9404 6792
rect 9263 6752 9404 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9600 6780 9628 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 11238 6848 11244 6860
rect 11199 6820 11244 6848
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 14160 6851 14218 6857
rect 14160 6817 14172 6851
rect 14206 6848 14218 6851
rect 14274 6848 14280 6860
rect 14206 6820 14280 6848
rect 14206 6817 14218 6820
rect 14160 6811 14218 6817
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 17678 6848 17684 6860
rect 14332 6820 17684 6848
rect 14332 6808 14338 6820
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 17862 6848 17868 6860
rect 17823 6820 17868 6848
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 18340 6857 18368 6888
rect 18601 6885 18613 6919
rect 18647 6916 18659 6919
rect 18690 6916 18696 6928
rect 18647 6888 18696 6916
rect 18647 6885 18659 6888
rect 18601 6879 18659 6885
rect 18690 6876 18696 6888
rect 18748 6916 18754 6928
rect 18877 6919 18935 6925
rect 18877 6916 18889 6919
rect 18748 6888 18889 6916
rect 18748 6876 18754 6888
rect 18877 6885 18889 6888
rect 18923 6885 18935 6919
rect 18877 6879 18935 6885
rect 21358 6876 21364 6928
rect 21416 6916 21422 6928
rect 24872 6916 24900 6956
rect 26237 6953 26249 6956
rect 26283 6984 26295 6987
rect 26326 6984 26332 6996
rect 26283 6956 26332 6984
rect 26283 6953 26295 6956
rect 26237 6947 26295 6953
rect 26326 6944 26332 6956
rect 26384 6944 26390 6996
rect 27522 6984 27528 6996
rect 27483 6956 27528 6984
rect 27522 6944 27528 6956
rect 27580 6944 27586 6996
rect 31110 6944 31116 6996
rect 31168 6984 31174 6996
rect 31481 6987 31539 6993
rect 31481 6984 31493 6987
rect 31168 6956 31493 6984
rect 31168 6944 31174 6956
rect 31481 6953 31493 6956
rect 31527 6984 31539 6987
rect 32217 6987 32275 6993
rect 32217 6984 32229 6987
rect 31527 6956 32229 6984
rect 31527 6953 31539 6956
rect 31481 6947 31539 6953
rect 32217 6953 32229 6956
rect 32263 6953 32275 6987
rect 32217 6947 32275 6953
rect 33229 6987 33287 6993
rect 33229 6953 33241 6987
rect 33275 6984 33287 6987
rect 33410 6984 33416 6996
rect 33275 6956 33416 6984
rect 33275 6953 33287 6956
rect 33229 6947 33287 6953
rect 33410 6944 33416 6956
rect 33468 6944 33474 6996
rect 34054 6984 34060 6996
rect 34015 6956 34060 6984
rect 34054 6944 34060 6956
rect 34112 6944 34118 6996
rect 34977 6987 35035 6993
rect 34977 6953 34989 6987
rect 35023 6984 35035 6987
rect 35066 6984 35072 6996
rect 35023 6956 35072 6984
rect 35023 6953 35035 6956
rect 34977 6947 35035 6953
rect 35066 6944 35072 6956
rect 35124 6984 35130 6996
rect 36357 6987 36415 6993
rect 36357 6984 36369 6987
rect 35124 6956 36369 6984
rect 35124 6944 35130 6956
rect 36357 6953 36369 6956
rect 36403 6953 36415 6987
rect 36357 6947 36415 6953
rect 25038 6916 25044 6928
rect 21416 6888 24900 6916
rect 24999 6888 25044 6916
rect 21416 6876 21422 6888
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 26694 6916 26700 6928
rect 26655 6888 26700 6916
rect 26694 6876 26700 6888
rect 26752 6876 26758 6928
rect 27246 6916 27252 6928
rect 27207 6888 27252 6916
rect 27246 6876 27252 6888
rect 27304 6876 27310 6928
rect 30098 6916 30104 6928
rect 28828 6888 30104 6916
rect 18325 6851 18383 6857
rect 18325 6817 18337 6851
rect 18371 6817 18383 6851
rect 19794 6848 19800 6860
rect 19755 6820 19800 6848
rect 18325 6811 18383 6817
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 22830 6848 22836 6860
rect 20548 6820 22836 6848
rect 11790 6780 11796 6792
rect 9600 6752 11796 6780
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 12345 6783 12403 6789
rect 12345 6749 12357 6783
rect 12391 6780 12403 6783
rect 12986 6780 12992 6792
rect 12391 6752 12992 6780
rect 12391 6749 12403 6752
rect 12345 6743 12403 6749
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16298 6780 16304 6792
rect 16163 6752 16304 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 17880 6780 17908 6808
rect 20548 6780 20576 6820
rect 22830 6808 22836 6820
rect 22888 6808 22894 6860
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6817 23167 6851
rect 23109 6811 23167 6817
rect 17880 6752 20576 6780
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20680 6752 20913 6780
rect 20680 6740 20686 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 23124 6780 23152 6811
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 28828 6857 28856 6888
rect 30098 6876 30104 6888
rect 30156 6876 30162 6928
rect 30837 6919 30895 6925
rect 30837 6885 30849 6919
rect 30883 6916 30895 6919
rect 33870 6916 33876 6928
rect 30883 6888 33876 6916
rect 30883 6885 30895 6888
rect 30837 6879 30895 6885
rect 33870 6876 33876 6888
rect 33928 6876 33934 6928
rect 35799 6919 35857 6925
rect 35799 6885 35811 6919
rect 35845 6916 35857 6919
rect 35894 6916 35900 6928
rect 35845 6888 35900 6916
rect 35845 6885 35857 6888
rect 35799 6879 35857 6885
rect 35894 6876 35900 6888
rect 35952 6876 35958 6928
rect 28813 6851 28871 6857
rect 28813 6848 28825 6851
rect 28684 6820 28825 6848
rect 28684 6808 28690 6820
rect 28813 6817 28825 6820
rect 28859 6817 28871 6851
rect 28994 6848 29000 6860
rect 28955 6820 29000 6848
rect 28813 6811 28871 6817
rect 28994 6808 29000 6820
rect 29052 6848 29058 6860
rect 29549 6851 29607 6857
rect 29549 6848 29561 6851
rect 29052 6820 29561 6848
rect 29052 6808 29058 6820
rect 29549 6817 29561 6820
rect 29595 6848 29607 6851
rect 29730 6848 29736 6860
rect 29595 6820 29736 6848
rect 29595 6817 29607 6820
rect 29549 6811 29607 6817
rect 29730 6808 29736 6820
rect 29788 6808 29794 6860
rect 29825 6851 29883 6857
rect 29825 6817 29837 6851
rect 29871 6848 29883 6851
rect 30374 6848 30380 6860
rect 29871 6820 30380 6848
rect 29871 6817 29883 6820
rect 29825 6811 29883 6817
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 30653 6851 30711 6857
rect 30653 6817 30665 6851
rect 30699 6848 30711 6851
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 30699 6820 30880 6848
rect 30699 6817 30711 6820
rect 30653 6811 30711 6817
rect 30852 6792 30880 6820
rect 31220 6820 32137 6848
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 22428 6752 24041 6780
rect 22428 6740 22434 6752
rect 24029 6749 24041 6752
rect 24075 6780 24087 6783
rect 24118 6780 24124 6792
rect 24075 6752 24124 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24946 6780 24952 6792
rect 24907 6752 24952 6780
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 25593 6783 25651 6789
rect 25593 6749 25605 6783
rect 25639 6780 25651 6783
rect 26605 6783 26663 6789
rect 26605 6780 26617 6783
rect 25639 6752 26617 6780
rect 25639 6749 25651 6752
rect 25593 6743 25651 6749
rect 26605 6749 26617 6752
rect 26651 6780 26663 6783
rect 28166 6780 28172 6792
rect 26651 6752 28172 6780
rect 26651 6749 26663 6752
rect 26605 6743 26663 6749
rect 7377 6715 7435 6721
rect 7377 6681 7389 6715
rect 7423 6712 7435 6715
rect 7910 6715 7968 6721
rect 7423 6684 7834 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 7064 6616 7205 6644
rect 7064 6604 7070 6616
rect 7193 6613 7205 6616
rect 7239 6613 7251 6647
rect 7193 6607 7251 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7524 6616 7573 6644
rect 7524 6604 7530 6616
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7806 6644 7834 6684
rect 7910 6681 7922 6715
rect 7956 6712 7968 6715
rect 8662 6712 8668 6724
rect 7956 6684 8668 6712
rect 7956 6681 7968 6684
rect 7910 6675 7968 6681
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 25608 6712 25636 6743
rect 28166 6740 28172 6752
rect 28224 6740 28230 6792
rect 29270 6780 29276 6792
rect 29231 6752 29276 6780
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 30834 6740 30840 6792
rect 30892 6780 30898 6792
rect 31113 6783 31171 6789
rect 31113 6780 31125 6783
rect 30892 6752 31125 6780
rect 30892 6740 30898 6752
rect 31113 6749 31125 6752
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 21876 6684 25636 6712
rect 21876 6672 21882 6684
rect 28902 6672 28908 6724
rect 28960 6712 28966 6724
rect 31220 6712 31248 6820
rect 32125 6817 32137 6820
rect 32171 6848 32183 6851
rect 32398 6848 32404 6860
rect 32171 6820 32404 6848
rect 32171 6817 32183 6820
rect 32125 6811 32183 6817
rect 32398 6808 32404 6820
rect 32456 6808 32462 6860
rect 32582 6848 32588 6860
rect 32543 6820 32588 6848
rect 32582 6808 32588 6820
rect 32640 6808 32646 6860
rect 34698 6808 34704 6860
rect 34756 6848 34762 6860
rect 36354 6848 36360 6860
rect 34756 6820 36360 6848
rect 34756 6808 34762 6820
rect 36354 6808 36360 6820
rect 36412 6848 36418 6860
rect 36633 6851 36691 6857
rect 36633 6848 36645 6851
rect 36412 6820 36645 6848
rect 36412 6808 36418 6820
rect 36633 6817 36645 6820
rect 36679 6817 36691 6851
rect 36633 6811 36691 6817
rect 33594 6740 33600 6792
rect 33652 6780 33658 6792
rect 33689 6783 33747 6789
rect 33689 6780 33701 6783
rect 33652 6752 33701 6780
rect 33652 6740 33658 6752
rect 33689 6749 33701 6752
rect 33735 6749 33747 6783
rect 35434 6780 35440 6792
rect 35395 6752 35440 6780
rect 33689 6743 33747 6749
rect 35434 6740 35440 6752
rect 35492 6740 35498 6792
rect 33505 6715 33563 6721
rect 33505 6712 33517 6715
rect 28960 6684 31248 6712
rect 33106 6684 33517 6712
rect 28960 6672 28966 6684
rect 33106 6656 33134 6684
rect 33505 6681 33517 6684
rect 33551 6681 33563 6715
rect 33505 6675 33563 6681
rect 34609 6715 34667 6721
rect 34609 6681 34621 6715
rect 34655 6712 34667 6715
rect 35066 6712 35072 6724
rect 34655 6684 35072 6712
rect 34655 6681 34667 6684
rect 34609 6675 34667 6681
rect 35066 6672 35072 6684
rect 35124 6712 35130 6724
rect 35253 6715 35311 6721
rect 35253 6712 35265 6715
rect 35124 6684 35265 6712
rect 35124 6672 35130 6684
rect 35253 6681 35265 6684
rect 35299 6681 35311 6715
rect 35253 6675 35311 6681
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 7806 6616 8033 6644
rect 7561 6607 7619 6613
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8021 6607 8079 6613
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 10134 6644 10140 6656
rect 10095 6616 10140 6644
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11379 6647 11437 6653
rect 11379 6644 11391 6647
rect 11204 6616 11391 6644
rect 11204 6604 11210 6616
rect 11379 6613 11391 6616
rect 11425 6613 11437 6647
rect 12158 6644 12164 6656
rect 12119 6616 12164 6644
rect 11379 6607 11437 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 13262 6644 13268 6656
rect 13223 6616 13268 6644
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 15102 6644 15108 6656
rect 14783 6616 15108 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 15102 6604 15108 6616
rect 15160 6644 15166 6656
rect 15470 6644 15476 6656
rect 15160 6616 15476 6644
rect 15160 6604 15166 6616
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16632 6616 17049 6644
rect 16632 6604 16638 6616
rect 17037 6613 17049 6616
rect 17083 6644 17095 6647
rect 18230 6644 18236 6656
rect 17083 6616 18236 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 18782 6604 18788 6656
rect 18840 6644 18846 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 18840 6616 19257 6644
rect 18840 6604 18846 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19245 6607 19303 6613
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20588 6616 20637 6644
rect 20588 6604 20594 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 22097 6647 22155 6653
rect 22097 6644 22109 6647
rect 20864 6616 22109 6644
rect 20864 6604 20870 6616
rect 22097 6613 22109 6616
rect 22143 6613 22155 6647
rect 22097 6607 22155 6613
rect 23753 6647 23811 6653
rect 23753 6613 23765 6647
rect 23799 6644 23811 6647
rect 23842 6644 23848 6656
rect 23799 6616 23848 6644
rect 23799 6613 23811 6616
rect 23753 6607 23811 6613
rect 23842 6604 23848 6616
rect 23900 6644 23906 6656
rect 25314 6644 25320 6656
rect 23900 6616 25320 6644
rect 23900 6604 23906 6616
rect 25314 6604 25320 6616
rect 25372 6644 25378 6656
rect 29825 6647 29883 6653
rect 29825 6644 29837 6647
rect 25372 6616 29837 6644
rect 25372 6604 25378 6616
rect 29825 6613 29837 6616
rect 29871 6613 29883 6647
rect 30006 6644 30012 6656
rect 29967 6616 30012 6644
rect 29825 6607 29883 6613
rect 30006 6604 30012 6616
rect 30064 6604 30070 6656
rect 31386 6604 31392 6656
rect 31444 6644 31450 6656
rect 33042 6644 33048 6656
rect 31444 6616 33048 6644
rect 31444 6604 31450 6616
rect 33042 6604 33048 6616
rect 33100 6616 33134 6656
rect 33100 6604 33106 6616
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 3200 6412 3617 6440
rect 3200 6400 3206 6412
rect 3605 6409 3617 6412
rect 3651 6440 3663 6443
rect 4338 6440 4344 6452
rect 3651 6412 4344 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5626 6440 5632 6452
rect 5587 6412 5632 6440
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 7929 6443 7987 6449
rect 5828 6412 7696 6440
rect 4065 6375 4123 6381
rect 4065 6341 4077 6375
rect 4111 6372 4123 6375
rect 4246 6372 4252 6384
rect 4111 6344 4252 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 4246 6332 4252 6344
rect 4304 6332 4310 6384
rect 4798 6372 4804 6384
rect 4711 6344 4804 6372
rect 4798 6332 4804 6344
rect 4856 6372 4862 6384
rect 5828 6372 5856 6412
rect 4856 6344 5856 6372
rect 5905 6375 5963 6381
rect 4856 6332 4862 6344
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 7006 6372 7012 6384
rect 5951 6344 7012 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7668 6372 7696 6412
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 8018 6440 8024 6452
rect 7975 6412 8024 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 12124 6412 12173 6440
rect 12124 6400 12130 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13412 6412 13645 6440
rect 13412 6400 13418 6412
rect 13633 6409 13645 6412
rect 13679 6440 13691 6443
rect 14366 6440 14372 6452
rect 13679 6412 14372 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 15565 6443 15623 6449
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 15930 6440 15936 6452
rect 15611 6412 15936 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 10318 6372 10324 6384
rect 7668 6344 10324 6372
rect 10318 6332 10324 6344
rect 10376 6332 10382 6384
rect 15580 6372 15608 6403
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 16908 6412 17417 6440
rect 16908 6400 16914 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 19935 6443 19993 6449
rect 19935 6409 19947 6443
rect 19981 6440 19993 6443
rect 20806 6440 20812 6452
rect 19981 6412 20812 6440
rect 19981 6409 19993 6412
rect 19935 6403 19993 6409
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21726 6400 21732 6452
rect 21784 6440 21790 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21784 6412 21833 6440
rect 21784 6400 21790 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 24949 6443 25007 6449
rect 24949 6409 24961 6443
rect 24995 6440 25007 6443
rect 25038 6440 25044 6452
rect 24995 6412 25044 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 25038 6400 25044 6412
rect 25096 6440 25102 6452
rect 26329 6443 26387 6449
rect 26329 6440 26341 6443
rect 25096 6412 26341 6440
rect 25096 6400 25102 6412
rect 26329 6409 26341 6412
rect 26375 6440 26387 6443
rect 27154 6440 27160 6452
rect 26375 6412 27160 6440
rect 26375 6409 26387 6412
rect 26329 6403 26387 6409
rect 27154 6400 27160 6412
rect 27212 6400 27218 6452
rect 28166 6440 28172 6452
rect 28127 6412 28172 6440
rect 28166 6400 28172 6412
rect 28224 6400 28230 6452
rect 28626 6440 28632 6452
rect 28587 6412 28632 6440
rect 28626 6400 28632 6412
rect 28684 6400 28690 6452
rect 29733 6443 29791 6449
rect 29733 6409 29745 6443
rect 29779 6440 29791 6443
rect 30834 6440 30840 6452
rect 29779 6412 30840 6440
rect 29779 6409 29791 6412
rect 29733 6403 29791 6409
rect 30834 6400 30840 6412
rect 30892 6400 30898 6452
rect 32493 6443 32551 6449
rect 32493 6409 32505 6443
rect 32539 6440 32551 6443
rect 32582 6440 32588 6452
rect 32539 6412 32588 6440
rect 32539 6409 32551 6412
rect 32493 6403 32551 6409
rect 32582 6400 32588 6412
rect 32640 6400 32646 6452
rect 34054 6400 34060 6452
rect 34112 6440 34118 6452
rect 34241 6443 34299 6449
rect 34241 6440 34253 6443
rect 34112 6412 34253 6440
rect 34112 6400 34118 6412
rect 34241 6409 34253 6412
rect 34287 6440 34299 6443
rect 35894 6440 35900 6452
rect 34287 6412 35900 6440
rect 34287 6409 34299 6412
rect 34241 6403 34299 6409
rect 35894 6400 35900 6412
rect 35952 6400 35958 6452
rect 36630 6440 36636 6452
rect 36591 6412 36636 6440
rect 36630 6400 36636 6412
rect 36688 6400 36694 6452
rect 37090 6440 37096 6452
rect 37051 6412 37096 6440
rect 37090 6400 37096 6412
rect 37148 6400 37154 6452
rect 13786 6344 15608 6372
rect 2682 6304 2688 6316
rect 2643 6276 2688 6304
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6304 3387 6307
rect 3786 6304 3792 6316
rect 3375 6276 3792 6304
rect 3375 6273 3387 6276
rect 3329 6267 3387 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 7190 6304 7196 6316
rect 6687 6276 7196 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2038 6236 2044 6248
rect 1443 6208 2044 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 6840 6245 6868 6276
rect 7190 6264 7196 6276
rect 7248 6304 7254 6316
rect 10045 6307 10103 6313
rect 7248 6276 8248 6304
rect 7248 6264 7254 6276
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5184 6208 5733 6236
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 3142 6168 3148 6180
rect 2823 6140 3148 6168
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 4246 6168 4252 6180
rect 4207 6140 4252 6168
rect 4246 6128 4252 6140
rect 4304 6128 4310 6180
rect 4338 6128 4344 6180
rect 4396 6168 4402 6180
rect 4396 6140 4441 6168
rect 4396 6128 4402 6140
rect 5184 6112 5212 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7098 6236 7104 6248
rect 6972 6208 7017 6236
rect 7059 6208 7104 6236
rect 6972 6196 6978 6208
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8220 6236 8248 6276
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 11146 6304 11152 6316
rect 10091 6276 11152 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 11296 6276 11341 6304
rect 11296 6264 11302 6276
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 8220 6208 8493 6236
rect 8220 6112 8248 6208
rect 8481 6205 8493 6208
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11931 6208 12449 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 12437 6205 12449 6208
rect 12483 6236 12495 6239
rect 13354 6236 13360 6248
rect 12483 6208 13360 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 10137 6171 10195 6177
rect 10137 6137 10149 6171
rect 10183 6137 10195 6171
rect 10137 6131 10195 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 10778 6168 10784 6180
rect 10735 6140 10784 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 6144 6072 6193 6100
rect 6144 6060 6150 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 7282 6100 7288 6112
rect 7243 6072 7288 6100
rect 6181 6063 6239 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 8202 6100 8208 6112
rect 8163 6072 8208 6100
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9861 6103 9919 6109
rect 9861 6069 9873 6103
rect 9907 6100 9919 6103
rect 9950 6100 9956 6112
rect 9907 6072 9956 6100
rect 9907 6069 9919 6072
rect 9861 6063 9919 6069
rect 9950 6060 9956 6072
rect 10008 6100 10014 6112
rect 10152 6100 10180 6131
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 12758 6171 12816 6177
rect 12758 6168 12770 6171
rect 12124 6140 12770 6168
rect 12124 6128 12130 6140
rect 12758 6137 12770 6140
rect 12804 6168 12816 6171
rect 13786 6168 13814 6344
rect 19242 6332 19248 6384
rect 19300 6372 19306 6384
rect 19300 6344 23474 6372
rect 19300 6332 19306 6344
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14274 6304 14280 6316
rect 14139 6276 14280 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 17773 6307 17831 6313
rect 17773 6304 17785 6307
rect 15804 6276 17785 6304
rect 15804 6264 15810 6276
rect 17773 6273 17785 6276
rect 17819 6304 17831 6307
rect 17862 6304 17868 6316
rect 17819 6276 17868 6304
rect 17819 6273 17831 6276
rect 17773 6267 17831 6273
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 18414 6304 18420 6316
rect 18375 6276 18420 6304
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 19879 6276 20361 6304
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6236 16083 6239
rect 16666 6236 16672 6248
rect 16071 6208 16672 6236
rect 16071 6205 16083 6208
rect 16025 6199 16083 6205
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 19879 6245 19907 6276
rect 20349 6273 20361 6276
rect 20395 6304 20407 6307
rect 21266 6304 21272 6316
rect 20395 6276 21272 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 21416 6276 21461 6304
rect 21416 6264 21422 6276
rect 19864 6239 19922 6245
rect 19864 6205 19876 6239
rect 19910 6205 19922 6239
rect 19864 6199 19922 6205
rect 22624 6239 22682 6245
rect 22624 6205 22636 6239
rect 22670 6236 22682 6239
rect 23014 6236 23020 6248
rect 22670 6208 23020 6236
rect 22670 6205 22682 6208
rect 22624 6199 22682 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 23446 6236 23474 6344
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 26881 6375 26939 6381
rect 26881 6372 26893 6375
rect 23624 6344 26893 6372
rect 23624 6332 23630 6344
rect 26881 6341 26893 6344
rect 26927 6372 26939 6375
rect 26973 6375 27031 6381
rect 26973 6372 26985 6375
rect 26927 6344 26985 6372
rect 26927 6341 26939 6344
rect 26881 6335 26939 6341
rect 26973 6341 26985 6344
rect 27019 6341 27031 6375
rect 26973 6335 27031 6341
rect 32398 6332 32404 6384
rect 32456 6372 32462 6384
rect 32769 6375 32827 6381
rect 32769 6372 32781 6375
rect 32456 6344 32781 6372
rect 32456 6332 32462 6344
rect 32769 6341 32781 6344
rect 32815 6341 32827 6375
rect 35526 6372 35532 6384
rect 35487 6344 35532 6372
rect 32769 6335 32827 6341
rect 35526 6332 35532 6344
rect 35584 6332 35590 6384
rect 26605 6307 26663 6313
rect 26605 6304 26617 6307
rect 24136 6276 26617 6304
rect 24136 6248 24164 6276
rect 26605 6273 26617 6276
rect 26651 6304 26663 6307
rect 28905 6307 28963 6313
rect 28905 6304 28917 6307
rect 26651 6276 28917 6304
rect 26651 6273 26663 6276
rect 26605 6267 26663 6273
rect 23842 6236 23848 6248
rect 23446 6208 23848 6236
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24118 6236 24124 6248
rect 24079 6208 24124 6236
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 25409 6239 25467 6245
rect 25409 6205 25421 6239
rect 25455 6236 25467 6239
rect 25498 6236 25504 6248
rect 25455 6208 25504 6236
rect 25455 6205 25467 6208
rect 25409 6199 25467 6205
rect 25498 6196 25504 6208
rect 25556 6196 25562 6248
rect 26881 6239 26939 6245
rect 26881 6205 26893 6239
rect 26927 6236 26939 6239
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 26927 6208 27169 6236
rect 26927 6205 26939 6208
rect 26881 6199 26939 6205
rect 27157 6205 27169 6208
rect 27203 6236 27215 6239
rect 27430 6236 27436 6248
rect 27203 6208 27436 6236
rect 27203 6205 27215 6208
rect 27157 6199 27215 6205
rect 27430 6196 27436 6208
rect 27488 6196 27494 6248
rect 27632 6245 27660 6276
rect 28905 6273 28917 6276
rect 28951 6304 28963 6307
rect 28994 6304 29000 6316
rect 28951 6276 29000 6304
rect 28951 6273 28963 6276
rect 28905 6267 28963 6273
rect 28994 6264 29000 6276
rect 29052 6304 29058 6316
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 29052 6276 31217 6304
rect 29052 6264 29058 6276
rect 31205 6273 31217 6276
rect 31251 6304 31263 6307
rect 33226 6304 33232 6316
rect 31251 6276 31892 6304
rect 33187 6276 33232 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 27617 6239 27675 6245
rect 27617 6205 27629 6239
rect 27663 6205 27675 6239
rect 31478 6236 31484 6248
rect 31439 6208 31484 6236
rect 27617 6199 27675 6205
rect 31478 6196 31484 6208
rect 31536 6196 31542 6248
rect 31864 6245 31892 6276
rect 33226 6264 33232 6276
rect 33284 6264 33290 6316
rect 33686 6304 33692 6316
rect 33647 6276 33692 6304
rect 33686 6264 33692 6276
rect 33744 6304 33750 6316
rect 34698 6304 34704 6316
rect 33744 6276 34704 6304
rect 33744 6264 33750 6276
rect 34698 6264 34704 6276
rect 34756 6264 34762 6316
rect 35434 6264 35440 6316
rect 35492 6304 35498 6316
rect 36265 6307 36323 6313
rect 36265 6304 36277 6307
rect 35492 6276 36277 6304
rect 35492 6264 35498 6276
rect 36265 6273 36277 6276
rect 36311 6273 36323 6307
rect 36265 6267 36323 6273
rect 31849 6239 31907 6245
rect 31849 6205 31861 6239
rect 31895 6205 31907 6239
rect 31849 6199 31907 6205
rect 36354 6196 36360 6248
rect 36412 6236 36418 6248
rect 36449 6239 36507 6245
rect 36449 6236 36461 6239
rect 36412 6208 36461 6236
rect 36412 6196 36418 6208
rect 36449 6205 36461 6208
rect 36495 6236 36507 6239
rect 37090 6236 37096 6248
rect 36495 6208 37096 6236
rect 36495 6205 36507 6208
rect 36449 6199 36507 6205
rect 37090 6196 37096 6208
rect 37148 6196 37154 6248
rect 37604 6239 37662 6245
rect 37604 6205 37616 6239
rect 37650 6236 37662 6239
rect 38010 6236 38016 6248
rect 37650 6208 38016 6236
rect 37650 6205 37662 6208
rect 37604 6199 37662 6205
rect 38010 6196 38016 6208
rect 38068 6196 38074 6248
rect 14277 6171 14335 6177
rect 14277 6168 14289 6171
rect 12804 6140 13814 6168
rect 14200 6140 14289 6168
rect 12804 6137 12816 6140
rect 12758 6131 12816 6137
rect 14200 6112 14228 6140
rect 14277 6137 14289 6140
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 14366 6128 14372 6180
rect 14424 6168 14430 6180
rect 14424 6140 14469 6168
rect 14424 6128 14430 6140
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 16346 6171 16404 6177
rect 16346 6168 16358 6171
rect 15988 6140 16358 6168
rect 15988 6128 15994 6140
rect 16346 6137 16358 6140
rect 16392 6137 16404 6171
rect 18138 6168 18144 6180
rect 18099 6140 18144 6168
rect 16346 6131 16404 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 18288 6140 19073 6168
rect 18288 6128 18294 6140
rect 19061 6137 19073 6140
rect 19107 6137 19119 6171
rect 19061 6131 19119 6137
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 20901 6171 20959 6177
rect 20901 6168 20913 6171
rect 20588 6140 20913 6168
rect 20588 6128 20594 6140
rect 20901 6137 20913 6140
rect 20947 6137 20959 6171
rect 20901 6131 20959 6137
rect 20993 6171 21051 6177
rect 20993 6137 21005 6171
rect 21039 6137 21051 6171
rect 20993 6131 21051 6137
rect 10008 6072 10180 6100
rect 10008 6060 10014 6072
rect 13170 6060 13176 6112
rect 13228 6100 13234 6112
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 13228 6072 13369 6100
rect 13228 6060 13234 6072
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 14182 6060 14188 6112
rect 14240 6060 14246 6112
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20625 6103 20683 6109
rect 20625 6100 20637 6103
rect 19852 6072 20637 6100
rect 19852 6060 19858 6072
rect 20625 6069 20637 6072
rect 20671 6069 20683 6103
rect 21008 6100 21036 6131
rect 22830 6128 22836 6180
rect 22888 6168 22894 6180
rect 23477 6171 23535 6177
rect 23477 6168 23489 6171
rect 22888 6140 23489 6168
rect 22888 6128 22894 6140
rect 23477 6137 23489 6140
rect 23523 6168 23535 6171
rect 23934 6168 23940 6180
rect 23523 6140 23940 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23934 6128 23940 6140
rect 23992 6168 23998 6180
rect 24854 6168 24860 6180
rect 23992 6140 24860 6168
rect 23992 6128 23998 6140
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 25317 6171 25375 6177
rect 25317 6137 25329 6171
rect 25363 6168 25375 6171
rect 25590 6168 25596 6180
rect 25363 6140 25596 6168
rect 25363 6137 25375 6140
rect 25317 6131 25375 6137
rect 25590 6128 25596 6140
rect 25648 6168 25654 6180
rect 25771 6171 25829 6177
rect 25771 6168 25783 6171
rect 25648 6140 25783 6168
rect 25648 6128 25654 6140
rect 25771 6137 25783 6140
rect 25817 6168 25829 6171
rect 27062 6168 27068 6180
rect 25817 6140 27068 6168
rect 25817 6137 25829 6140
rect 25771 6131 25829 6137
rect 27062 6128 27068 6140
rect 27120 6128 27126 6180
rect 29730 6128 29736 6180
rect 29788 6168 29794 6180
rect 29917 6171 29975 6177
rect 29917 6168 29929 6171
rect 29788 6140 29929 6168
rect 29788 6128 29794 6140
rect 29917 6137 29929 6140
rect 29963 6137 29975 6171
rect 29917 6131 29975 6137
rect 30006 6128 30012 6180
rect 30064 6168 30070 6180
rect 30558 6168 30564 6180
rect 30064 6140 30109 6168
rect 30519 6140 30564 6168
rect 30064 6128 30070 6140
rect 30558 6128 30564 6140
rect 30616 6128 30622 6180
rect 32122 6168 32128 6180
rect 32083 6140 32128 6168
rect 32122 6128 32128 6140
rect 32180 6128 32186 6180
rect 33321 6171 33379 6177
rect 33321 6137 33333 6171
rect 33367 6168 33379 6171
rect 33410 6168 33416 6180
rect 33367 6140 33416 6168
rect 33367 6137 33379 6140
rect 33321 6131 33379 6137
rect 33410 6128 33416 6140
rect 33468 6128 33474 6180
rect 34701 6171 34759 6177
rect 34701 6137 34713 6171
rect 34747 6168 34759 6171
rect 34790 6168 34796 6180
rect 34747 6140 34796 6168
rect 34747 6137 34759 6140
rect 34701 6131 34759 6137
rect 34790 6128 34796 6140
rect 34848 6168 34854 6180
rect 34977 6171 35035 6177
rect 34977 6168 34989 6171
rect 34848 6140 34989 6168
rect 34848 6128 34854 6140
rect 34977 6137 34989 6140
rect 35023 6137 35035 6171
rect 34977 6131 35035 6137
rect 35066 6128 35072 6180
rect 35124 6168 35130 6180
rect 35124 6140 35169 6168
rect 35124 6128 35130 6140
rect 35250 6128 35256 6180
rect 35308 6168 35314 6180
rect 37691 6171 37749 6177
rect 37691 6168 37703 6171
rect 35308 6140 37703 6168
rect 35308 6128 35314 6140
rect 37691 6137 37703 6140
rect 37737 6137 37749 6171
rect 37691 6131 37749 6137
rect 21726 6100 21732 6112
rect 21008 6072 21732 6100
rect 20625 6063 20683 6069
rect 21726 6060 21732 6072
rect 21784 6060 21790 6112
rect 22370 6100 22376 6112
rect 22331 6072 22376 6100
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 22695 6103 22753 6109
rect 22695 6069 22707 6103
rect 22741 6100 22753 6103
rect 22922 6100 22928 6112
rect 22741 6072 22928 6100
rect 22741 6069 22753 6072
rect 22695 6063 22753 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23750 6100 23756 6112
rect 23711 6072 23756 6100
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 27246 6100 27252 6112
rect 27207 6072 27252 6100
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 30374 6060 30380 6112
rect 30432 6100 30438 6112
rect 30929 6103 30987 6109
rect 30929 6100 30941 6103
rect 30432 6072 30941 6100
rect 30432 6060 30438 6072
rect 30929 6069 30941 6072
rect 30975 6100 30987 6103
rect 31202 6100 31208 6112
rect 30975 6072 31208 6100
rect 30975 6069 30987 6072
rect 30929 6063 30987 6069
rect 31202 6060 31208 6072
rect 31260 6060 31266 6112
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1452 5868 1593 5896
rect 1452 5856 1458 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2406 5896 2412 5908
rect 1820 5868 2412 5896
rect 1820 5856 1826 5868
rect 2406 5856 2412 5868
rect 2464 5896 2470 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2464 5868 2881 5896
rect 2464 5856 2470 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3237 5899 3295 5905
rect 3237 5896 3249 5899
rect 3200 5868 3249 5896
rect 3200 5856 3206 5868
rect 3237 5865 3249 5868
rect 3283 5865 3295 5899
rect 3602 5896 3608 5908
rect 3563 5868 3608 5896
rect 3237 5859 3295 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 4154 5856 4160 5908
rect 4212 5905 4218 5908
rect 4212 5899 4261 5905
rect 4212 5865 4215 5899
rect 4249 5896 4261 5899
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4249 5868 4537 5896
rect 4249 5865 4261 5868
rect 4212 5859 4261 5865
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 4525 5859 4583 5865
rect 4212 5856 4218 5859
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6914 5896 6920 5908
rect 6595 5868 6920 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 8386 5896 8392 5908
rect 7208 5868 8392 5896
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 6825 5831 6883 5837
rect 6825 5828 6837 5831
rect 5224 5800 6837 5828
rect 5224 5788 5230 5800
rect 6825 5797 6837 5800
rect 6871 5828 6883 5831
rect 7098 5828 7104 5840
rect 6871 5800 7104 5828
rect 6871 5797 6883 5800
rect 6825 5791 6883 5797
rect 7098 5788 7104 5800
rect 7156 5788 7162 5840
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1912 5732 1961 5760
rect 1912 5720 1918 5732
rect 1949 5729 1961 5732
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 4132 5763 4190 5769
rect 4132 5729 4144 5763
rect 4178 5760 4190 5763
rect 4982 5760 4988 5772
rect 4178 5732 4988 5760
rect 4178 5729 4190 5732
rect 4132 5723 4190 5729
rect 1964 5692 1992 5723
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5442 5720 5448 5772
rect 5500 5760 5506 5772
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5500 5732 6009 5760
rect 5500 5720 5506 5732
rect 5997 5729 6009 5732
rect 6043 5760 6055 5763
rect 7208 5760 7236 5868
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 11146 5896 11152 5908
rect 11107 5868 11152 5896
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12437 5899 12495 5905
rect 12437 5896 12449 5899
rect 12124 5868 12449 5896
rect 12124 5856 12130 5868
rect 12437 5865 12449 5868
rect 12483 5865 12495 5899
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 12437 5859 12495 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18598 5896 18604 5908
rect 18196 5868 18604 5896
rect 18196 5856 18202 5868
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 22922 5856 22928 5908
rect 22980 5896 22986 5908
rect 24857 5899 24915 5905
rect 24857 5896 24869 5899
rect 22980 5868 24869 5896
rect 22980 5856 22986 5868
rect 24857 5865 24869 5868
rect 24903 5896 24915 5899
rect 24946 5896 24952 5908
rect 24903 5868 24952 5896
rect 24903 5865 24915 5868
rect 24857 5859 24915 5865
rect 24946 5856 24952 5868
rect 25004 5856 25010 5908
rect 26694 5896 26700 5908
rect 26655 5868 26700 5896
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 33226 5856 33232 5908
rect 33284 5896 33290 5908
rect 34057 5899 34115 5905
rect 34057 5896 34069 5899
rect 33284 5868 34069 5896
rect 33284 5856 33290 5868
rect 34057 5865 34069 5868
rect 34103 5865 34115 5899
rect 34057 5859 34115 5865
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 8662 5828 8668 5840
rect 7432 5800 8668 5828
rect 7432 5788 7438 5800
rect 8662 5788 8668 5800
rect 8720 5828 8726 5840
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8720 5800 8953 5828
rect 8720 5788 8726 5800
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10229 5831 10287 5837
rect 10229 5828 10241 5831
rect 10192 5800 10241 5828
rect 10192 5788 10198 5800
rect 10229 5797 10241 5800
rect 10275 5797 10287 5831
rect 10778 5828 10784 5840
rect 10739 5800 10784 5828
rect 10229 5791 10287 5797
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 13170 5828 13176 5840
rect 13131 5800 13176 5828
rect 13170 5788 13176 5800
rect 13228 5828 13234 5840
rect 15102 5828 15108 5840
rect 13228 5800 15108 5828
rect 13228 5788 13234 5800
rect 15102 5788 15108 5800
rect 15160 5828 15166 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 15160 5800 15485 5828
rect 15160 5788 15166 5800
rect 15473 5797 15485 5800
rect 15519 5797 15531 5831
rect 15473 5791 15531 5797
rect 16942 5788 16948 5840
rect 17000 5828 17006 5840
rect 17402 5828 17408 5840
rect 17000 5800 17408 5828
rect 17000 5788 17006 5800
rect 17402 5788 17408 5800
rect 17460 5828 17466 5840
rect 17773 5831 17831 5837
rect 17773 5828 17785 5831
rect 17460 5800 17785 5828
rect 17460 5788 17466 5800
rect 17773 5797 17785 5800
rect 17819 5797 17831 5831
rect 17773 5791 17831 5797
rect 18046 5788 18052 5840
rect 18104 5828 18110 5840
rect 19981 5831 20039 5837
rect 18104 5800 19288 5828
rect 18104 5788 18110 5800
rect 19260 5772 19288 5800
rect 19981 5797 19993 5831
rect 20027 5828 20039 5831
rect 20622 5828 20628 5840
rect 20027 5800 20628 5828
rect 20027 5797 20039 5800
rect 19981 5791 20039 5797
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 21174 5828 21180 5840
rect 21087 5800 21180 5828
rect 21174 5788 21180 5800
rect 21232 5828 21238 5840
rect 21815 5831 21873 5837
rect 21815 5828 21827 5831
rect 21232 5800 21827 5828
rect 21232 5788 21238 5800
rect 21815 5797 21827 5800
rect 21861 5828 21873 5831
rect 21910 5828 21916 5840
rect 21861 5800 21916 5828
rect 21861 5797 21873 5800
rect 21815 5791 21873 5797
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 23290 5788 23296 5840
rect 23348 5828 23354 5840
rect 23563 5831 23621 5837
rect 23563 5828 23575 5831
rect 23348 5800 23575 5828
rect 23348 5788 23354 5800
rect 23563 5797 23575 5800
rect 23609 5828 23621 5831
rect 25590 5828 25596 5840
rect 23609 5800 25596 5828
rect 23609 5797 23621 5800
rect 23563 5791 23621 5797
rect 25590 5788 25596 5800
rect 25648 5788 25654 5840
rect 27154 5788 27160 5840
rect 27212 5828 27218 5840
rect 27427 5831 27485 5837
rect 27427 5828 27439 5831
rect 27212 5800 27439 5828
rect 27212 5788 27218 5800
rect 27427 5797 27439 5800
rect 27473 5828 27485 5831
rect 28994 5828 29000 5840
rect 27473 5800 29000 5828
rect 27473 5797 27485 5800
rect 27427 5791 27485 5797
rect 28994 5788 29000 5800
rect 29052 5828 29058 5840
rect 29778 5831 29836 5837
rect 29778 5828 29790 5831
rect 29052 5800 29790 5828
rect 29052 5788 29058 5800
rect 29778 5797 29790 5800
rect 29824 5797 29836 5831
rect 29778 5791 29836 5797
rect 32490 5788 32496 5840
rect 32548 5828 32554 5840
rect 32630 5831 32688 5837
rect 32630 5828 32642 5831
rect 32548 5800 32642 5828
rect 32548 5788 32554 5800
rect 32630 5797 32642 5800
rect 32676 5797 32688 5831
rect 34606 5828 34612 5840
rect 34567 5800 34612 5828
rect 32630 5791 32688 5797
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 6043 5732 7236 5760
rect 7837 5763 7895 5769
rect 6043 5729 6055 5732
rect 5997 5723 6055 5729
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8018 5760 8024 5772
rect 7883 5732 8024 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8478 5760 8484 5772
rect 8435 5732 8484 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 11606 5760 11612 5772
rect 11567 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 11790 5760 11796 5772
rect 11751 5732 11796 5760
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 19242 5760 19248 5772
rect 19155 5732 19248 5760
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 6638 5692 6644 5704
rect 1964 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5692 6702 5704
rect 7190 5692 7196 5704
rect 6696 5664 7196 5692
rect 6696 5652 6702 5664
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7466 5692 7472 5704
rect 7379 5664 7472 5692
rect 2130 5624 2136 5636
rect 2091 5596 2136 5624
rect 2130 5584 2136 5596
rect 2188 5584 2194 5636
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4304 5528 4905 5556
rect 4304 5516 4310 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 4893 5519 4951 5525
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7392 5565 7420 5664
rect 7466 5652 7472 5664
rect 7524 5692 7530 5704
rect 8110 5692 8116 5704
rect 7524 5664 8116 5692
rect 7524 5652 7530 5664
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 8168 5664 8309 5692
rect 8168 5652 8174 5664
rect 8297 5661 8309 5664
rect 8343 5661 8355 5695
rect 8662 5692 8668 5704
rect 8623 5664 8668 5692
rect 8297 5655 8355 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10226 5692 10232 5704
rect 10183 5664 10232 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 13078 5692 13084 5704
rect 13039 5664 13084 5692
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 14884 5664 15393 5692
rect 14884 5652 14890 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15381 5655 15439 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 17497 5695 17555 5701
rect 15856 5664 16988 5692
rect 13630 5624 13636 5636
rect 13543 5596 13636 5624
rect 13630 5584 13636 5596
rect 13688 5624 13694 5636
rect 15856 5624 15884 5664
rect 13688 5596 15884 5624
rect 16960 5624 16988 5664
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 17543 5664 17693 5692
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 17681 5661 17693 5664
rect 17727 5692 17739 5695
rect 18322 5692 18328 5704
rect 17727 5664 18328 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 19702 5652 19708 5704
rect 19760 5692 19766 5704
rect 19812 5692 19840 5723
rect 20806 5720 20812 5772
rect 20864 5760 20870 5772
rect 21453 5763 21511 5769
rect 21453 5760 21465 5763
rect 20864 5732 21465 5760
rect 20864 5720 20870 5732
rect 21453 5729 21465 5732
rect 21499 5760 21511 5763
rect 22738 5760 22744 5772
rect 21499 5732 22744 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 22738 5720 22744 5732
rect 22796 5720 22802 5772
rect 23201 5763 23259 5769
rect 23201 5729 23213 5763
rect 23247 5760 23259 5763
rect 23750 5760 23756 5772
rect 23247 5732 23756 5760
rect 23247 5729 23259 5732
rect 23201 5723 23259 5729
rect 23750 5720 23756 5732
rect 23808 5720 23814 5772
rect 25016 5763 25074 5769
rect 25016 5729 25028 5763
rect 25062 5760 25074 5763
rect 25130 5760 25136 5772
rect 25062 5732 25136 5760
rect 25062 5729 25074 5732
rect 25016 5723 25074 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 27065 5763 27123 5769
rect 27065 5729 27077 5763
rect 27111 5760 27123 5763
rect 27246 5760 27252 5772
rect 27111 5732 27252 5760
rect 27111 5729 27123 5732
rect 27065 5723 27123 5729
rect 27246 5720 27252 5732
rect 27304 5720 27310 5772
rect 29270 5720 29276 5772
rect 29328 5760 29334 5772
rect 29457 5763 29515 5769
rect 29457 5760 29469 5763
rect 29328 5732 29469 5760
rect 29328 5720 29334 5732
rect 29457 5729 29469 5732
rect 29503 5729 29515 5763
rect 29457 5723 29515 5729
rect 32122 5720 32128 5772
rect 32180 5760 32186 5772
rect 32309 5763 32367 5769
rect 32309 5760 32321 5763
rect 32180 5732 32321 5760
rect 32180 5720 32186 5732
rect 32309 5729 32321 5732
rect 32355 5729 32367 5763
rect 32309 5723 32367 5729
rect 35526 5720 35532 5772
rect 35584 5760 35590 5772
rect 36024 5763 36082 5769
rect 36024 5760 36036 5763
rect 35584 5732 36036 5760
rect 35584 5720 35590 5732
rect 36024 5729 36036 5732
rect 36070 5760 36082 5763
rect 36722 5760 36728 5772
rect 36070 5732 36728 5760
rect 36070 5729 36082 5732
rect 36024 5723 36082 5729
rect 36722 5720 36728 5732
rect 36780 5720 36786 5772
rect 24670 5692 24676 5704
rect 19760 5664 24676 5692
rect 19760 5652 19766 5664
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 33134 5652 33140 5704
rect 33192 5692 33198 5704
rect 34146 5692 34152 5704
rect 33192 5664 34152 5692
rect 33192 5652 33198 5664
rect 34146 5652 34152 5664
rect 34204 5692 34210 5704
rect 34517 5695 34575 5701
rect 34517 5692 34529 5695
rect 34204 5664 34529 5692
rect 34204 5652 34210 5664
rect 34517 5661 34529 5664
rect 34563 5661 34575 5695
rect 34517 5655 34575 5661
rect 34698 5652 34704 5704
rect 34756 5692 34762 5704
rect 34793 5695 34851 5701
rect 34793 5692 34805 5695
rect 34756 5664 34805 5692
rect 34756 5652 34762 5664
rect 34793 5661 34805 5664
rect 34839 5661 34851 5695
rect 34793 5655 34851 5661
rect 18233 5627 18291 5633
rect 18233 5624 18245 5627
rect 16960 5596 18245 5624
rect 13688 5584 13694 5596
rect 18233 5593 18245 5596
rect 18279 5624 18291 5627
rect 18414 5624 18420 5636
rect 18279 5596 18420 5624
rect 18279 5593 18291 5596
rect 18233 5587 18291 5593
rect 18414 5584 18420 5596
rect 18472 5584 18478 5636
rect 29730 5584 29736 5636
rect 29788 5624 29794 5636
rect 30653 5627 30711 5633
rect 30653 5624 30665 5627
rect 29788 5596 30665 5624
rect 29788 5584 29794 5596
rect 30653 5593 30665 5596
rect 30699 5593 30711 5627
rect 30653 5587 30711 5593
rect 7377 5559 7435 5565
rect 7377 5556 7389 5559
rect 6604 5528 7389 5556
rect 6604 5516 6610 5528
rect 7377 5525 7389 5528
rect 7423 5525 7435 5559
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 7377 5519 7435 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 11882 5556 11888 5568
rect 11843 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5556 12955 5559
rect 12986 5556 12992 5568
rect 12943 5528 12992 5556
rect 12943 5525 12955 5528
rect 12897 5519 12955 5525
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 14182 5556 14188 5568
rect 13504 5528 14188 5556
rect 13504 5516 13510 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 16298 5556 16304 5568
rect 16259 5528 16304 5556
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 16666 5556 16672 5568
rect 16627 5528 16672 5556
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 22186 5516 22192 5568
rect 22244 5556 22250 5568
rect 22373 5559 22431 5565
rect 22373 5556 22385 5559
rect 22244 5528 22385 5556
rect 22244 5516 22250 5528
rect 22373 5525 22385 5528
rect 22419 5525 22431 5559
rect 24118 5556 24124 5568
rect 24079 5528 24124 5556
rect 22373 5519 22431 5525
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 24394 5556 24400 5568
rect 24355 5528 24400 5556
rect 24394 5516 24400 5528
rect 24452 5516 24458 5568
rect 25087 5559 25145 5565
rect 25087 5525 25099 5559
rect 25133 5556 25145 5559
rect 25314 5556 25320 5568
rect 25133 5528 25320 5556
rect 25133 5525 25145 5528
rect 25087 5519 25145 5525
rect 25314 5516 25320 5528
rect 25372 5516 25378 5568
rect 25498 5556 25504 5568
rect 25459 5528 25504 5556
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 27982 5556 27988 5568
rect 27943 5528 27988 5556
rect 27982 5516 27988 5528
rect 28040 5516 28046 5568
rect 29914 5516 29920 5568
rect 29972 5556 29978 5568
rect 30377 5559 30435 5565
rect 30377 5556 30389 5559
rect 29972 5528 30389 5556
rect 29972 5516 29978 5528
rect 30377 5525 30389 5528
rect 30423 5525 30435 5559
rect 31478 5556 31484 5568
rect 31391 5528 31484 5556
rect 30377 5519 30435 5525
rect 31478 5516 31484 5528
rect 31536 5556 31542 5568
rect 32214 5556 32220 5568
rect 31536 5528 32220 5556
rect 31536 5516 31542 5528
rect 32214 5516 32220 5528
rect 32272 5516 32278 5568
rect 33229 5559 33287 5565
rect 33229 5525 33241 5559
rect 33275 5556 33287 5559
rect 33318 5556 33324 5568
rect 33275 5528 33324 5556
rect 33275 5525 33287 5528
rect 33229 5519 33287 5525
rect 33318 5516 33324 5528
rect 33376 5516 33382 5568
rect 33594 5516 33600 5568
rect 33652 5556 33658 5568
rect 33689 5559 33747 5565
rect 33689 5556 33701 5559
rect 33652 5528 33701 5556
rect 33652 5516 33658 5528
rect 33689 5525 33701 5528
rect 33735 5525 33747 5559
rect 33689 5519 33747 5525
rect 35894 5516 35900 5568
rect 35952 5556 35958 5568
rect 36127 5559 36185 5565
rect 36127 5556 36139 5559
rect 35952 5528 36139 5556
rect 35952 5516 35958 5528
rect 36127 5525 36139 5528
rect 36173 5525 36185 5559
rect 36127 5519 36185 5525
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2924 5324 3157 5352
rect 2924 5312 2930 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 5442 5352 5448 5364
rect 5403 5324 5448 5352
rect 3145 5315 3203 5321
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 7282 5352 7288 5364
rect 6319 5324 7288 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 4982 5284 4988 5296
rect 4895 5256 4988 5284
rect 4982 5244 4988 5256
rect 5040 5284 5046 5296
rect 5810 5284 5816 5296
rect 5040 5256 5816 5284
rect 5040 5244 5046 5256
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5166 5216 5172 5228
rect 4663 5188 5172 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 2406 5148 2412 5160
rect 2367 5120 2412 5148
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 2866 5148 2872 5160
rect 2731 5120 2872 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6288 5148 6316 5315
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 9180 5324 9229 5352
rect 9180 5312 9186 5324
rect 9217 5321 9229 5324
rect 9263 5321 9275 5355
rect 9217 5315 9275 5321
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10192 5324 10609 5352
rect 10192 5312 10198 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 10597 5315 10655 5321
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 11977 5355 12035 5361
rect 11977 5352 11989 5355
rect 11664 5324 11989 5352
rect 11664 5312 11670 5324
rect 11977 5321 11989 5324
rect 12023 5321 12035 5355
rect 11977 5315 12035 5321
rect 13081 5355 13139 5361
rect 13081 5321 13093 5355
rect 13127 5352 13139 5355
rect 13170 5352 13176 5364
rect 13127 5324 13176 5352
rect 13127 5321 13139 5324
rect 13081 5315 13139 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13722 5352 13728 5364
rect 13311 5324 13728 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 14826 5352 14832 5364
rect 14787 5324 14832 5352
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 15102 5352 15108 5364
rect 15063 5324 15108 5352
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 17954 5352 17960 5364
rect 17911 5324 17960 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 20027 5355 20085 5361
rect 20027 5321 20039 5355
rect 20073 5352 20085 5355
rect 20530 5352 20536 5364
rect 20073 5324 20536 5352
rect 20073 5321 20085 5324
rect 20027 5315 20085 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20806 5352 20812 5364
rect 20767 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21910 5352 21916 5364
rect 21823 5324 21916 5352
rect 21910 5312 21916 5324
rect 21968 5352 21974 5364
rect 23290 5352 23296 5364
rect 21968 5324 23296 5352
rect 21968 5312 21974 5324
rect 23290 5312 23296 5324
rect 23348 5312 23354 5364
rect 25041 5355 25099 5361
rect 25041 5321 25053 5355
rect 25087 5352 25099 5355
rect 25130 5352 25136 5364
rect 25087 5324 25136 5352
rect 25087 5321 25099 5324
rect 25041 5315 25099 5321
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 26789 5355 26847 5361
rect 26789 5321 26801 5355
rect 26835 5352 26847 5355
rect 27246 5352 27252 5364
rect 26835 5324 27252 5352
rect 26835 5321 26847 5324
rect 26789 5315 26847 5321
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 28721 5355 28779 5361
rect 28721 5321 28733 5355
rect 28767 5352 28779 5355
rect 29270 5352 29276 5364
rect 28767 5324 29276 5352
rect 28767 5321 28779 5324
rect 28721 5315 28779 5321
rect 29270 5312 29276 5324
rect 29328 5312 29334 5364
rect 30006 5312 30012 5364
rect 30064 5352 30070 5364
rect 30377 5355 30435 5361
rect 30377 5352 30389 5355
rect 30064 5324 30389 5352
rect 30064 5312 30070 5324
rect 30377 5321 30389 5324
rect 30423 5321 30435 5355
rect 30377 5315 30435 5321
rect 34517 5355 34575 5361
rect 34517 5321 34529 5355
rect 34563 5352 34575 5355
rect 34606 5352 34612 5364
rect 34563 5324 34612 5352
rect 34563 5321 34575 5324
rect 34517 5315 34575 5321
rect 34606 5312 34612 5324
rect 34664 5312 34670 5364
rect 36035 5355 36093 5361
rect 36035 5321 36047 5355
rect 36081 5352 36093 5355
rect 36538 5352 36544 5364
rect 36081 5324 36544 5352
rect 36081 5321 36093 5324
rect 36035 5315 36093 5321
rect 36538 5312 36544 5324
rect 36596 5312 36602 5364
rect 36722 5352 36728 5364
rect 36683 5324 36728 5352
rect 36722 5312 36728 5324
rect 36780 5312 36786 5364
rect 8294 5284 8300 5296
rect 8036 5256 8300 5284
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7248 5188 7297 5216
rect 7248 5176 7254 5188
rect 7285 5185 7297 5188
rect 7331 5216 7343 5219
rect 8036 5216 8064 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10321 5287 10379 5293
rect 10321 5284 10333 5287
rect 10008 5256 10333 5284
rect 10008 5244 10014 5256
rect 10321 5253 10333 5256
rect 10367 5253 10379 5287
rect 10321 5247 10379 5253
rect 12667 5287 12725 5293
rect 12667 5253 12679 5287
rect 12713 5284 12725 5287
rect 15378 5284 15384 5296
rect 12713 5256 15384 5284
rect 12713 5253 12725 5256
rect 12667 5247 12725 5253
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 15473 5287 15531 5293
rect 15473 5253 15485 5287
rect 15519 5284 15531 5287
rect 18230 5284 18236 5296
rect 15519 5256 18236 5284
rect 15519 5253 15531 5256
rect 15473 5247 15531 5253
rect 18230 5244 18236 5256
rect 18288 5244 18294 5296
rect 20622 5244 20628 5296
rect 20680 5284 20686 5296
rect 21085 5287 21143 5293
rect 21085 5284 21097 5287
rect 20680 5256 21097 5284
rect 20680 5244 20686 5256
rect 21085 5253 21097 5256
rect 21131 5253 21143 5287
rect 21085 5247 21143 5253
rect 22649 5287 22707 5293
rect 22649 5253 22661 5287
rect 22695 5284 22707 5287
rect 26973 5287 27031 5293
rect 22695 5256 25636 5284
rect 22695 5253 22707 5256
rect 22649 5247 22707 5253
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 7331 5188 8064 5216
rect 8128 5188 8861 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 8128 5160 8156 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 13630 5216 13636 5228
rect 13591 5188 13636 5216
rect 8849 5179 8907 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 13906 5216 13912 5228
rect 13780 5188 13912 5216
rect 13780 5176 13786 5188
rect 13906 5176 13912 5188
rect 13964 5216 13970 5228
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 13964 5188 14289 5216
rect 13964 5176 13970 5188
rect 14277 5185 14289 5188
rect 14323 5216 14335 5219
rect 14642 5216 14648 5228
rect 14323 5188 14648 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 14918 5176 14924 5228
rect 14976 5176 14982 5228
rect 15654 5176 15660 5228
rect 15712 5216 15718 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 15712 5188 16773 5216
rect 15712 5176 15718 5188
rect 16761 5185 16773 5188
rect 16807 5216 16819 5219
rect 17586 5216 17592 5228
rect 16807 5188 17592 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 18782 5216 18788 5228
rect 18743 5188 18788 5216
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 22094 5216 22100 5228
rect 21468 5188 22100 5216
rect 5767 5120 6316 5148
rect 7745 5151 7803 5157
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 7745 5117 7757 5151
rect 7791 5117 7803 5151
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 7745 5111 7803 5117
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 1728 5052 3709 5080
rect 1728 5040 1734 5052
rect 3697 5049 3709 5052
rect 3743 5080 3755 5083
rect 3988 5080 4016 5111
rect 3743 5052 4016 5080
rect 6641 5083 6699 5089
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7190 5080 7196 5092
rect 6687 5052 7196 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6656 5012 6684 5043
rect 7190 5040 7196 5052
rect 7248 5080 7254 5092
rect 7760 5080 7788 5111
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8294 5148 8300 5160
rect 8255 5120 8300 5148
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 9398 5148 9404 5160
rect 8619 5120 9404 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 11200 5151 11258 5157
rect 11200 5117 11212 5151
rect 11246 5148 11258 5151
rect 11246 5120 11744 5148
rect 11246 5117 11258 5120
rect 11200 5111 11258 5117
rect 8018 5080 8024 5092
rect 7248 5052 8024 5080
rect 7248 5040 7254 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9722 5083 9780 5089
rect 9722 5080 9734 5083
rect 9180 5052 9734 5080
rect 9180 5040 9186 5052
rect 9722 5049 9734 5052
rect 9768 5049 9780 5083
rect 9722 5043 9780 5049
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 11287 5083 11345 5089
rect 11287 5080 11299 5083
rect 10284 5052 11299 5080
rect 10284 5040 10290 5052
rect 11287 5049 11299 5052
rect 11333 5049 11345 5083
rect 11287 5043 11345 5049
rect 11716 5024 11744 5120
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 12596 5151 12654 5157
rect 12596 5148 12608 5151
rect 12124 5120 12608 5148
rect 12124 5108 12130 5120
rect 12596 5117 12608 5120
rect 12642 5148 12654 5151
rect 13265 5151 13323 5157
rect 13265 5148 13277 5151
rect 12642 5120 13277 5148
rect 12642 5117 12654 5120
rect 12596 5111 12654 5117
rect 13265 5117 13277 5120
rect 13311 5117 13323 5151
rect 14936 5148 14964 5176
rect 15277 5151 15335 5157
rect 15277 5148 15289 5151
rect 14936 5120 15289 5148
rect 13265 5111 13323 5117
rect 15277 5117 15289 5120
rect 15323 5148 15335 5151
rect 15838 5148 15844 5160
rect 15323 5120 15844 5148
rect 15323 5117 15335 5120
rect 15277 5111 15335 5117
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 17954 5148 17960 5160
rect 17736 5120 17960 5148
rect 17736 5108 17742 5120
rect 17954 5108 17960 5120
rect 18012 5148 18018 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 18012 5120 18061 5148
rect 18012 5108 18018 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18506 5148 18512 5160
rect 18467 5120 18512 5148
rect 18049 5111 18107 5117
rect 18506 5108 18512 5120
rect 18564 5148 18570 5160
rect 19702 5148 19708 5160
rect 18564 5120 19708 5148
rect 18564 5108 18570 5120
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 21468 5157 21496 5188
rect 22094 5176 22100 5188
rect 22152 5176 22158 5228
rect 23198 5176 23204 5228
rect 23256 5216 23262 5228
rect 23753 5219 23811 5225
rect 23753 5216 23765 5219
rect 23256 5188 23765 5216
rect 23256 5176 23262 5188
rect 23753 5185 23765 5188
rect 23799 5216 23811 5219
rect 24394 5216 24400 5228
rect 23799 5188 24400 5216
rect 23799 5185 23811 5188
rect 23753 5179 23811 5185
rect 24394 5176 24400 5188
rect 24452 5176 24458 5228
rect 25314 5216 25320 5228
rect 25275 5188 25320 5216
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 25608 5225 25636 5256
rect 26973 5253 26985 5287
rect 27019 5284 27031 5287
rect 28261 5287 28319 5293
rect 28261 5284 28273 5287
rect 27019 5256 28273 5284
rect 27019 5253 27031 5256
rect 26973 5247 27031 5253
rect 28261 5253 28273 5256
rect 28307 5284 28319 5287
rect 29730 5284 29736 5296
rect 28307 5256 29736 5284
rect 28307 5253 28319 5256
rect 28261 5247 28319 5253
rect 29730 5244 29736 5256
rect 29788 5244 29794 5296
rect 30558 5244 30564 5296
rect 30616 5284 30622 5296
rect 36446 5284 36452 5296
rect 30616 5256 33548 5284
rect 36407 5256 36452 5284
rect 30616 5244 30622 5256
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5216 25651 5219
rect 28166 5216 28172 5228
rect 25639 5188 28172 5216
rect 25639 5185 25651 5188
rect 25593 5179 25651 5185
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 28994 5216 29000 5228
rect 28955 5188 29000 5216
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 29457 5219 29515 5225
rect 29457 5185 29469 5219
rect 29503 5216 29515 5219
rect 29546 5216 29552 5228
rect 29503 5188 29552 5216
rect 29503 5185 29515 5188
rect 29457 5179 29515 5185
rect 29546 5176 29552 5188
rect 29604 5216 29610 5228
rect 33520 5225 33548 5256
rect 36446 5244 36452 5256
rect 36504 5244 36510 5296
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 29604 5188 30665 5216
rect 29604 5176 29610 5188
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 31113 5219 31171 5225
rect 31113 5185 31125 5219
rect 31159 5216 31171 5219
rect 33505 5219 33563 5225
rect 31159 5188 31800 5216
rect 31159 5185 31171 5188
rect 31113 5179 31171 5185
rect 19935 5151 19993 5157
rect 19935 5117 19947 5151
rect 19981 5117 19993 5151
rect 19935 5111 19993 5117
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5148 20959 5151
rect 21453 5151 21511 5157
rect 21453 5148 21465 5151
rect 20947 5120 21465 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21453 5117 21465 5120
rect 21499 5117 21511 5151
rect 27154 5148 27160 5160
rect 27115 5120 27160 5148
rect 21453 5111 21511 5117
rect 13725 5083 13783 5089
rect 13725 5049 13737 5083
rect 13771 5080 13783 5083
rect 13814 5080 13820 5092
rect 13771 5052 13820 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 11698 5012 11704 5024
rect 5951 4984 6684 5012
rect 11659 4984 11704 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 13449 5015 13507 5021
rect 13449 4981 13461 5015
rect 13495 5012 13507 5015
rect 13740 5012 13768 5043
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 16482 5080 16488 5092
rect 16443 5052 16488 5080
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16632 5052 16677 5080
rect 16632 5040 16638 5052
rect 17218 5040 17224 5092
rect 17276 5080 17282 5092
rect 19950 5080 19978 5111
rect 27154 5108 27160 5120
rect 27212 5108 27218 5160
rect 20349 5083 20407 5089
rect 20349 5080 20361 5083
rect 17276 5052 20361 5080
rect 17276 5040 17282 5052
rect 20349 5049 20361 5052
rect 20395 5080 20407 5083
rect 21358 5080 21364 5092
rect 20395 5052 21364 5080
rect 20395 5049 20407 5052
rect 20349 5043 20407 5049
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 22094 5080 22100 5092
rect 22055 5052 22100 5080
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 22186 5040 22192 5092
rect 22244 5080 22250 5092
rect 22244 5052 23474 5080
rect 22244 5040 22250 5052
rect 13495 4984 13768 5012
rect 16301 5015 16359 5021
rect 13495 4981 13507 4984
rect 13449 4975 13507 4981
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16592 5012 16620 5040
rect 16347 4984 16620 5012
rect 23446 5012 23474 5052
rect 23842 5040 23848 5092
rect 23900 5080 23906 5092
rect 24394 5080 24400 5092
rect 23900 5052 23945 5080
rect 24355 5052 24400 5080
rect 23900 5040 23906 5052
rect 24394 5040 24400 5052
rect 24452 5080 24458 5092
rect 25406 5080 25412 5092
rect 24452 5052 25268 5080
rect 25367 5052 25412 5080
rect 24452 5040 24458 5052
rect 23860 5012 23888 5040
rect 23446 4984 23888 5012
rect 25240 5012 25268 5052
rect 25406 5040 25412 5052
rect 25464 5040 25470 5092
rect 27522 5040 27528 5092
rect 27580 5080 27586 5092
rect 27709 5083 27767 5089
rect 27709 5080 27721 5083
rect 27580 5052 27721 5080
rect 27580 5040 27586 5052
rect 27709 5049 27721 5052
rect 27755 5049 27767 5083
rect 27709 5043 27767 5049
rect 27801 5083 27859 5089
rect 27801 5049 27813 5083
rect 27847 5080 27859 5083
rect 27982 5080 27988 5092
rect 27847 5052 27988 5080
rect 27847 5049 27859 5052
rect 27801 5043 27859 5049
rect 26973 5015 27031 5021
rect 26973 5012 26985 5015
rect 25240 4984 26985 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 26973 4981 26985 4984
rect 27019 4981 27031 5015
rect 26973 4975 27031 4981
rect 27433 5015 27491 5021
rect 27433 4981 27445 5015
rect 27479 5012 27491 5015
rect 27816 5012 27844 5043
rect 27982 5040 27988 5052
rect 28040 5040 28046 5092
rect 29012 5080 29040 5176
rect 31202 5148 31208 5160
rect 31163 5120 31208 5148
rect 31202 5108 31208 5120
rect 31260 5108 31266 5160
rect 31772 5157 31800 5188
rect 33505 5185 33517 5219
rect 33551 5216 33563 5219
rect 34606 5216 34612 5228
rect 33551 5188 34612 5216
rect 33551 5185 33563 5188
rect 33505 5179 33563 5185
rect 34606 5176 34612 5188
rect 34664 5176 34670 5228
rect 34790 5176 34796 5228
rect 34848 5216 34854 5228
rect 34885 5219 34943 5225
rect 34885 5216 34897 5219
rect 34848 5188 34897 5216
rect 34848 5176 34854 5188
rect 34885 5185 34897 5188
rect 34931 5185 34943 5219
rect 34885 5179 34943 5185
rect 31757 5151 31815 5157
rect 31757 5117 31769 5151
rect 31803 5148 31815 5151
rect 32582 5148 32588 5160
rect 31803 5120 32588 5148
rect 31803 5117 31815 5120
rect 31757 5111 31815 5117
rect 32582 5108 32588 5120
rect 32640 5108 32646 5160
rect 35964 5151 36022 5157
rect 35964 5117 35976 5151
rect 36010 5148 36022 5151
rect 36464 5148 36492 5244
rect 36010 5120 36492 5148
rect 36010 5117 36022 5120
rect 35964 5111 36022 5117
rect 29454 5080 29460 5092
rect 29012 5052 29460 5080
rect 29454 5040 29460 5052
rect 29512 5080 29518 5092
rect 29778 5083 29836 5089
rect 29778 5080 29790 5083
rect 29512 5052 29790 5080
rect 29512 5040 29518 5052
rect 29778 5049 29790 5052
rect 29824 5080 29836 5083
rect 32309 5083 32367 5089
rect 32309 5080 32321 5083
rect 29824 5052 32321 5080
rect 29824 5049 29836 5052
rect 29778 5043 29836 5049
rect 32309 5049 32321 5052
rect 32355 5080 32367 5083
rect 32490 5080 32496 5092
rect 32355 5052 32496 5080
rect 32355 5049 32367 5052
rect 32309 5043 32367 5049
rect 32490 5040 32496 5052
rect 32548 5040 32554 5092
rect 33045 5083 33103 5089
rect 33045 5049 33057 5083
rect 33091 5080 33103 5083
rect 33226 5080 33232 5092
rect 33091 5052 33232 5080
rect 33091 5049 33103 5052
rect 33045 5043 33103 5049
rect 33226 5040 33232 5052
rect 33284 5040 33290 5092
rect 33318 5040 33324 5092
rect 33376 5080 33382 5092
rect 33376 5052 33421 5080
rect 33376 5040 33382 5052
rect 31294 5012 31300 5024
rect 27479 4984 27844 5012
rect 31255 4984 31300 5012
rect 27479 4981 27491 4984
rect 27433 4975 27491 4981
rect 31294 4972 31300 4984
rect 31352 4972 31358 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 2866 4808 2872 4820
rect 2792 4780 2872 4808
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2590 4672 2596 4684
rect 2547 4644 2596 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 2792 4681 2820 4780
rect 2866 4768 2872 4780
rect 2924 4808 2930 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 2924 4780 5089 4808
rect 2924 4768 2930 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 5077 4771 5135 4777
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7282 4808 7288 4820
rect 7064 4780 7288 4808
rect 7064 4768 7070 4780
rect 7282 4768 7288 4780
rect 7340 4808 7346 4820
rect 8662 4808 8668 4820
rect 7340 4780 7604 4808
rect 8623 4780 8668 4808
rect 7340 4768 7346 4780
rect 2958 4740 2964 4752
rect 2919 4712 2964 4740
rect 2958 4700 2964 4712
rect 3016 4700 3022 4752
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 5500 4712 5917 4740
rect 5500 4700 5506 4712
rect 5905 4709 5917 4712
rect 5951 4740 5963 4743
rect 5994 4740 6000 4752
rect 5951 4712 6000 4740
rect 5951 4709 5963 4712
rect 5905 4703 5963 4709
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4641 2835 4675
rect 4890 4672 4896 4684
rect 4803 4644 4896 4672
rect 2777 4635 2835 4641
rect 4890 4632 4896 4644
rect 4948 4672 4954 4684
rect 5350 4672 5356 4684
rect 4948 4644 5356 4672
rect 4948 4632 4954 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 6972 4644 7297 4672
rect 6972 4632 6978 4644
rect 7285 4641 7297 4644
rect 7331 4672 7343 4675
rect 7374 4672 7380 4684
rect 7331 4644 7380 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 7576 4681 7604 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 9398 4808 9404 4820
rect 9359 4780 9404 4808
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10226 4808 10232 4820
rect 10183 4780 10232 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 11606 4808 11612 4820
rect 10704 4780 11612 4808
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 8076 4712 8401 4740
rect 8076 4700 8082 4712
rect 8389 4709 8401 4712
rect 8435 4740 8447 4743
rect 10704 4740 10732 4780
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 11790 4808 11796 4820
rect 11747 4780 11796 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12710 4808 12716 4820
rect 12671 4780 12716 4808
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13078 4808 13084 4820
rect 13039 4780 13084 4808
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 14826 4808 14832 4820
rect 13188 4780 14832 4808
rect 8435 4712 10732 4740
rect 10781 4743 10839 4749
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 10781 4709 10793 4743
rect 10827 4740 10839 4743
rect 10870 4740 10876 4752
rect 10827 4712 10876 4740
rect 10827 4709 10839 4712
rect 10781 4703 10839 4709
rect 10870 4700 10876 4712
rect 10928 4700 10934 4752
rect 12299 4743 12357 4749
rect 12299 4709 12311 4743
rect 12345 4740 12357 4743
rect 13188 4740 13216 4780
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 16482 4808 16488 4820
rect 16443 4780 16488 4808
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 18233 4811 18291 4817
rect 18233 4777 18245 4811
rect 18279 4808 18291 4811
rect 18506 4808 18512 4820
rect 18279 4780 18512 4808
rect 18279 4777 18291 4780
rect 18233 4771 18291 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 18598 4768 18604 4820
rect 18656 4808 18662 4820
rect 18831 4811 18889 4817
rect 18831 4808 18843 4811
rect 18656 4780 18843 4808
rect 18656 4768 18662 4780
rect 18831 4777 18843 4780
rect 18877 4777 18889 4811
rect 18831 4771 18889 4777
rect 21407 4811 21465 4817
rect 21407 4777 21419 4811
rect 21453 4808 21465 4811
rect 22094 4808 22100 4820
rect 21453 4780 22100 4808
rect 21453 4777 21465 4780
rect 21407 4771 21465 4777
rect 22094 4768 22100 4780
rect 22152 4808 22158 4820
rect 22373 4811 22431 4817
rect 22373 4808 22385 4811
rect 22152 4780 22385 4808
rect 22152 4768 22158 4780
rect 22373 4777 22385 4780
rect 22419 4777 22431 4811
rect 23198 4808 23204 4820
rect 23159 4780 23204 4808
rect 22373 4771 22431 4777
rect 23198 4768 23204 4780
rect 23256 4768 23262 4820
rect 23842 4808 23848 4820
rect 23803 4780 23848 4808
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 25314 4768 25320 4820
rect 25372 4808 25378 4820
rect 25593 4811 25651 4817
rect 25593 4808 25605 4811
rect 25372 4780 25605 4808
rect 25372 4768 25378 4780
rect 25593 4777 25605 4780
rect 25639 4777 25651 4811
rect 25593 4771 25651 4777
rect 27019 4811 27077 4817
rect 27019 4777 27031 4811
rect 27065 4808 27077 4811
rect 27522 4808 27528 4820
rect 27065 4780 27528 4808
rect 27065 4777 27077 4780
rect 27019 4771 27077 4777
rect 27522 4768 27528 4780
rect 27580 4808 27586 4820
rect 27617 4811 27675 4817
rect 27617 4808 27629 4811
rect 27580 4780 27629 4808
rect 27580 4768 27586 4780
rect 27617 4777 27629 4780
rect 27663 4777 27675 4811
rect 29454 4808 29460 4820
rect 29415 4780 29460 4808
rect 27617 4771 27675 4777
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 31202 4808 31208 4820
rect 31163 4780 31208 4808
rect 31202 4768 31208 4780
rect 31260 4768 31266 4820
rect 31941 4811 31999 4817
rect 31941 4777 31953 4811
rect 31987 4808 31999 4811
rect 32122 4808 32128 4820
rect 31987 4780 32128 4808
rect 31987 4777 31999 4780
rect 31941 4771 31999 4777
rect 32122 4768 32128 4780
rect 32180 4768 32186 4820
rect 33229 4811 33287 4817
rect 33229 4777 33241 4811
rect 33275 4808 33287 4811
rect 33318 4808 33324 4820
rect 33275 4780 33324 4808
rect 33275 4777 33287 4780
rect 33229 4771 33287 4777
rect 33318 4768 33324 4780
rect 33376 4768 33382 4820
rect 34146 4768 34152 4820
rect 34204 4808 34210 4820
rect 34425 4811 34483 4817
rect 34425 4808 34437 4811
rect 34204 4780 34437 4808
rect 34204 4768 34210 4780
rect 34425 4777 34437 4780
rect 34471 4777 34483 4811
rect 34425 4771 34483 4777
rect 12345 4712 13216 4740
rect 12345 4709 12357 4712
rect 12299 4703 12357 4709
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 13357 4743 13415 4749
rect 13357 4740 13369 4743
rect 13320 4712 13369 4740
rect 13320 4700 13326 4712
rect 13357 4709 13369 4712
rect 13403 4709 13415 4743
rect 13906 4740 13912 4752
rect 13867 4712 13912 4740
rect 13357 4703 13415 4709
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 16025 4743 16083 4749
rect 16025 4709 16037 4743
rect 16071 4740 16083 4743
rect 16666 4740 16672 4752
rect 16071 4712 16672 4740
rect 16071 4709 16083 4712
rect 16025 4703 16083 4709
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 17313 4743 17371 4749
rect 17313 4709 17325 4743
rect 17359 4740 17371 4743
rect 17402 4740 17408 4752
rect 17359 4712 17408 4740
rect 17359 4709 17371 4712
rect 17313 4703 17371 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 19935 4743 19993 4749
rect 19935 4709 19947 4743
rect 19981 4740 19993 4743
rect 22002 4740 22008 4752
rect 19981 4712 22008 4740
rect 19981 4709 19993 4712
rect 19935 4703 19993 4709
rect 22002 4700 22008 4712
rect 22060 4700 22066 4752
rect 23477 4743 23535 4749
rect 23477 4709 23489 4743
rect 23523 4740 23535 4743
rect 23750 4740 23756 4752
rect 23523 4712 23756 4740
rect 23523 4709 23535 4712
rect 23477 4703 23535 4709
rect 23750 4700 23756 4712
rect 23808 4700 23814 4752
rect 24118 4740 24124 4752
rect 24079 4712 24124 4740
rect 24118 4700 24124 4712
rect 24176 4740 24182 4752
rect 25225 4743 25283 4749
rect 25225 4740 25237 4743
rect 24176 4712 25237 4740
rect 24176 4700 24182 4712
rect 25225 4709 25237 4712
rect 25271 4740 25283 4743
rect 25406 4740 25412 4752
rect 25271 4712 25412 4740
rect 25271 4709 25283 4712
rect 25225 4703 25283 4709
rect 25406 4700 25412 4712
rect 25464 4700 25470 4752
rect 27982 4700 27988 4752
rect 28040 4740 28046 4752
rect 28077 4743 28135 4749
rect 28077 4740 28089 4743
rect 28040 4712 28089 4740
rect 28040 4700 28046 4712
rect 28077 4709 28089 4712
rect 28123 4709 28135 4743
rect 29914 4740 29920 4752
rect 29875 4712 29920 4740
rect 28077 4703 28135 4709
rect 29914 4700 29920 4712
rect 29972 4700 29978 4752
rect 30469 4743 30527 4749
rect 30469 4709 30481 4743
rect 30515 4740 30527 4743
rect 30558 4740 30564 4752
rect 30515 4712 30564 4740
rect 30515 4709 30527 4712
rect 30469 4703 30527 4709
rect 30558 4700 30564 4712
rect 30616 4700 30622 4752
rect 32858 4740 32864 4752
rect 32819 4712 32864 4740
rect 32858 4700 32864 4712
rect 32916 4700 32922 4752
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 12212 4675 12270 4681
rect 12212 4641 12224 4675
rect 12258 4672 12270 4675
rect 12434 4672 12440 4684
rect 12258 4644 12440 4672
rect 12258 4641 12270 4644
rect 12212 4635 12270 4641
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 15470 4672 15476 4684
rect 15431 4644 15476 4672
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4672 15899 4675
rect 15930 4672 15936 4684
rect 15887 4644 15936 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 18693 4675 18751 4681
rect 18693 4641 18705 4675
rect 18739 4672 18751 4675
rect 18782 4672 18788 4684
rect 18739 4644 18788 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 19794 4672 19800 4684
rect 19852 4681 19858 4684
rect 19852 4675 19890 4681
rect 18892 4644 19800 4672
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7524 4576 7757 4604
rect 7524 4564 7530 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 10778 4604 10784 4616
rect 10735 4576 10784 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 13265 4607 13323 4613
rect 13265 4573 13277 4607
rect 13311 4604 13323 4607
rect 15654 4604 15660 4616
rect 13311 4576 15660 4604
rect 13311 4573 13323 4576
rect 13265 4567 13323 4573
rect 6454 4496 6460 4548
rect 6512 4536 6518 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6512 4508 7389 4536
rect 6512 4496 6518 4508
rect 7377 4505 7389 4508
rect 7423 4536 7435 4539
rect 8018 4536 8024 4548
rect 7423 4508 8024 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8018 4496 8024 4508
rect 8076 4496 8082 4548
rect 11238 4536 11244 4548
rect 11199 4508 11244 4536
rect 11238 4496 11244 4508
rect 11296 4496 11302 4548
rect 13170 4496 13176 4548
rect 13228 4536 13234 4548
rect 13280 4536 13308 4567
rect 15654 4564 15660 4576
rect 15712 4564 15718 4616
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4604 17279 4607
rect 17494 4604 17500 4616
rect 17267 4576 17500 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 17586 4564 17592 4616
rect 17644 4604 17650 4616
rect 17644 4576 17689 4604
rect 17644 4564 17650 4576
rect 13228 4508 13308 4536
rect 13228 4496 13234 4508
rect 13630 4496 13636 4548
rect 13688 4536 13694 4548
rect 13688 4508 13814 4536
rect 13688 4496 13694 4508
rect 7193 4471 7251 4477
rect 7193 4437 7205 4471
rect 7239 4468 7251 4471
rect 8478 4468 8484 4480
rect 7239 4440 8484 4468
rect 7239 4437 7251 4440
rect 7193 4431 7251 4437
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 13786 4468 13814 4508
rect 15838 4496 15844 4548
rect 15896 4536 15902 4548
rect 18892 4536 18920 4644
rect 19794 4632 19800 4644
rect 19878 4641 19890 4675
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 19852 4635 19890 4641
rect 19852 4632 19858 4635
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4672 22155 4675
rect 22186 4672 22192 4684
rect 22143 4644 22192 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 22992 4675 23050 4681
rect 22992 4641 23004 4675
rect 23038 4672 23050 4675
rect 23106 4672 23112 4684
rect 23038 4644 23112 4672
rect 23038 4641 23050 4644
rect 22992 4635 23050 4641
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 26948 4675 27006 4681
rect 26948 4672 26960 4675
rect 24688 4644 26960 4672
rect 24026 4604 24032 4616
rect 23987 4576 24032 4604
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 24394 4604 24400 4616
rect 24355 4576 24400 4604
rect 24394 4564 24400 4576
rect 24452 4564 24458 4616
rect 24688 4604 24716 4644
rect 26948 4641 26960 4644
rect 26994 4672 27006 4675
rect 27614 4672 27620 4684
rect 26994 4644 27620 4672
rect 26994 4641 27006 4644
rect 26948 4635 27006 4641
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 32125 4675 32183 4681
rect 32125 4641 32137 4675
rect 32171 4641 32183 4675
rect 32582 4672 32588 4684
rect 32543 4644 32588 4672
rect 32125 4635 32183 4641
rect 27982 4604 27988 4616
rect 24504 4576 24716 4604
rect 27943 4576 27988 4604
rect 15896 4508 18920 4536
rect 15896 4496 15902 4508
rect 23014 4496 23020 4548
rect 23072 4536 23078 4548
rect 24504 4536 24532 4576
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 28166 4564 28172 4616
rect 28224 4604 28230 4616
rect 28261 4607 28319 4613
rect 28261 4604 28273 4607
rect 28224 4576 28273 4604
rect 28224 4564 28230 4576
rect 28261 4573 28273 4576
rect 28307 4604 28319 4607
rect 28994 4604 29000 4616
rect 28307 4576 29000 4604
rect 28307 4573 28319 4576
rect 28261 4567 28319 4573
rect 28994 4564 29000 4576
rect 29052 4604 29058 4616
rect 29825 4607 29883 4613
rect 29825 4604 29837 4607
rect 29052 4576 29837 4604
rect 29052 4564 29058 4576
rect 29825 4573 29837 4576
rect 29871 4573 29883 4607
rect 29825 4567 29883 4573
rect 30098 4564 30104 4616
rect 30156 4604 30162 4616
rect 32030 4604 32036 4616
rect 30156 4576 32036 4604
rect 30156 4564 30162 4576
rect 32030 4564 32036 4576
rect 32088 4604 32094 4616
rect 32140 4604 32168 4635
rect 32582 4632 32588 4644
rect 32640 4632 32646 4684
rect 33226 4632 33232 4684
rect 33284 4672 33290 4684
rect 33689 4675 33747 4681
rect 33689 4672 33701 4675
rect 33284 4644 33701 4672
rect 33284 4632 33290 4644
rect 33689 4641 33701 4644
rect 33735 4641 33747 4675
rect 33689 4635 33747 4641
rect 34606 4632 34612 4684
rect 34664 4672 34670 4684
rect 34736 4675 34794 4681
rect 34736 4672 34748 4675
rect 34664 4644 34748 4672
rect 34664 4632 34670 4644
rect 34736 4641 34748 4644
rect 34782 4641 34794 4675
rect 34736 4635 34794 4641
rect 32088 4576 32168 4604
rect 32088 4564 32094 4576
rect 23072 4508 24532 4536
rect 23072 4496 23078 4508
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 13786 4440 14197 4468
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 14185 4431 14243 4437
rect 14918 4428 14924 4480
rect 14976 4468 14982 4480
rect 18782 4468 18788 4480
rect 14976 4440 18788 4468
rect 14976 4428 14982 4440
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 34839 4471 34897 4477
rect 34839 4437 34851 4471
rect 34885 4468 34897 4471
rect 38562 4468 38568 4480
rect 34885 4440 38568 4468
rect 34885 4437 34897 4440
rect 34839 4431 34897 4437
rect 38562 4428 38568 4440
rect 38620 4428 38626 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 2409 4267 2467 4273
rect 2409 4233 2421 4267
rect 2455 4264 2467 4267
rect 2590 4264 2596 4276
rect 2455 4236 2596 4264
rect 2455 4233 2467 4236
rect 2409 4227 2467 4233
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 2777 4267 2835 4273
rect 2777 4264 2789 4267
rect 2740 4236 2789 4264
rect 2740 4224 2746 4236
rect 2777 4233 2789 4236
rect 2823 4233 2835 4267
rect 3050 4264 3056 4276
rect 3011 4236 3056 4264
rect 2777 4227 2835 4233
rect 3050 4224 3056 4236
rect 3108 4224 3114 4276
rect 3651 4267 3709 4273
rect 3651 4233 3663 4267
rect 3697 4264 3709 4267
rect 4246 4264 4252 4276
rect 3697 4236 4252 4264
rect 3697 4233 3709 4236
rect 3651 4227 3709 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5261 4267 5319 4273
rect 5261 4233 5273 4267
rect 5307 4264 5319 4267
rect 5626 4264 5632 4276
rect 5307 4236 5632 4264
rect 5307 4233 5319 4236
rect 5261 4227 5319 4233
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2568 4063 2626 4069
rect 1443 4032 2084 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2056 3933 2084 4032
rect 2568 4029 2580 4063
rect 2614 4060 2626 4063
rect 3068 4060 3096 4224
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 2614 4032 3096 4060
rect 3580 4063 3638 4069
rect 2614 4029 2626 4032
rect 2568 4023 2626 4029
rect 3580 4029 3592 4063
rect 3626 4060 3638 4063
rect 3988 4060 4016 4088
rect 5368 4069 5396 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 7006 4264 7012 4276
rect 6420 4236 7012 4264
rect 6420 4224 6426 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 8018 4264 8024 4276
rect 7979 4236 8024 4264
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12253 4267 12311 4273
rect 12253 4264 12265 4267
rect 11756 4236 12265 4264
rect 11756 4224 11762 4236
rect 12253 4233 12265 4236
rect 12299 4264 12311 4267
rect 12434 4264 12440 4276
rect 12299 4236 12440 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12434 4224 12440 4236
rect 12492 4264 12498 4276
rect 12492 4236 13032 4264
rect 12492 4224 12498 4236
rect 9953 4199 10011 4205
rect 9953 4196 9965 4199
rect 9863 4168 9965 4196
rect 9953 4165 9965 4168
rect 9999 4196 10011 4199
rect 10778 4196 10784 4208
rect 9999 4168 10784 4196
rect 9999 4165 10011 4168
rect 9953 4159 10011 4165
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8662 4128 8668 4140
rect 8619 4100 8668 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 3626 4032 4016 4060
rect 5353 4063 5411 4069
rect 3626 4029 3638 4032
rect 3580 4023 3638 4029
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5353 4023 5411 4029
rect 5534 4020 5540 4032
rect 5592 4060 5598 4072
rect 6086 4060 6092 4072
rect 5592 4032 6092 4060
rect 5592 4020 5598 4032
rect 6086 4020 6092 4032
rect 6144 4060 6150 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 6144 4032 6193 4060
rect 6144 4020 6150 4032
rect 6181 4029 6193 4032
rect 6227 4060 6239 4063
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6227 4032 6561 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 6549 4023 6607 4029
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7064 4032 7389 4060
rect 7064 4020 7070 4032
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 7742 4060 7748 4072
rect 7423 4032 7748 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9968 4060 9996 4159
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 12894 4156 12900 4208
rect 12952 4156 12958 4208
rect 13004 4196 13032 4236
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 13320 4236 13461 4264
rect 13320 4224 13326 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 17218 4264 17224 4276
rect 13449 4227 13507 4233
rect 13786 4236 17224 4264
rect 13786 4196 13814 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 17494 4264 17500 4276
rect 17455 4236 17500 4264
rect 17494 4224 17500 4236
rect 17552 4264 17558 4276
rect 18187 4267 18245 4273
rect 18187 4264 18199 4267
rect 17552 4236 18199 4264
rect 17552 4224 17558 4236
rect 18187 4233 18199 4236
rect 18233 4233 18245 4267
rect 18187 4227 18245 4233
rect 18322 4224 18328 4276
rect 18380 4264 18386 4276
rect 19199 4267 19257 4273
rect 19199 4264 19211 4267
rect 18380 4236 19211 4264
rect 18380 4224 18386 4236
rect 19199 4233 19211 4236
rect 19245 4233 19257 4267
rect 19794 4264 19800 4276
rect 19755 4236 19800 4264
rect 19199 4227 19257 4233
rect 19794 4224 19800 4236
rect 19852 4224 19858 4276
rect 21637 4267 21695 4273
rect 21637 4233 21649 4267
rect 21683 4264 21695 4267
rect 22370 4264 22376 4276
rect 21683 4236 22376 4264
rect 21683 4233 21695 4236
rect 21637 4227 21695 4233
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 23477 4267 23535 4273
rect 23477 4233 23489 4267
rect 23523 4264 23535 4267
rect 23799 4267 23857 4273
rect 23799 4264 23811 4267
rect 23523 4236 23811 4264
rect 23523 4233 23535 4236
rect 23477 4227 23535 4233
rect 23799 4233 23811 4236
rect 23845 4264 23857 4267
rect 24026 4264 24032 4276
rect 23845 4236 24032 4264
rect 23845 4233 23857 4236
rect 23799 4227 23857 4233
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 26418 4264 26424 4276
rect 26379 4236 26424 4264
rect 26418 4224 26424 4236
rect 26476 4224 26482 4276
rect 27614 4264 27620 4276
rect 27575 4236 27620 4264
rect 27614 4224 27620 4236
rect 27672 4224 27678 4276
rect 27890 4264 27896 4276
rect 27851 4236 27896 4264
rect 27890 4224 27896 4236
rect 27948 4224 27954 4276
rect 27982 4224 27988 4276
rect 28040 4264 28046 4276
rect 28215 4267 28273 4273
rect 28215 4264 28227 4267
rect 28040 4236 28227 4264
rect 28040 4224 28046 4236
rect 28215 4233 28227 4236
rect 28261 4233 28273 4267
rect 28994 4264 29000 4276
rect 28955 4236 29000 4264
rect 28215 4227 28273 4233
rect 28994 4224 29000 4236
rect 29052 4224 29058 4276
rect 34606 4224 34612 4276
rect 34664 4264 34670 4276
rect 35069 4267 35127 4273
rect 35069 4264 35081 4267
rect 34664 4236 35081 4264
rect 34664 4224 34670 4236
rect 35069 4233 35081 4236
rect 35115 4233 35127 4267
rect 35069 4227 35127 4233
rect 13004 4168 13814 4196
rect 14090 4156 14096 4208
rect 14148 4196 14154 4208
rect 15286 4196 15292 4208
rect 14148 4168 15292 4196
rect 14148 4156 14154 4168
rect 15286 4156 15292 4168
rect 15344 4196 15350 4208
rect 15381 4199 15439 4205
rect 15381 4196 15393 4199
rect 15344 4168 15393 4196
rect 15344 4156 15350 4168
rect 15381 4165 15393 4168
rect 15427 4165 15439 4199
rect 15381 4159 15439 4165
rect 15470 4156 15476 4208
rect 15528 4196 15534 4208
rect 16577 4199 16635 4205
rect 16577 4196 16589 4199
rect 15528 4168 16589 4196
rect 15528 4156 15534 4168
rect 16577 4165 16589 4168
rect 16623 4165 16635 4199
rect 16577 4159 16635 4165
rect 24670 4156 24676 4208
rect 24728 4196 24734 4208
rect 25406 4196 25412 4208
rect 24728 4168 25412 4196
rect 24728 4156 24734 4168
rect 25406 4156 25412 4168
rect 25464 4196 25470 4208
rect 25961 4199 26019 4205
rect 25961 4196 25973 4199
rect 25464 4168 25973 4196
rect 25464 4156 25470 4168
rect 25961 4165 25973 4168
rect 26007 4196 26019 4199
rect 26237 4199 26295 4205
rect 26237 4196 26249 4199
rect 26007 4168 26249 4196
rect 26007 4165 26019 4168
rect 25961 4159 26019 4165
rect 26237 4165 26249 4168
rect 26283 4165 26295 4199
rect 26436 4196 26464 4224
rect 28074 4196 28080 4208
rect 26436 4168 28080 4196
rect 26237 4159 26295 4165
rect 28074 4156 28080 4168
rect 28132 4156 28138 4208
rect 29457 4199 29515 4205
rect 29457 4165 29469 4199
rect 29503 4196 29515 4199
rect 29549 4199 29607 4205
rect 29549 4196 29561 4199
rect 29503 4168 29561 4196
rect 29503 4165 29515 4168
rect 29457 4159 29515 4165
rect 29549 4165 29561 4168
rect 29595 4165 29607 4199
rect 29549 4159 29607 4165
rect 11238 4128 11244 4140
rect 11199 4100 11244 4128
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 12912 4128 12940 4156
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12912 4100 13001 4128
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 13412 4100 14565 4128
rect 13412 4088 13418 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 16298 4128 16304 4140
rect 15068 4100 16160 4128
rect 16259 4100 16304 4128
rect 15068 4088 15074 4100
rect 12710 4060 12716 4072
rect 9539 4032 9996 4060
rect 12671 4032 12716 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 12897 4023 12955 4029
rect 5902 3992 5908 4004
rect 5863 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7190 3992 7196 4004
rect 7151 3964 7196 3992
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8894 3995 8952 4001
rect 8894 3992 8906 3995
rect 8435 3964 8906 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 8894 3961 8906 3964
rect 8940 3992 8952 3995
rect 9122 3992 9128 4004
rect 8940 3964 9128 3992
rect 8940 3961 8952 3964
rect 8894 3955 8952 3961
rect 9122 3952 9128 3964
rect 9180 3952 9186 4004
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3992 10379 3995
rect 10502 3992 10508 4004
rect 10367 3964 10508 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10502 3952 10508 3964
rect 10560 3992 10566 4004
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 10560 3964 10885 3992
rect 10560 3952 10566 3964
rect 10873 3961 10885 3964
rect 10919 3961 10931 3995
rect 10873 3955 10931 3961
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3961 11023 3995
rect 12912 3992 12940 4023
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 13909 3995 13967 4001
rect 13909 3992 13921 3995
rect 10965 3955 11023 3961
rect 12360 3964 13921 3992
rect 2041 3927 2099 3933
rect 2041 3893 2053 3927
rect 2087 3924 2099 3927
rect 2406 3924 2412 3936
rect 2087 3896 2412 3924
rect 2087 3893 2099 3896
rect 2041 3887 2099 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 7469 3927 7527 3933
rect 7469 3893 7481 3927
rect 7515 3924 7527 3927
rect 8294 3924 8300 3936
rect 7515 3896 8300 3924
rect 7515 3893 7527 3896
rect 7469 3887 7527 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 10980 3924 11008 3955
rect 12360 3936 12388 3964
rect 13909 3961 13921 3964
rect 13955 3992 13967 3995
rect 14476 3992 14504 4023
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 15565 4063 15623 4069
rect 15565 4060 15577 4063
rect 15344 4032 15577 4060
rect 15344 4020 15350 4032
rect 15565 4029 15577 4032
rect 15611 4029 15623 4063
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 15565 4023 15623 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16132 4060 16160 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 17221 4131 17279 4137
rect 17221 4097 17233 4131
rect 17267 4128 17279 4131
rect 17402 4128 17408 4140
rect 17267 4100 17408 4128
rect 17267 4097 17279 4100
rect 17221 4091 17279 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 18877 4131 18935 4137
rect 18877 4128 18889 4131
rect 18840 4100 18889 4128
rect 18840 4088 18846 4100
rect 18877 4097 18889 4100
rect 18923 4097 18935 4131
rect 21266 4128 21272 4140
rect 21227 4100 21272 4128
rect 18877 4091 18935 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 25498 4128 25504 4140
rect 25459 4100 25504 4128
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 30193 4131 30251 4137
rect 30193 4128 30205 4131
rect 25608 4100 30205 4128
rect 18116 4063 18174 4069
rect 18116 4060 18128 4063
rect 16132 4032 18128 4060
rect 18116 4029 18128 4032
rect 18162 4060 18174 4063
rect 19061 4063 19119 4069
rect 18162 4032 18644 4060
rect 18162 4029 18174 4032
rect 18116 4023 18174 4029
rect 15105 3995 15163 4001
rect 15105 3992 15117 3995
rect 13955 3964 15117 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 15105 3961 15117 3964
rect 15151 3992 15163 3995
rect 16040 3992 16068 4020
rect 15151 3964 16068 3992
rect 15151 3961 15163 3964
rect 15105 3955 15163 3961
rect 18616 3936 18644 4032
rect 19061 4029 19073 4063
rect 19107 4060 19119 4063
rect 19150 4060 19156 4072
rect 19107 4032 19156 4060
rect 19107 4029 19119 4032
rect 19061 4023 19119 4029
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 20772 4032 21465 4060
rect 20772 4020 20778 4032
rect 21453 4029 21465 4032
rect 21499 4060 21511 4063
rect 21913 4063 21971 4069
rect 21913 4060 21925 4063
rect 21499 4032 21925 4060
rect 21499 4029 21511 4032
rect 21453 4023 21511 4029
rect 21913 4029 21925 4032
rect 21959 4029 21971 4063
rect 21913 4023 21971 4029
rect 22462 4020 22468 4072
rect 22520 4060 22526 4072
rect 23728 4063 23786 4069
rect 23728 4060 23740 4063
rect 22520 4032 23740 4060
rect 22520 4020 22526 4032
rect 23728 4029 23740 4032
rect 23774 4060 23786 4063
rect 24854 4060 24860 4072
rect 23774 4032 24256 4060
rect 24767 4032 24860 4060
rect 23774 4029 23786 4032
rect 23728 4023 23786 4029
rect 24228 3936 24256 4032
rect 24854 4020 24860 4032
rect 24912 4060 24918 4072
rect 25225 4063 25283 4069
rect 25225 4060 25237 4063
rect 24912 4032 25237 4060
rect 24912 4020 24918 4032
rect 25225 4029 25237 4032
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 25240 3992 25268 4023
rect 25406 4020 25412 4072
rect 25464 4060 25470 4072
rect 25464 4032 25509 4060
rect 25464 4020 25470 4032
rect 25608 3992 25636 4100
rect 30193 4097 30205 4100
rect 30239 4128 30251 4131
rect 30466 4128 30472 4140
rect 30239 4100 30472 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 30466 4088 30472 4100
rect 30524 4128 30530 4140
rect 31386 4128 31392 4140
rect 30524 4100 30696 4128
rect 31347 4100 31392 4128
rect 30524 4088 30530 4100
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26513 4063 26571 4069
rect 26513 4060 26525 4063
rect 26384 4032 26525 4060
rect 26384 4020 26390 4032
rect 26513 4029 26525 4032
rect 26559 4029 26571 4063
rect 26513 4023 26571 4029
rect 26973 4063 27031 4069
rect 26973 4029 26985 4063
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 25240 3964 25636 3992
rect 26237 3995 26295 4001
rect 26237 3961 26249 3995
rect 26283 3992 26295 3995
rect 26988 3992 27016 4023
rect 27522 4020 27528 4072
rect 27580 4060 27586 4072
rect 28112 4063 28170 4069
rect 28112 4060 28124 4063
rect 27580 4032 28124 4060
rect 27580 4020 27586 4032
rect 28112 4029 28124 4032
rect 28158 4060 28170 4063
rect 28537 4063 28595 4069
rect 28537 4060 28549 4063
rect 28158 4032 28549 4060
rect 28158 4029 28170 4032
rect 28112 4023 28170 4029
rect 28537 4029 28549 4032
rect 28583 4029 28595 4063
rect 29270 4060 29276 4072
rect 29231 4032 29276 4060
rect 28537 4023 28595 4029
rect 26283 3964 27016 3992
rect 26283 3961 26295 3964
rect 26237 3955 26295 3961
rect 10652 3896 11008 3924
rect 11885 3927 11943 3933
rect 10652 3884 10658 3896
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12342 3924 12348 3936
rect 11931 3896 12348 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 18598 3924 18604 3936
rect 18559 3896 18604 3924
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 23106 3924 23112 3936
rect 23063 3896 23112 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 23106 3884 23112 3896
rect 23164 3924 23170 3936
rect 24026 3924 24032 3936
rect 23164 3896 24032 3924
rect 23164 3884 23170 3896
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24210 3924 24216 3936
rect 24171 3896 24216 3924
rect 24210 3884 24216 3896
rect 24268 3884 24274 3936
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 28552 3924 28580 4023
rect 29270 4020 29276 4032
rect 29328 4060 29334 4072
rect 30668 4069 30696 4100
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 31757 4131 31815 4137
rect 31757 4097 31769 4131
rect 31803 4128 31815 4131
rect 32125 4131 32183 4137
rect 32125 4128 32137 4131
rect 31803 4100 32137 4128
rect 31803 4097 31815 4100
rect 31757 4091 31815 4097
rect 32125 4097 32137 4100
rect 32171 4128 32183 4131
rect 32953 4131 33011 4137
rect 32171 4100 32628 4128
rect 32171 4097 32183 4100
rect 32125 4091 32183 4097
rect 29733 4063 29791 4069
rect 29733 4060 29745 4063
rect 29328 4032 29745 4060
rect 29328 4020 29334 4032
rect 29733 4029 29745 4032
rect 29779 4029 29791 4063
rect 29733 4023 29791 4029
rect 30653 4063 30711 4069
rect 30653 4029 30665 4063
rect 30699 4029 30711 4063
rect 30653 4023 30711 4029
rect 31205 4063 31263 4069
rect 31205 4029 31217 4063
rect 31251 4060 31263 4063
rect 31772 4060 31800 4091
rect 32600 4072 32628 4100
rect 32953 4097 32965 4131
rect 32999 4128 33011 4131
rect 33594 4128 33600 4140
rect 32999 4100 33600 4128
rect 32999 4097 33011 4100
rect 32953 4091 33011 4097
rect 33594 4088 33600 4100
rect 33652 4088 33658 4140
rect 31251 4032 31800 4060
rect 31251 4029 31263 4032
rect 31205 4023 31263 4029
rect 29549 3995 29607 4001
rect 29549 3961 29561 3995
rect 29595 3992 29607 3995
rect 30561 3995 30619 4001
rect 30561 3992 30573 3995
rect 29595 3964 30573 3992
rect 29595 3961 29607 3964
rect 29549 3955 29607 3961
rect 30561 3961 30573 3964
rect 30607 3992 30619 3995
rect 30926 3992 30932 4004
rect 30607 3964 30932 3992
rect 30607 3961 30619 3964
rect 30561 3955 30619 3961
rect 30926 3952 30932 3964
rect 30984 3992 30990 4004
rect 31220 3992 31248 4023
rect 32214 4020 32220 4072
rect 32272 4060 32278 4072
rect 32490 4060 32496 4072
rect 32272 4032 32496 4060
rect 32272 4020 32278 4032
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 32582 4020 32588 4072
rect 32640 4060 32646 4072
rect 32677 4063 32735 4069
rect 32677 4060 32689 4063
rect 32640 4032 32689 4060
rect 32640 4020 32646 4032
rect 32677 4029 32689 4032
rect 32723 4029 32735 4063
rect 32677 4023 32735 4029
rect 30984 3964 31248 3992
rect 30984 3952 30990 3964
rect 30466 3924 30472 3936
rect 28552 3896 30472 3924
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2685 3723 2743 3729
rect 2685 3689 2697 3723
rect 2731 3720 2743 3723
rect 2866 3720 2872 3732
rect 2731 3692 2872 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 5994 3720 6000 3732
rect 5955 3692 6000 3720
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6546 3720 6552 3732
rect 6507 3692 6552 3720
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 6914 3720 6920 3732
rect 6875 3692 6920 3720
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 10594 3720 10600 3732
rect 10555 3692 10600 3720
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 10744 3692 11345 3720
rect 10744 3680 10750 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 12158 3720 12164 3732
rect 12119 3692 12164 3720
rect 11333 3683 11391 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12860 3692 12909 3720
rect 12860 3680 12866 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13265 3723 13323 3729
rect 13265 3720 13277 3723
rect 13228 3692 13277 3720
rect 13228 3680 13234 3692
rect 13265 3689 13277 3692
rect 13311 3689 13323 3723
rect 13446 3720 13452 3732
rect 13407 3692 13452 3720
rect 13265 3683 13323 3689
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 15746 3720 15752 3732
rect 15703 3692 15752 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16022 3720 16028 3732
rect 15983 3692 16028 3720
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16899 3723 16957 3729
rect 16899 3720 16911 3723
rect 16540 3692 16911 3720
rect 16540 3680 16546 3692
rect 16899 3689 16911 3692
rect 16945 3689 16957 3723
rect 16899 3683 16957 3689
rect 17911 3723 17969 3729
rect 17911 3689 17923 3723
rect 17957 3720 17969 3723
rect 18874 3720 18880 3732
rect 17957 3692 18880 3720
rect 17957 3689 17969 3692
rect 17911 3683 17969 3689
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19150 3720 19156 3732
rect 19063 3692 19156 3720
rect 19150 3680 19156 3692
rect 19208 3720 19214 3732
rect 23014 3720 23020 3732
rect 19208 3692 23020 3720
rect 19208 3680 19214 3692
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 24029 3723 24087 3729
rect 24029 3689 24041 3723
rect 24075 3720 24087 3723
rect 24118 3720 24124 3732
rect 24075 3692 24124 3720
rect 24075 3689 24087 3692
rect 24029 3683 24087 3689
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 24670 3680 24676 3732
rect 24728 3720 24734 3732
rect 24949 3723 25007 3729
rect 24949 3720 24961 3723
rect 24728 3692 24961 3720
rect 24728 3680 24734 3692
rect 24949 3689 24961 3692
rect 24995 3689 25007 3723
rect 27982 3720 27988 3732
rect 27943 3692 27988 3720
rect 24949 3683 25007 3689
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 29825 3723 29883 3729
rect 29825 3689 29837 3723
rect 29871 3720 29883 3723
rect 29914 3720 29920 3732
rect 29871 3692 29920 3720
rect 29871 3689 29883 3692
rect 29825 3683 29883 3689
rect 29914 3680 29920 3692
rect 29972 3680 29978 3732
rect 32030 3680 32036 3732
rect 32088 3720 32094 3732
rect 32309 3723 32367 3729
rect 32309 3720 32321 3723
rect 32088 3692 32321 3720
rect 32088 3680 32094 3692
rect 32309 3689 32321 3692
rect 32355 3689 32367 3723
rect 32309 3683 32367 3689
rect 32490 3680 32496 3732
rect 32548 3720 32554 3732
rect 32677 3723 32735 3729
rect 32677 3720 32689 3723
rect 32548 3692 32689 3720
rect 32548 3680 32554 3692
rect 32677 3689 32689 3692
rect 32723 3689 32735 3723
rect 32677 3683 32735 3689
rect 2271 3655 2329 3661
rect 2271 3621 2283 3655
rect 2317 3652 2329 3655
rect 3602 3652 3608 3664
rect 2317 3624 3608 3652
rect 2317 3621 2329 3624
rect 2271 3615 2329 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 7742 3652 7748 3664
rect 7703 3624 7748 3652
rect 7742 3612 7748 3624
rect 7800 3652 7806 3664
rect 8478 3652 8484 3664
rect 7800 3624 8484 3652
rect 7800 3612 7806 3624
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 28810 3652 28816 3664
rect 24268 3624 28816 3652
rect 24268 3612 24274 3624
rect 28810 3612 28816 3624
rect 28868 3612 28874 3664
rect 31113 3655 31171 3661
rect 31113 3621 31125 3655
rect 31159 3652 31171 3655
rect 35434 3652 35440 3664
rect 31159 3624 35440 3652
rect 31159 3621 31171 3624
rect 31113 3615 31171 3621
rect 35434 3612 35440 3624
rect 35492 3612 35498 3664
rect 2184 3587 2242 3593
rect 2184 3553 2196 3587
rect 2230 3584 2242 3587
rect 2406 3584 2412 3596
rect 2230 3556 2412 3584
rect 2230 3553 2242 3556
rect 2184 3547 2242 3553
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 5902 3544 5908 3596
rect 5960 3584 5966 3596
rect 6362 3584 6368 3596
rect 5960 3556 6368 3584
rect 5960 3544 5966 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 10778 3584 10784 3596
rect 10739 3556 10784 3584
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12250 3584 12256 3596
rect 12207 3556 12256 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 15470 3584 15476 3596
rect 12400 3556 12445 3584
rect 15431 3556 15476 3584
rect 12400 3544 12406 3556
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15562 3544 15568 3596
rect 15620 3584 15626 3596
rect 16758 3584 16764 3596
rect 16816 3593 16822 3596
rect 16816 3587 16854 3593
rect 15620 3556 16764 3584
rect 15620 3544 15626 3556
rect 16758 3544 16764 3556
rect 16842 3584 16854 3587
rect 17808 3587 17866 3593
rect 17808 3584 17820 3587
rect 16842 3556 17820 3584
rect 16842 3553 16854 3556
rect 16816 3547 16854 3553
rect 17808 3553 17820 3556
rect 17854 3553 17866 3587
rect 17808 3547 17866 3553
rect 16816 3544 16822 3547
rect 28074 3544 28080 3596
rect 28132 3584 28138 3596
rect 30653 3587 30711 3593
rect 30653 3584 30665 3587
rect 28132 3556 30665 3584
rect 28132 3544 28138 3556
rect 30653 3553 30665 3556
rect 30699 3584 30711 3587
rect 30742 3584 30748 3596
rect 30699 3556 30748 3584
rect 30699 3553 30711 3556
rect 30653 3547 30711 3553
rect 30742 3544 30748 3556
rect 30800 3544 30806 3596
rect 30926 3584 30932 3596
rect 30887 3556 30932 3584
rect 30926 3544 30932 3556
rect 30984 3544 30990 3596
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7576 3488 8125 3516
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 7576 3457 7604 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 7432 3420 7573 3448
rect 7432 3408 7438 3420
rect 7561 3417 7573 3420
rect 7607 3417 7619 3451
rect 8018 3448 8024 3460
rect 7979 3420 8024 3448
rect 7561 3411 7619 3417
rect 8018 3408 8024 3420
rect 8076 3408 8082 3460
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 7883 3383 7941 3389
rect 7883 3380 7895 3383
rect 7340 3352 7895 3380
rect 7340 3340 7346 3352
rect 7883 3349 7895 3352
rect 7929 3349 7941 3383
rect 7883 3343 7941 3349
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 8168 3352 8217 3380
rect 8168 3340 8174 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 8205 3343 8263 3349
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 2406 3176 2412 3188
rect 2271 3148 2412 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7466 3176 7472 3188
rect 7331 3148 7472 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7392 2981 7420 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8076 3148 8217 3176
rect 8076 3136 8082 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8536 3148 8585 3176
rect 8536 3136 8542 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 8573 3139 8631 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10778 3176 10784 3188
rect 10551 3148 10784 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 12250 3176 12256 3188
rect 11563 3148 12256 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14139 3179 14197 3185
rect 14139 3176 14151 3179
rect 13136 3148 14151 3176
rect 13136 3136 13142 3148
rect 14139 3145 14151 3148
rect 14185 3145 14197 3179
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 14139 3139 14197 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15841 3179 15899 3185
rect 15841 3145 15853 3179
rect 15887 3176 15899 3179
rect 17678 3176 17684 3188
rect 15887 3148 17684 3176
rect 15887 3145 15899 3148
rect 15841 3139 15899 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 30742 3176 30748 3188
rect 30703 3148 30748 3176
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 10137 3111 10195 3117
rect 10137 3077 10149 3111
rect 10183 3108 10195 3111
rect 11054 3108 11060 3120
rect 10183 3080 11060 3108
rect 10183 3077 10195 3080
rect 10137 3071 10195 3077
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 9585 2975 9643 2981
rect 9585 2941 9597 2975
rect 9631 2972 9643 2975
rect 10152 2972 10180 3071
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 16758 3108 16764 3120
rect 16719 3080 16764 3108
rect 16758 3068 16764 3080
rect 16816 3108 16822 3120
rect 17773 3111 17831 3117
rect 17773 3108 17785 3111
rect 16816 3080 17785 3108
rect 16816 3068 16822 3080
rect 17773 3077 17785 3080
rect 17819 3077 17831 3111
rect 17773 3071 17831 3077
rect 30469 3111 30527 3117
rect 30469 3077 30481 3111
rect 30515 3108 30527 3111
rect 30926 3108 30932 3120
rect 30515 3080 30932 3108
rect 30515 3077 30527 3080
rect 30469 3071 30527 3077
rect 30926 3068 30932 3080
rect 30984 3068 30990 3120
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10560 3012 10609 3040
rect 10560 3000 10566 3012
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 10597 3003 10655 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 21266 3040 21272 3052
rect 14476 3012 21272 3040
rect 9631 2944 10180 2972
rect 12713 2975 12771 2981
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 12802 2972 12808 2984
rect 12759 2944 12808 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 14090 2981 14096 2984
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2941 12955 2975
rect 14036 2975 14096 2981
rect 14036 2972 14048 2975
rect 12897 2935 12955 2941
rect 14016 2941 14048 2972
rect 14082 2941 14096 2975
rect 14016 2935 14096 2941
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 7466 2904 7472 2916
rect 7340 2876 7472 2904
rect 7340 2864 7346 2876
rect 7466 2864 7472 2876
rect 7524 2904 7530 2916
rect 7837 2907 7895 2913
rect 7837 2904 7849 2907
rect 7524 2876 7849 2904
rect 7524 2864 7530 2876
rect 7837 2873 7849 2876
rect 7883 2904 7895 2907
rect 8202 2904 8208 2916
rect 7883 2876 8208 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 12342 2904 12348 2916
rect 12176 2876 12348 2904
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 6880 2808 7573 2836
rect 6880 2796 6886 2808
rect 7561 2805 7573 2808
rect 7607 2805 7619 2839
rect 7561 2799 7619 2805
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 12176 2845 12204 2876
rect 12342 2864 12348 2876
rect 12400 2904 12406 2916
rect 12912 2904 12940 2935
rect 12400 2876 12940 2904
rect 14016 2904 14044 2935
rect 14090 2932 14096 2935
rect 14148 2972 14154 2984
rect 14476 2981 14504 3012
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14148 2944 14473 2972
rect 14148 2932 14154 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 15344 2944 15669 2972
rect 15344 2932 15350 2944
rect 15657 2941 15669 2944
rect 15703 2972 15715 2975
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15703 2944 16129 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 14108 2904 14136 2932
rect 14016 2876 14136 2904
rect 12400 2864 12406 2876
rect 11793 2839 11851 2845
rect 11793 2836 11805 2839
rect 10468 2808 11805 2836
rect 10468 2796 10474 2808
rect 11793 2805 11805 2808
rect 11839 2836 11851 2839
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 11839 2808 12173 2836
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 12161 2805 12173 2808
rect 12207 2805 12219 2839
rect 12161 2799 12219 2805
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 7432 2604 7757 2632
rect 7432 2592 7438 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 10410 2632 10416 2644
rect 10371 2604 10416 2632
rect 7745 2595 7803 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11882 2632 11888 2644
rect 10827 2604 11888 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 10796 2496 10824 2595
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 14918 2632 14924 2644
rect 13311 2604 14924 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 10275 2468 10824 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11552 2499 11610 2505
rect 11552 2496 11564 2499
rect 11296 2468 11564 2496
rect 11296 2456 11302 2468
rect 11552 2465 11564 2468
rect 11598 2496 11610 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11598 2468 11989 2496
rect 11598 2465 11610 2468
rect 11552 2459 11610 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13280 2496 13308 2595
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 12667 2468 13308 2496
rect 28169 2499 28227 2505
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 28169 2465 28181 2499
rect 28215 2496 28227 2499
rect 28828 2496 28856 2592
rect 28215 2468 28856 2496
rect 28215 2465 28227 2468
rect 28169 2459 28227 2465
rect 28353 2363 28411 2369
rect 28353 2329 28365 2363
rect 28399 2360 28411 2363
rect 29638 2360 29644 2372
rect 28399 2332 29644 2360
rect 28399 2329 28411 2332
rect 28353 2323 28411 2329
rect 29638 2320 29644 2332
rect 29696 2320 29702 2372
rect 11655 2295 11713 2301
rect 11655 2261 11667 2295
rect 11701 2292 11713 2295
rect 11882 2292 11888 2304
rect 11701 2264 11888 2292
rect 11701 2261 11713 2264
rect 11655 2255 11713 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12894 2292 12900 2304
rect 12851 2264 12900 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 2498 280 2504 332
rect 2556 320 2562 332
rect 7006 320 7012 332
rect 2556 292 7012 320
rect 2556 280 2562 292
rect 7006 280 7012 292
rect 7064 280 7070 332
rect 15654 76 15660 128
rect 15712 116 15718 128
rect 20622 116 20628 128
rect 15712 88 20628 116
rect 15712 76 15718 88
rect 20622 76 20628 88
rect 20680 76 20686 128
<< via1 >>
rect 11152 15580 11204 15632
rect 19156 15580 19208 15632
rect 15476 15512 15528 15564
rect 16212 15512 16264 15564
rect 27988 15512 28040 15564
rect 28724 15512 28776 15564
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 20812 13336 20864 13388
rect 11888 13268 11940 13320
rect 20444 13268 20496 13320
rect 112 13132 164 13184
rect 12348 13132 12400 13184
rect 15844 13132 15896 13184
rect 20076 13132 20128 13184
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 7196 12928 7248 12980
rect 13360 12928 13412 12980
rect 23756 12928 23808 12980
rect 25780 12928 25832 12980
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 35900 12860 35952 12912
rect 2780 12724 2832 12776
rect 13268 12792 13320 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 3148 12588 3200 12640
rect 8668 12588 8720 12640
rect 10416 12724 10468 12776
rect 13360 12724 13412 12776
rect 24492 12792 24544 12844
rect 15844 12656 15896 12708
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 15752 12588 15804 12640
rect 20444 12767 20496 12776
rect 20444 12733 20453 12767
rect 20453 12733 20487 12767
rect 20487 12733 20496 12767
rect 20444 12724 20496 12733
rect 21456 12724 21508 12776
rect 20720 12699 20772 12708
rect 20720 12665 20729 12699
rect 20729 12665 20763 12699
rect 20763 12665 20772 12699
rect 20720 12656 20772 12665
rect 24400 12724 24452 12776
rect 32772 12792 32824 12844
rect 33876 12724 33928 12776
rect 31300 12656 31352 12708
rect 18236 12588 18288 12640
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 19800 12588 19852 12597
rect 20812 12588 20864 12640
rect 26424 12588 26476 12640
rect 29092 12631 29144 12640
rect 29092 12597 29101 12631
rect 29101 12597 29135 12631
rect 29135 12597 29144 12631
rect 29092 12588 29144 12597
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 15568 12384 15620 12436
rect 18788 12384 18840 12436
rect 23296 12384 23348 12436
rect 20 12316 72 12368
rect 16212 12359 16264 12368
rect 16212 12325 16221 12359
rect 16221 12325 16255 12359
rect 16255 12325 16264 12359
rect 16212 12316 16264 12325
rect 21272 12316 21324 12368
rect 26332 12316 26384 12368
rect 29092 12316 29144 12368
rect 2320 12248 2372 12300
rect 3424 12248 3476 12300
rect 4988 12248 5040 12300
rect 6552 12291 6604 12300
rect 6552 12257 6561 12291
rect 6561 12257 6595 12291
rect 6595 12257 6604 12291
rect 6552 12248 6604 12257
rect 7472 12248 7524 12300
rect 10968 12291 11020 12300
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 10600 12112 10652 12164
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 19524 12248 19576 12300
rect 22284 12248 22336 12300
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 27436 12248 27488 12300
rect 28080 12248 28132 12300
rect 33600 12248 33652 12300
rect 35348 12248 35400 12300
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 21272 12180 21324 12232
rect 16488 12112 16540 12164
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 16672 12112 16724 12121
rect 21916 12112 21968 12164
rect 2228 12044 2280 12096
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 8116 12044 8168 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 13452 12044 13504 12096
rect 19800 12044 19852 12096
rect 21732 12044 21784 12096
rect 22928 12044 22980 12096
rect 24676 12087 24728 12096
rect 24676 12053 24685 12087
rect 24685 12053 24719 12087
rect 24719 12053 24728 12087
rect 24676 12044 24728 12053
rect 25320 12087 25372 12096
rect 25320 12053 25329 12087
rect 25329 12053 25363 12087
rect 25363 12053 25372 12087
rect 25320 12044 25372 12053
rect 26516 12044 26568 12096
rect 29000 12044 29052 12096
rect 34704 12044 34756 12096
rect 36544 12044 36596 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 15844 11840 15896 11892
rect 16212 11840 16264 11892
rect 21272 11840 21324 11892
rect 24492 11883 24544 11892
rect 2044 11815 2096 11824
rect 2044 11781 2053 11815
rect 2053 11781 2087 11815
rect 2087 11781 2096 11815
rect 2044 11772 2096 11781
rect 2320 11772 2372 11824
rect 2872 11772 2924 11824
rect 3700 11772 3752 11824
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 8576 11704 8628 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 10416 11704 10468 11756
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2320 11636 2372 11688
rect 2872 11500 2924 11552
rect 3792 11636 3844 11688
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 4436 11636 4488 11688
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 4620 11568 4672 11620
rect 6552 11611 6604 11620
rect 6552 11577 6561 11611
rect 6561 11577 6595 11611
rect 6595 11577 6604 11611
rect 6552 11568 6604 11577
rect 8300 11611 8352 11620
rect 8300 11577 8309 11611
rect 8309 11577 8343 11611
rect 8343 11577 8352 11611
rect 8300 11568 8352 11577
rect 3516 11500 3568 11509
rect 4068 11500 4120 11552
rect 4988 11500 5040 11552
rect 5264 11543 5316 11552
rect 5264 11509 5273 11543
rect 5273 11509 5307 11543
rect 5307 11509 5316 11543
rect 5264 11500 5316 11509
rect 5816 11500 5868 11552
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 7472 11500 7524 11509
rect 8944 11500 8996 11552
rect 11152 11636 11204 11688
rect 12808 11772 12860 11824
rect 13084 11772 13136 11824
rect 13728 11772 13780 11824
rect 16672 11772 16724 11824
rect 12072 11704 12124 11756
rect 19248 11704 19300 11756
rect 11520 11611 11572 11620
rect 11520 11577 11529 11611
rect 11529 11577 11563 11611
rect 11563 11577 11572 11611
rect 11520 11568 11572 11577
rect 12532 11611 12584 11620
rect 12532 11577 12541 11611
rect 12541 11577 12575 11611
rect 12575 11577 12584 11611
rect 12532 11568 12584 11577
rect 12624 11611 12676 11620
rect 12624 11577 12633 11611
rect 12633 11577 12667 11611
rect 12667 11577 12676 11611
rect 13176 11611 13228 11620
rect 12624 11568 12676 11577
rect 13176 11577 13185 11611
rect 13185 11577 13219 11611
rect 13219 11577 13228 11611
rect 13176 11568 13228 11577
rect 10968 11500 11020 11552
rect 14924 11636 14976 11688
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 17684 11636 17736 11688
rect 19524 11679 19576 11688
rect 19524 11645 19533 11679
rect 19533 11645 19567 11679
rect 19567 11645 19576 11679
rect 19524 11636 19576 11645
rect 20444 11704 20496 11756
rect 24492 11849 24501 11883
rect 24501 11849 24535 11883
rect 24535 11849 24544 11883
rect 24492 11840 24544 11849
rect 30104 11840 30156 11892
rect 31300 11883 31352 11892
rect 31300 11849 31309 11883
rect 31309 11849 31343 11883
rect 31343 11849 31352 11883
rect 31300 11840 31352 11849
rect 33600 11883 33652 11892
rect 33600 11849 33609 11883
rect 33609 11849 33643 11883
rect 33643 11849 33652 11883
rect 33600 11840 33652 11849
rect 35716 11840 35768 11892
rect 25136 11772 25188 11824
rect 27988 11772 28040 11824
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 32128 11704 32180 11756
rect 16304 11611 16356 11620
rect 16304 11577 16313 11611
rect 16313 11577 16347 11611
rect 16347 11577 16356 11611
rect 16304 11568 16356 11577
rect 16488 11568 16540 11620
rect 15016 11500 15068 11552
rect 16120 11500 16172 11552
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 24492 11636 24544 11688
rect 24768 11636 24820 11688
rect 26056 11679 26108 11688
rect 26056 11645 26065 11679
rect 26065 11645 26099 11679
rect 26099 11645 26108 11679
rect 26056 11636 26108 11645
rect 26700 11679 26752 11688
rect 20444 11611 20496 11620
rect 20444 11577 20453 11611
rect 20453 11577 20487 11611
rect 20487 11577 20496 11611
rect 20444 11568 20496 11577
rect 21548 11568 21600 11620
rect 22008 11611 22060 11620
rect 22008 11577 22017 11611
rect 22017 11577 22051 11611
rect 22051 11577 22060 11611
rect 22008 11568 22060 11577
rect 22100 11568 22152 11620
rect 23020 11611 23072 11620
rect 23020 11577 23029 11611
rect 23029 11577 23063 11611
rect 23063 11577 23072 11611
rect 23020 11568 23072 11577
rect 25412 11611 25464 11620
rect 25412 11577 25421 11611
rect 25421 11577 25455 11611
rect 25455 11577 25464 11611
rect 25412 11568 25464 11577
rect 26700 11645 26709 11679
rect 26709 11645 26743 11679
rect 26743 11645 26752 11679
rect 26700 11636 26752 11645
rect 31300 11636 31352 11688
rect 33968 11636 34020 11688
rect 35164 11636 35216 11688
rect 19800 11500 19852 11552
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 23204 11500 23256 11552
rect 26608 11568 26660 11620
rect 26976 11611 27028 11620
rect 26976 11577 26985 11611
rect 26985 11577 27019 11611
rect 27019 11577 27028 11611
rect 26976 11568 27028 11577
rect 27436 11500 27488 11552
rect 27528 11500 27580 11552
rect 28080 11500 28132 11552
rect 31116 11500 31168 11552
rect 31760 11543 31812 11552
rect 31760 11509 31769 11543
rect 31769 11509 31803 11543
rect 31803 11509 31812 11543
rect 31760 11500 31812 11509
rect 32772 11500 32824 11552
rect 33600 11500 33652 11552
rect 34152 11500 34204 11552
rect 35348 11500 35400 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 3700 11339 3752 11348
rect 3700 11305 3709 11339
rect 3709 11305 3743 11339
rect 3743 11305 3752 11339
rect 3700 11296 3752 11305
rect 4252 11296 4304 11348
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 9220 11339 9272 11348
rect 7656 11296 7708 11305
rect 8116 11271 8168 11280
rect 8116 11237 8125 11271
rect 8125 11237 8159 11271
rect 8159 11237 8168 11271
rect 8116 11228 8168 11237
rect 9220 11305 9229 11339
rect 9229 11305 9263 11339
rect 9263 11305 9272 11339
rect 9220 11296 9272 11305
rect 12532 11296 12584 11348
rect 8944 11228 8996 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 11980 11271 12032 11280
rect 11980 11237 11989 11271
rect 11989 11237 12023 11271
rect 12023 11237 12032 11271
rect 11980 11228 12032 11237
rect 13544 11271 13596 11280
rect 13544 11237 13553 11271
rect 13553 11237 13587 11271
rect 13587 11237 13596 11271
rect 13544 11228 13596 11237
rect 16212 11228 16264 11280
rect 18696 11296 18748 11348
rect 18236 11271 18288 11280
rect 18236 11237 18245 11271
rect 18245 11237 18279 11271
rect 18279 11237 18288 11271
rect 18236 11228 18288 11237
rect 19156 11296 19208 11348
rect 20536 11296 20588 11348
rect 21640 11228 21692 11280
rect 1768 11160 1820 11212
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2228 11203 2280 11212
rect 2044 11160 2096 11169
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4436 11160 4488 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 15292 11160 15344 11212
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 27988 11296 28040 11348
rect 30380 11339 30432 11348
rect 30380 11305 30389 11339
rect 30389 11305 30423 11339
rect 30423 11305 30432 11339
rect 30380 11296 30432 11305
rect 33324 11296 33376 11348
rect 26240 11271 26292 11280
rect 26240 11237 26249 11271
rect 26249 11237 26283 11271
rect 26283 11237 26292 11271
rect 26240 11228 26292 11237
rect 26424 11228 26476 11280
rect 26700 11271 26752 11280
rect 26700 11237 26709 11271
rect 26709 11237 26743 11271
rect 26743 11237 26752 11271
rect 26700 11228 26752 11237
rect 30840 11228 30892 11280
rect 34152 11228 34204 11280
rect 34612 11228 34664 11280
rect 1400 11092 1452 11144
rect 2504 11092 2556 11144
rect 8484 11092 8536 11144
rect 10140 11092 10192 11144
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 13636 11092 13688 11144
rect 16580 11135 16632 11144
rect 4252 11024 4304 11076
rect 13176 11024 13228 11076
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 19064 11092 19116 11144
rect 19524 11024 19576 11076
rect 21824 11135 21876 11144
rect 21824 11101 21833 11135
rect 21833 11101 21867 11135
rect 21867 11101 21876 11135
rect 21824 11092 21876 11101
rect 22008 11092 22060 11144
rect 23020 11092 23072 11144
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 2872 10956 2924 11008
rect 4896 10956 4948 11008
rect 10968 10956 11020 11008
rect 11152 10999 11204 11008
rect 11152 10965 11161 10999
rect 11161 10965 11195 10999
rect 11195 10965 11204 10999
rect 11152 10956 11204 10965
rect 15844 10956 15896 11008
rect 21548 10956 21600 11008
rect 23296 11160 23348 11212
rect 23940 11160 23992 11212
rect 24768 11203 24820 11212
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 28172 11160 28224 11212
rect 30104 11203 30156 11212
rect 30104 11169 30113 11203
rect 30113 11169 30147 11203
rect 30147 11169 30156 11203
rect 30104 11160 30156 11169
rect 32128 11203 32180 11212
rect 26608 11092 26660 11144
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 29000 11092 29052 11144
rect 32128 11169 32137 11203
rect 32137 11169 32171 11203
rect 32171 11169 32180 11203
rect 32128 11160 32180 11169
rect 35992 11160 36044 11212
rect 31024 11092 31076 11144
rect 26240 11024 26292 11076
rect 31392 11024 31444 11076
rect 34980 11067 35032 11076
rect 34980 11033 34989 11067
rect 34989 11033 35023 11067
rect 35023 11033 35032 11067
rect 34980 11024 35032 11033
rect 23572 10956 23624 11008
rect 25780 10999 25832 11008
rect 25780 10965 25789 10999
rect 25789 10965 25823 10999
rect 25823 10965 25832 10999
rect 25780 10956 25832 10965
rect 29828 10999 29880 11008
rect 29828 10965 29837 10999
rect 29837 10965 29871 10999
rect 29871 10965 29880 10999
rect 29828 10956 29880 10965
rect 32956 10956 33008 11008
rect 35072 10956 35124 11008
rect 35808 10956 35860 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 2044 10752 2096 10804
rect 4436 10795 4488 10804
rect 4436 10761 4445 10795
rect 4445 10761 4479 10795
rect 4479 10761 4488 10795
rect 4436 10752 4488 10761
rect 6920 10752 6972 10804
rect 8300 10752 8352 10804
rect 1584 10684 1636 10736
rect 2964 10727 3016 10736
rect 2964 10693 2973 10727
rect 2973 10693 3007 10727
rect 3007 10693 3016 10727
rect 2964 10684 3016 10693
rect 3976 10684 4028 10736
rect 4988 10684 5040 10736
rect 6736 10684 6788 10736
rect 8024 10684 8076 10736
rect 8944 10727 8996 10736
rect 8944 10693 8953 10727
rect 8953 10693 8987 10727
rect 8987 10693 8996 10727
rect 8944 10684 8996 10693
rect 1676 10548 1728 10600
rect 2136 10548 2188 10600
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 3516 10616 3568 10668
rect 4620 10616 4672 10668
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 5264 10616 5316 10668
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 4896 10523 4948 10532
rect 4896 10489 4905 10523
rect 4905 10489 4939 10523
rect 4939 10489 4948 10523
rect 4896 10480 4948 10489
rect 112 10412 164 10464
rect 1768 10412 1820 10464
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 7012 10412 7064 10464
rect 7932 10480 7984 10532
rect 9864 10752 9916 10804
rect 13544 10752 13596 10804
rect 16120 10752 16172 10804
rect 16212 10752 16264 10804
rect 18236 10752 18288 10804
rect 19064 10795 19116 10804
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 21824 10752 21876 10804
rect 25228 10752 25280 10804
rect 26884 10752 26936 10804
rect 31024 10795 31076 10804
rect 10140 10727 10192 10736
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 13728 10684 13780 10736
rect 15292 10727 15344 10736
rect 15292 10693 15301 10727
rect 15301 10693 15335 10727
rect 15335 10693 15344 10727
rect 18696 10727 18748 10736
rect 15292 10684 15344 10693
rect 10600 10616 10652 10668
rect 11520 10616 11572 10668
rect 12532 10616 12584 10668
rect 14188 10616 14240 10668
rect 18696 10693 18705 10727
rect 18705 10693 18739 10727
rect 18739 10693 18748 10727
rect 18696 10684 18748 10693
rect 19524 10727 19576 10736
rect 19524 10693 19533 10727
rect 19533 10693 19567 10727
rect 19567 10693 19576 10727
rect 19524 10684 19576 10693
rect 20444 10616 20496 10668
rect 23572 10616 23624 10668
rect 25228 10616 25280 10668
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 31024 10761 31033 10795
rect 31033 10761 31067 10795
rect 31067 10761 31076 10795
rect 31024 10752 31076 10761
rect 31116 10752 31168 10804
rect 32864 10752 32916 10804
rect 33968 10752 34020 10804
rect 32128 10684 32180 10736
rect 33508 10684 33560 10736
rect 28448 10616 28500 10668
rect 29828 10659 29880 10668
rect 29828 10625 29837 10659
rect 29837 10625 29871 10659
rect 29871 10625 29880 10659
rect 29828 10616 29880 10625
rect 31760 10616 31812 10668
rect 35164 10684 35216 10736
rect 34980 10659 35032 10668
rect 34980 10625 34989 10659
rect 34989 10625 35023 10659
rect 35023 10625 35032 10659
rect 34980 10616 35032 10625
rect 10232 10548 10284 10600
rect 13636 10548 13688 10600
rect 11980 10480 12032 10532
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 9864 10412 9916 10464
rect 10600 10412 10652 10464
rect 11336 10412 11388 10464
rect 16304 10548 16356 10600
rect 15844 10480 15896 10532
rect 14740 10412 14792 10464
rect 21456 10548 21508 10600
rect 22376 10548 22428 10600
rect 23940 10591 23992 10600
rect 23940 10557 23949 10591
rect 23949 10557 23983 10591
rect 23983 10557 23992 10591
rect 23940 10548 23992 10557
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 18144 10523 18196 10532
rect 18144 10489 18153 10523
rect 18153 10489 18187 10523
rect 18187 10489 18196 10523
rect 18144 10480 18196 10489
rect 21272 10480 21324 10532
rect 24860 10523 24912 10532
rect 24860 10489 24869 10523
rect 24869 10489 24903 10523
rect 24903 10489 24912 10523
rect 24860 10480 24912 10489
rect 24952 10480 25004 10532
rect 25780 10523 25832 10532
rect 25780 10489 25789 10523
rect 25789 10489 25823 10523
rect 25823 10489 25832 10523
rect 25780 10480 25832 10489
rect 32404 10548 32456 10600
rect 39580 10752 39632 10804
rect 37924 10659 37976 10668
rect 37924 10625 37933 10659
rect 37933 10625 37967 10659
rect 37967 10625 37976 10659
rect 37924 10616 37976 10625
rect 21640 10412 21692 10464
rect 24768 10412 24820 10464
rect 25320 10412 25372 10464
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 26700 10455 26752 10464
rect 25596 10412 25648 10421
rect 26700 10421 26709 10455
rect 26709 10421 26743 10455
rect 26743 10421 26752 10455
rect 26700 10412 26752 10421
rect 28172 10412 28224 10464
rect 31668 10480 31720 10532
rect 32496 10480 32548 10532
rect 33416 10480 33468 10532
rect 34612 10480 34664 10532
rect 35072 10523 35124 10532
rect 35072 10489 35081 10523
rect 35081 10489 35115 10523
rect 35115 10489 35124 10523
rect 35072 10480 35124 10489
rect 35992 10523 36044 10532
rect 35992 10489 36001 10523
rect 36001 10489 36035 10523
rect 36035 10489 36044 10523
rect 35992 10480 36044 10489
rect 36084 10480 36136 10532
rect 30656 10412 30708 10464
rect 33140 10412 33192 10464
rect 33508 10412 33560 10464
rect 35256 10412 35308 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 4896 10208 4948 10260
rect 7104 10208 7156 10260
rect 7748 10208 7800 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8116 10208 8168 10260
rect 10140 10208 10192 10260
rect 10600 10208 10652 10260
rect 2228 10140 2280 10192
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 4712 10072 4764 10124
rect 8944 10072 8996 10124
rect 9036 10072 9088 10124
rect 11060 10208 11112 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11980 10208 12032 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 12624 10208 12676 10260
rect 15844 10251 15896 10260
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 16304 10208 16356 10260
rect 16580 10208 16632 10260
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 18144 10208 18196 10260
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 20444 10208 20496 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 24124 10251 24176 10260
rect 24124 10217 24133 10251
rect 24133 10217 24167 10251
rect 24167 10217 24176 10251
rect 24124 10208 24176 10217
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 26424 10208 26476 10260
rect 26516 10208 26568 10260
rect 12992 10183 13044 10192
rect 12992 10149 13001 10183
rect 13001 10149 13035 10183
rect 13035 10149 13044 10183
rect 12992 10140 13044 10149
rect 22836 10183 22888 10192
rect 22836 10149 22845 10183
rect 22845 10149 22879 10183
rect 22879 10149 22888 10183
rect 22836 10140 22888 10149
rect 25044 10183 25096 10192
rect 25044 10149 25053 10183
rect 25053 10149 25087 10183
rect 25087 10149 25096 10183
rect 25044 10140 25096 10149
rect 27344 10208 27396 10260
rect 30104 10251 30156 10260
rect 30104 10217 30113 10251
rect 30113 10217 30147 10251
rect 30147 10217 30156 10251
rect 30104 10208 30156 10217
rect 30656 10251 30708 10260
rect 30656 10217 30665 10251
rect 30665 10217 30699 10251
rect 30699 10217 30708 10251
rect 30656 10208 30708 10217
rect 31668 10251 31720 10260
rect 31668 10217 31677 10251
rect 31677 10217 31711 10251
rect 31711 10217 31720 10251
rect 31668 10208 31720 10217
rect 34152 10208 34204 10260
rect 34704 10208 34756 10260
rect 26700 10183 26752 10192
rect 26700 10149 26709 10183
rect 26709 10149 26743 10183
rect 26743 10149 26752 10183
rect 28264 10183 28316 10192
rect 26700 10140 26752 10149
rect 28264 10149 28273 10183
rect 28273 10149 28307 10183
rect 28307 10149 28316 10183
rect 28264 10140 28316 10149
rect 33416 10140 33468 10192
rect 34612 10183 34664 10192
rect 34612 10149 34621 10183
rect 34621 10149 34655 10183
rect 34655 10149 34664 10183
rect 34612 10140 34664 10149
rect 35164 10183 35216 10192
rect 35164 10149 35173 10183
rect 35173 10149 35207 10183
rect 35207 10149 35216 10183
rect 35164 10140 35216 10149
rect 36084 10183 36136 10192
rect 36084 10149 36093 10183
rect 36093 10149 36127 10183
rect 36127 10149 36136 10183
rect 36084 10140 36136 10149
rect 36176 10183 36228 10192
rect 36176 10149 36185 10183
rect 36185 10149 36219 10183
rect 36219 10149 36228 10183
rect 36176 10140 36228 10149
rect 11888 10072 11940 10124
rect 18236 10072 18288 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 7472 10004 7524 10056
rect 11520 10004 11572 10056
rect 15200 10004 15252 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 19064 10004 19116 10056
rect 19248 10004 19300 10056
rect 20720 10072 20772 10124
rect 21916 10072 21968 10124
rect 30380 10072 30432 10124
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 25228 10047 25280 10056
rect 24768 9936 24820 9988
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 27988 10004 28040 10056
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 32956 10047 33008 10056
rect 32956 10013 32965 10047
rect 32965 10013 32999 10047
rect 32999 10013 33008 10047
rect 32956 10004 33008 10013
rect 34888 10004 34940 10056
rect 34980 10004 35032 10056
rect 25872 9936 25924 9988
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 10968 9868 11020 9920
rect 13728 9868 13780 9920
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 16672 9868 16724 9877
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 23388 9868 23440 9920
rect 24124 9868 24176 9920
rect 31208 9911 31260 9920
rect 31208 9877 31217 9911
rect 31217 9877 31251 9911
rect 31251 9877 31260 9911
rect 31208 9868 31260 9877
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 2136 9596 2188 9648
rect 1676 9528 1728 9580
rect 4896 9528 4948 9580
rect 5172 9460 5224 9512
rect 3516 9392 3568 9444
rect 6920 9460 6972 9512
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 8208 9528 8260 9580
rect 10232 9664 10284 9716
rect 9956 9596 10008 9648
rect 8576 9503 8628 9512
rect 7380 9392 7432 9444
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 11336 9528 11388 9580
rect 12992 9664 13044 9716
rect 15844 9664 15896 9716
rect 17592 9664 17644 9716
rect 18788 9664 18840 9716
rect 21640 9707 21692 9716
rect 21640 9673 21649 9707
rect 21649 9673 21683 9707
rect 21683 9673 21692 9707
rect 21640 9664 21692 9673
rect 21916 9707 21968 9716
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 22744 9664 22796 9716
rect 22836 9664 22888 9716
rect 24952 9664 25004 9716
rect 25044 9664 25096 9716
rect 28264 9664 28316 9716
rect 29000 9707 29052 9716
rect 29000 9673 29009 9707
rect 29009 9673 29043 9707
rect 29043 9673 29052 9707
rect 29000 9664 29052 9673
rect 31208 9664 31260 9716
rect 34612 9664 34664 9716
rect 36176 9664 36228 9716
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 10968 9460 11020 9512
rect 13728 9596 13780 9648
rect 14188 9528 14240 9580
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 18420 9596 18472 9648
rect 19340 9639 19392 9648
rect 19340 9605 19349 9639
rect 19349 9605 19383 9639
rect 19383 9605 19392 9639
rect 19340 9596 19392 9605
rect 17224 9528 17276 9580
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 19984 9528 20036 9580
rect 21456 9528 21508 9580
rect 23664 9596 23716 9648
rect 24400 9639 24452 9648
rect 24400 9605 24409 9639
rect 24409 9605 24443 9639
rect 24443 9605 24452 9639
rect 24400 9596 24452 9605
rect 26700 9596 26752 9648
rect 27988 9596 28040 9648
rect 24584 9528 24636 9580
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 26608 9571 26660 9580
rect 26608 9537 26617 9571
rect 26617 9537 26651 9571
rect 26651 9537 26660 9571
rect 26608 9528 26660 9537
rect 35072 9596 35124 9648
rect 29828 9571 29880 9580
rect 13360 9460 13412 9469
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 2596 9324 2648 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 7012 9367 7064 9376
rect 4712 9324 4764 9333
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 7104 9324 7156 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 9772 9324 9824 9376
rect 12164 9392 12216 9444
rect 10876 9324 10928 9376
rect 10968 9324 11020 9376
rect 11336 9324 11388 9376
rect 11520 9324 11572 9376
rect 14096 9392 14148 9444
rect 15384 9460 15436 9512
rect 16672 9460 16724 9512
rect 16028 9392 16080 9444
rect 18144 9435 18196 9444
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 18420 9392 18472 9444
rect 21272 9392 21324 9444
rect 14004 9324 14056 9376
rect 14648 9324 14700 9376
rect 19340 9324 19392 9376
rect 24400 9460 24452 9512
rect 27344 9460 27396 9512
rect 29276 9503 29328 9512
rect 29276 9469 29285 9503
rect 29285 9469 29319 9503
rect 29319 9469 29328 9503
rect 29276 9460 29328 9469
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 32864 9528 32916 9580
rect 34980 9528 35032 9580
rect 36544 9571 36596 9580
rect 36544 9537 36553 9571
rect 36553 9537 36587 9571
rect 36587 9537 36596 9571
rect 36544 9528 36596 9537
rect 31484 9460 31536 9512
rect 24768 9392 24820 9444
rect 23112 9367 23164 9376
rect 23112 9333 23121 9367
rect 23121 9333 23155 9367
rect 23155 9333 23164 9367
rect 23112 9324 23164 9333
rect 25044 9324 25096 9376
rect 26516 9367 26568 9376
rect 26516 9333 26525 9367
rect 26525 9333 26559 9367
rect 26559 9333 26568 9367
rect 30656 9392 30708 9444
rect 31576 9392 31628 9444
rect 26516 9324 26568 9333
rect 32312 9324 32364 9376
rect 32496 9324 32548 9376
rect 33692 9435 33744 9444
rect 33692 9401 33701 9435
rect 33701 9401 33735 9435
rect 33735 9401 33744 9435
rect 33692 9392 33744 9401
rect 34796 9392 34848 9444
rect 34428 9324 34480 9376
rect 34520 9324 34572 9376
rect 36636 9435 36688 9444
rect 36636 9401 36645 9435
rect 36645 9401 36679 9435
rect 36679 9401 36688 9435
rect 37188 9435 37240 9444
rect 36636 9392 36688 9401
rect 37188 9401 37197 9435
rect 37197 9401 37231 9435
rect 37231 9401 37240 9435
rect 37188 9392 37240 9401
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1676 9120 1728 9172
rect 3976 9120 4028 9172
rect 7472 9120 7524 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 10692 9120 10744 9172
rect 13360 9120 13412 9172
rect 14648 9120 14700 9172
rect 21456 9163 21508 9172
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 24216 9120 24268 9172
rect 24860 9120 24912 9172
rect 25044 9163 25096 9172
rect 25044 9129 25053 9163
rect 25053 9129 25087 9163
rect 25087 9129 25096 9163
rect 25044 9120 25096 9129
rect 25596 9163 25648 9172
rect 25596 9129 25605 9163
rect 25605 9129 25639 9163
rect 25639 9129 25648 9163
rect 25596 9120 25648 9129
rect 25872 9163 25924 9172
rect 25872 9129 25881 9163
rect 25881 9129 25915 9163
rect 25915 9129 25924 9163
rect 25872 9120 25924 9129
rect 26700 9120 26752 9172
rect 26976 9120 27028 9172
rect 29276 9163 29328 9172
rect 1952 9052 2004 9104
rect 3792 9052 3844 9104
rect 3884 9052 3936 9104
rect 4804 9095 4856 9104
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 10968 9052 11020 9104
rect 15936 9052 15988 9104
rect 17500 9095 17552 9104
rect 17500 9061 17509 9095
rect 17509 9061 17543 9095
rect 17543 9061 17552 9095
rect 17500 9052 17552 9061
rect 19432 9095 19484 9104
rect 19432 9061 19441 9095
rect 19441 9061 19475 9095
rect 19475 9061 19484 9095
rect 19432 9052 19484 9061
rect 21916 9095 21968 9104
rect 21916 9061 21925 9095
rect 21925 9061 21959 9095
rect 21959 9061 21968 9095
rect 21916 9052 21968 9061
rect 29276 9129 29285 9163
rect 29285 9129 29319 9163
rect 29319 9129 29328 9163
rect 29276 9120 29328 9129
rect 30380 9120 30432 9172
rect 34520 9163 34572 9172
rect 34520 9129 34529 9163
rect 34529 9129 34563 9163
rect 34563 9129 34572 9163
rect 34520 9120 34572 9129
rect 34980 9163 35032 9172
rect 34980 9129 34989 9163
rect 34989 9129 35023 9163
rect 35023 9129 35032 9163
rect 34980 9120 35032 9129
rect 35808 9120 35860 9172
rect 36176 9120 36228 9172
rect 36636 9163 36688 9172
rect 36636 9129 36645 9163
rect 36645 9129 36679 9163
rect 36679 9129 36688 9163
rect 36636 9120 36688 9129
rect 2320 8984 2372 9036
rect 3516 8984 3568 9036
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 6184 8984 6236 9036
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7472 8984 7524 9036
rect 11796 9027 11848 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 7288 8916 7340 8968
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 14188 9027 14240 9036
rect 14188 8993 14197 9027
rect 14197 8993 14231 9027
rect 14231 8993 14240 9027
rect 14188 8984 14240 8993
rect 23480 8984 23532 9036
rect 27528 9052 27580 9104
rect 27988 9052 28040 9104
rect 30656 9052 30708 9104
rect 34612 9052 34664 9104
rect 35900 9052 35952 9104
rect 26332 8984 26384 9036
rect 26700 8984 26752 9036
rect 32496 8984 32548 9036
rect 34428 8984 34480 9036
rect 36636 8984 36688 9036
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 15292 8959 15344 8968
rect 3976 8780 4028 8832
rect 12624 8848 12676 8900
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 17592 8916 17644 8968
rect 13268 8891 13320 8900
rect 13268 8857 13277 8891
rect 13277 8857 13311 8891
rect 13311 8857 13320 8891
rect 18512 8916 18564 8968
rect 20076 8916 20128 8968
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 13268 8848 13320 8857
rect 18144 8848 18196 8900
rect 24032 8916 24084 8968
rect 5172 8823 5224 8832
rect 5172 8789 5181 8823
rect 5181 8789 5215 8823
rect 5215 8789 5224 8823
rect 5172 8780 5224 8789
rect 5356 8780 5408 8832
rect 15200 8780 15252 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 21272 8780 21324 8832
rect 21364 8780 21416 8832
rect 27252 8916 27304 8968
rect 28172 8916 28224 8968
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 33048 8916 33100 8968
rect 33876 8916 33928 8968
rect 36268 8916 36320 8968
rect 22560 8780 22612 8832
rect 24124 8823 24176 8832
rect 24124 8789 24133 8823
rect 24133 8789 24167 8823
rect 24167 8789 24176 8823
rect 24124 8780 24176 8789
rect 26976 8780 27028 8832
rect 31484 8823 31536 8832
rect 31484 8789 31493 8823
rect 31493 8789 31527 8823
rect 31527 8789 31536 8823
rect 31484 8780 31536 8789
rect 32496 8823 32548 8832
rect 32496 8789 32505 8823
rect 32505 8789 32539 8823
rect 32539 8789 32548 8823
rect 32496 8780 32548 8789
rect 33140 8780 33192 8832
rect 33416 8780 33468 8832
rect 33600 8780 33652 8832
rect 35348 8780 35400 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3516 8576 3568 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9128 8576 9180 8628
rect 3884 8508 3936 8560
rect 5540 8508 5592 8560
rect 10876 8576 10928 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 13452 8576 13504 8628
rect 17500 8619 17552 8628
rect 10968 8551 11020 8560
rect 3148 8440 3200 8492
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 7656 8440 7708 8492
rect 8484 8440 8536 8492
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 12072 8508 12124 8560
rect 14188 8551 14240 8560
rect 14188 8517 14197 8551
rect 14197 8517 14231 8551
rect 14231 8517 14240 8551
rect 14188 8508 14240 8517
rect 4436 8415 4488 8424
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 2412 8236 2464 8288
rect 3608 8279 3660 8288
rect 3608 8245 3617 8279
rect 3617 8245 3651 8279
rect 3651 8245 3660 8279
rect 3608 8236 3660 8245
rect 4712 8304 4764 8356
rect 5724 8304 5776 8356
rect 7196 8304 7248 8356
rect 8024 8304 8076 8356
rect 9128 8304 9180 8356
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 6184 8279 6236 8288
rect 4344 8236 4396 8245
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 6644 8236 6696 8288
rect 7288 8236 7340 8288
rect 8576 8236 8628 8288
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 10048 8347 10100 8356
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 11152 8304 11204 8356
rect 12716 8304 12768 8356
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 17592 8576 17644 8628
rect 21364 8576 21416 8628
rect 21824 8576 21876 8628
rect 22928 8576 22980 8628
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16488 8440 16540 8492
rect 21916 8508 21968 8560
rect 22560 8551 22612 8560
rect 22560 8517 22569 8551
rect 22569 8517 22603 8551
rect 22603 8517 22612 8551
rect 22560 8508 22612 8517
rect 23480 8551 23532 8560
rect 23480 8517 23489 8551
rect 23489 8517 23523 8551
rect 23523 8517 23532 8551
rect 23480 8508 23532 8517
rect 19432 8440 19484 8492
rect 26332 8576 26384 8628
rect 27528 8576 27580 8628
rect 29000 8619 29052 8628
rect 29000 8585 29009 8619
rect 29009 8585 29043 8619
rect 29043 8585 29052 8619
rect 29000 8576 29052 8585
rect 32312 8619 32364 8628
rect 32312 8585 32321 8619
rect 32321 8585 32355 8619
rect 32355 8585 32364 8619
rect 32312 8576 32364 8585
rect 32496 8576 32548 8628
rect 33600 8576 33652 8628
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 17132 8372 17184 8424
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 15292 8304 15344 8356
rect 15936 8304 15988 8356
rect 20444 8347 20496 8356
rect 20444 8313 20453 8347
rect 20453 8313 20487 8347
rect 20487 8313 20496 8347
rect 20444 8304 20496 8313
rect 20536 8347 20588 8356
rect 20536 8313 20545 8347
rect 20545 8313 20579 8347
rect 20579 8313 20588 8347
rect 20536 8304 20588 8313
rect 18604 8236 18656 8288
rect 20260 8279 20312 8288
rect 20260 8245 20269 8279
rect 20269 8245 20303 8279
rect 20303 8245 20312 8279
rect 20260 8236 20312 8245
rect 21364 8304 21416 8356
rect 21732 8304 21784 8356
rect 21916 8236 21968 8288
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 25412 8440 25464 8492
rect 27068 8483 27120 8492
rect 27068 8449 27077 8483
rect 27077 8449 27111 8483
rect 27111 8449 27120 8483
rect 27068 8440 27120 8449
rect 24584 8372 24636 8424
rect 26424 8372 26476 8424
rect 29092 8372 29144 8424
rect 30012 8372 30064 8424
rect 31484 8440 31536 8492
rect 32956 8440 33008 8492
rect 35256 8576 35308 8628
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 34612 8508 34664 8560
rect 34888 8508 34940 8560
rect 37188 8508 37240 8560
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 35716 8440 35768 8492
rect 30840 8372 30892 8424
rect 31300 8372 31352 8424
rect 23756 8304 23808 8356
rect 25044 8304 25096 8356
rect 26516 8304 26568 8356
rect 24400 8236 24452 8288
rect 26240 8279 26292 8288
rect 26240 8245 26249 8279
rect 26249 8245 26283 8279
rect 26283 8245 26292 8279
rect 26240 8236 26292 8245
rect 27068 8236 27120 8288
rect 27988 8279 28040 8288
rect 27988 8245 27997 8279
rect 27997 8245 28031 8279
rect 28031 8245 28040 8279
rect 27988 8236 28040 8245
rect 31576 8304 31628 8356
rect 33324 8304 33376 8356
rect 33416 8347 33468 8356
rect 33416 8313 33425 8347
rect 33425 8313 33459 8347
rect 33459 8313 33468 8347
rect 33968 8347 34020 8356
rect 33416 8304 33468 8313
rect 33968 8313 33977 8347
rect 33977 8313 34011 8347
rect 34011 8313 34020 8347
rect 33968 8304 34020 8313
rect 33048 8279 33100 8288
rect 33048 8245 33057 8279
rect 33057 8245 33091 8279
rect 33091 8245 33100 8279
rect 33048 8236 33100 8245
rect 36176 8304 36228 8356
rect 36544 8347 36596 8356
rect 36544 8313 36553 8347
rect 36553 8313 36587 8347
rect 36587 8313 36596 8347
rect 36544 8304 36596 8313
rect 36636 8347 36688 8356
rect 36636 8313 36645 8347
rect 36645 8313 36679 8347
rect 36679 8313 36688 8347
rect 36636 8304 36688 8313
rect 35900 8279 35952 8288
rect 35900 8245 35909 8279
rect 35909 8245 35943 8279
rect 35943 8245 35952 8279
rect 35900 8236 35952 8245
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4436 8032 4488 8084
rect 6828 8032 6880 8084
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 12624 8075 12676 8084
rect 7196 8032 7248 8041
rect 1860 7964 1912 8016
rect 2504 7964 2556 8016
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 3056 7964 3108 8016
rect 3608 7964 3660 8016
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 4804 8007 4856 8016
rect 4804 7973 4813 8007
rect 4813 7973 4847 8007
rect 4847 7973 4856 8007
rect 4804 7964 4856 7973
rect 10048 7964 10100 8016
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3516 7896 3568 7948
rect 6092 7896 6144 7948
rect 7472 7896 7524 7948
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 15292 8032 15344 8084
rect 22468 8032 22520 8084
rect 12072 7964 12124 8016
rect 13544 7964 13596 8016
rect 15108 7964 15160 8016
rect 11612 7896 11664 7948
rect 11796 7896 11848 7948
rect 15752 7896 15804 7948
rect 16488 7964 16540 8016
rect 18604 7964 18656 8016
rect 20076 7964 20128 8016
rect 20260 7964 20312 8016
rect 20536 7964 20588 8016
rect 21916 8007 21968 8016
rect 21916 7973 21925 8007
rect 21925 7973 21959 8007
rect 21959 7973 21968 8007
rect 21916 7964 21968 7973
rect 23204 8032 23256 8084
rect 25412 8075 25464 8084
rect 23756 8007 23808 8016
rect 23756 7973 23765 8007
rect 23765 7973 23799 8007
rect 23799 7973 23808 8007
rect 23756 7964 23808 7973
rect 25412 8041 25421 8075
rect 25421 8041 25455 8075
rect 25455 8041 25464 8075
rect 25412 8032 25464 8041
rect 27988 8032 28040 8084
rect 29000 8032 29052 8084
rect 30012 8075 30064 8084
rect 30012 8041 30021 8075
rect 30021 8041 30055 8075
rect 30055 8041 30064 8075
rect 30012 8032 30064 8041
rect 32956 8075 33008 8084
rect 32956 8041 32965 8075
rect 32965 8041 32999 8075
rect 32999 8041 33008 8075
rect 32956 8032 33008 8041
rect 33324 8032 33376 8084
rect 37740 8032 37792 8084
rect 24400 7964 24452 8016
rect 26240 7964 26292 8016
rect 26792 7964 26844 8016
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 17316 7896 17368 7948
rect 21732 7896 21784 7948
rect 28908 7939 28960 7948
rect 28908 7905 28917 7939
rect 28917 7905 28951 7939
rect 28951 7905 28960 7939
rect 28908 7896 28960 7905
rect 29920 7964 29972 8016
rect 33048 7964 33100 8016
rect 35072 8007 35124 8016
rect 35072 7973 35081 8007
rect 35081 7973 35115 8007
rect 35115 7973 35124 8007
rect 35072 7964 35124 7973
rect 30472 7939 30524 7948
rect 30472 7905 30481 7939
rect 30481 7905 30515 7939
rect 30515 7905 30524 7939
rect 30472 7896 30524 7905
rect 30840 7896 30892 7948
rect 36268 7896 36320 7948
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 5540 7828 5592 7880
rect 6920 7828 6972 7880
rect 8116 7828 8168 7880
rect 8852 7828 8904 7880
rect 10140 7828 10192 7880
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 20352 7828 20404 7880
rect 21824 7828 21876 7880
rect 22008 7828 22060 7880
rect 22652 7828 22704 7880
rect 2320 7760 2372 7812
rect 7196 7760 7248 7812
rect 18880 7760 18932 7812
rect 20444 7803 20496 7812
rect 20444 7769 20453 7803
rect 20453 7769 20487 7803
rect 20487 7769 20496 7803
rect 20444 7760 20496 7769
rect 24032 7760 24084 7812
rect 26332 7828 26384 7880
rect 27252 7871 27304 7880
rect 27252 7837 27261 7871
rect 27261 7837 27295 7871
rect 27295 7837 27304 7871
rect 27252 7828 27304 7837
rect 33048 7871 33100 7880
rect 33048 7837 33057 7871
rect 33057 7837 33091 7871
rect 33091 7837 33100 7871
rect 33048 7828 33100 7837
rect 33968 7828 34020 7880
rect 35716 7828 35768 7880
rect 35532 7803 35584 7812
rect 35532 7769 35541 7803
rect 35541 7769 35575 7803
rect 35575 7769 35584 7803
rect 35532 7760 35584 7769
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 8024 7692 8076 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8760 7692 8812 7744
rect 9312 7692 9364 7744
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 11060 7692 11112 7744
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 18512 7692 18564 7744
rect 34152 7692 34204 7744
rect 35256 7692 35308 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 2964 7488 3016 7540
rect 3056 7488 3108 7540
rect 4252 7488 4304 7540
rect 8576 7488 8628 7540
rect 9036 7488 9088 7540
rect 11244 7488 11296 7540
rect 15476 7488 15528 7540
rect 15752 7488 15804 7540
rect 18052 7488 18104 7540
rect 19064 7488 19116 7540
rect 20260 7488 20312 7540
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 23204 7488 23256 7540
rect 26792 7531 26844 7540
rect 26792 7497 26801 7531
rect 26801 7497 26835 7531
rect 26835 7497 26844 7531
rect 26792 7488 26844 7497
rect 29092 7531 29144 7540
rect 29092 7497 29101 7531
rect 29101 7497 29135 7531
rect 29135 7497 29144 7531
rect 29092 7488 29144 7497
rect 30472 7531 30524 7540
rect 30472 7497 30481 7531
rect 30481 7497 30515 7531
rect 30515 7497 30524 7531
rect 30472 7488 30524 7497
rect 34152 7488 34204 7540
rect 6092 7420 6144 7472
rect 6460 7420 6512 7472
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 9312 7420 9364 7472
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2964 7284 3016 7336
rect 4344 7259 4396 7268
rect 4344 7225 4347 7259
rect 4347 7225 4381 7259
rect 4381 7225 4396 7259
rect 4344 7216 4396 7225
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 8116 7352 8168 7404
rect 9220 7352 9272 7404
rect 9588 7395 9640 7404
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 9588 7352 9640 7361
rect 13728 7420 13780 7472
rect 17776 7463 17828 7472
rect 11520 7395 11572 7404
rect 8208 7284 8260 7336
rect 8668 7284 8720 7336
rect 7656 7259 7708 7268
rect 7656 7225 7665 7259
rect 7665 7225 7699 7259
rect 7699 7225 7708 7259
rect 7656 7216 7708 7225
rect 8852 7216 8904 7268
rect 10876 7284 10928 7336
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11152 7284 11204 7336
rect 12164 7284 12216 7336
rect 17776 7429 17785 7463
rect 17785 7429 17819 7463
rect 17819 7429 17828 7463
rect 17776 7420 17828 7429
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 15108 7327 15160 7336
rect 15108 7293 15117 7327
rect 15117 7293 15151 7327
rect 15151 7293 15160 7327
rect 15108 7284 15160 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 18788 7284 18840 7336
rect 7196 7148 7248 7157
rect 11704 7148 11756 7200
rect 12072 7148 12124 7200
rect 12900 7216 12952 7268
rect 21272 7352 21324 7404
rect 26332 7420 26384 7472
rect 26976 7352 27028 7404
rect 27528 7352 27580 7404
rect 33416 7420 33468 7472
rect 36636 7420 36688 7472
rect 30656 7352 30708 7404
rect 33784 7352 33836 7404
rect 35256 7352 35308 7404
rect 35624 7352 35676 7404
rect 20812 7216 20864 7268
rect 21824 7259 21876 7268
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 17316 7148 17368 7200
rect 21824 7225 21833 7259
rect 21833 7225 21867 7259
rect 21867 7225 21876 7259
rect 21824 7216 21876 7225
rect 26608 7284 26660 7336
rect 29092 7284 29144 7336
rect 29736 7327 29788 7336
rect 29736 7293 29745 7327
rect 29745 7293 29779 7327
rect 29779 7293 29788 7327
rect 29736 7284 29788 7293
rect 31116 7327 31168 7336
rect 31116 7293 31125 7327
rect 31125 7293 31159 7327
rect 31159 7293 31168 7327
rect 31116 7284 31168 7293
rect 32864 7284 32916 7336
rect 21732 7148 21784 7200
rect 22008 7148 22060 7200
rect 23940 7191 23992 7200
rect 23940 7157 23949 7191
rect 23949 7157 23983 7191
rect 23983 7157 23992 7191
rect 23940 7148 23992 7157
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 25596 7148 25648 7200
rect 26700 7148 26752 7200
rect 27160 7191 27212 7200
rect 27160 7157 27169 7191
rect 27169 7157 27203 7191
rect 27203 7157 27212 7191
rect 27160 7148 27212 7157
rect 27436 7148 27488 7200
rect 28908 7148 28960 7200
rect 29552 7191 29604 7200
rect 29552 7157 29561 7191
rect 29561 7157 29595 7191
rect 29595 7157 29604 7191
rect 29552 7148 29604 7157
rect 33324 7148 33376 7200
rect 34060 7148 34112 7200
rect 34612 7148 34664 7200
rect 35716 7216 35768 7268
rect 36360 7216 36412 7268
rect 36636 7259 36688 7268
rect 36636 7225 36645 7259
rect 36645 7225 36679 7259
rect 36679 7225 36688 7259
rect 36636 7216 36688 7225
rect 36268 7191 36320 7200
rect 36268 7157 36277 7191
rect 36277 7157 36311 7191
rect 36311 7157 36320 7191
rect 36268 7148 36320 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1860 6987 1912 6996
rect 1860 6953 1869 6987
rect 1869 6953 1903 6987
rect 1903 6953 1912 6987
rect 1860 6944 1912 6953
rect 3792 6944 3844 6996
rect 4160 6944 4212 6996
rect 4436 6944 4488 6996
rect 6184 6944 6236 6996
rect 7656 6944 7708 6996
rect 9496 6944 9548 6996
rect 10140 6944 10192 6996
rect 16856 6944 16908 6996
rect 20352 6987 20404 6996
rect 20352 6953 20361 6987
rect 20361 6953 20395 6987
rect 20395 6953 20404 6987
rect 20352 6944 20404 6953
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 21732 6944 21784 6996
rect 22744 6987 22796 6996
rect 22744 6953 22753 6987
rect 22753 6953 22787 6987
rect 22787 6953 22796 6987
rect 22744 6944 22796 6953
rect 24400 6987 24452 6996
rect 24400 6953 24409 6987
rect 24409 6953 24443 6987
rect 24443 6953 24452 6987
rect 24400 6944 24452 6953
rect 2504 6876 2556 6928
rect 4252 6919 4304 6928
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 4896 6876 4948 6928
rect 6920 6876 6972 6928
rect 8760 6919 8812 6928
rect 8760 6885 8769 6919
rect 8769 6885 8803 6919
rect 8803 6885 8812 6919
rect 8760 6876 8812 6885
rect 10876 6919 10928 6928
rect 10876 6885 10885 6919
rect 10885 6885 10919 6919
rect 10919 6885 10928 6919
rect 10876 6876 10928 6885
rect 11612 6876 11664 6928
rect 12072 6876 12124 6928
rect 16028 6876 16080 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 6092 6808 6144 6860
rect 3608 6740 3660 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4436 6783 4488 6792
rect 4160 6740 4212 6749
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6368 6740 6420 6792
rect 8024 6808 8076 6860
rect 9956 6851 10008 6860
rect 8116 6783 8168 6792
rect 3976 6672 4028 6724
rect 4804 6672 4856 6724
rect 1768 6604 1820 6656
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2688 6604 2740 6656
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 7012 6604 7064 6656
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 9404 6740 9456 6792
rect 9956 6817 9965 6851
rect 9965 6817 9999 6851
rect 9999 6817 10008 6851
rect 9956 6808 10008 6817
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 14280 6808 14332 6860
rect 17684 6808 17736 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 18696 6876 18748 6928
rect 21364 6876 21416 6928
rect 26332 6944 26384 6996
rect 27528 6987 27580 6996
rect 27528 6953 27537 6987
rect 27537 6953 27571 6987
rect 27571 6953 27580 6987
rect 27528 6944 27580 6953
rect 31116 6944 31168 6996
rect 33416 6944 33468 6996
rect 34060 6987 34112 6996
rect 34060 6953 34069 6987
rect 34069 6953 34103 6987
rect 34103 6953 34112 6987
rect 34060 6944 34112 6953
rect 35072 6944 35124 6996
rect 25044 6919 25096 6928
rect 25044 6885 25053 6919
rect 25053 6885 25087 6919
rect 25087 6885 25096 6919
rect 25044 6876 25096 6885
rect 26700 6919 26752 6928
rect 26700 6885 26709 6919
rect 26709 6885 26743 6919
rect 26743 6885 26752 6919
rect 26700 6876 26752 6885
rect 27252 6919 27304 6928
rect 27252 6885 27261 6919
rect 27261 6885 27295 6919
rect 27295 6885 27304 6919
rect 27252 6876 27304 6885
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 22836 6851 22888 6860
rect 11796 6740 11848 6792
rect 12992 6740 13044 6792
rect 16304 6740 16356 6792
rect 22836 6817 22845 6851
rect 22845 6817 22879 6851
rect 22879 6817 22888 6851
rect 22836 6808 22888 6817
rect 20628 6740 20680 6792
rect 22376 6740 22428 6792
rect 28632 6808 28684 6860
rect 30104 6876 30156 6928
rect 33876 6876 33928 6928
rect 35900 6876 35952 6928
rect 29000 6851 29052 6860
rect 29000 6817 29009 6851
rect 29009 6817 29043 6851
rect 29043 6817 29052 6851
rect 29000 6808 29052 6817
rect 29736 6808 29788 6860
rect 30380 6851 30432 6860
rect 30380 6817 30389 6851
rect 30389 6817 30423 6851
rect 30423 6817 30432 6851
rect 30380 6808 30432 6817
rect 24124 6740 24176 6792
rect 24952 6783 25004 6792
rect 24952 6749 24961 6783
rect 24961 6749 24995 6783
rect 24995 6749 25004 6783
rect 24952 6740 25004 6749
rect 7472 6604 7524 6656
rect 8668 6672 8720 6724
rect 21824 6672 21876 6724
rect 28172 6740 28224 6792
rect 29276 6783 29328 6792
rect 29276 6749 29285 6783
rect 29285 6749 29319 6783
rect 29319 6749 29328 6783
rect 29276 6740 29328 6749
rect 30840 6740 30892 6792
rect 28908 6672 28960 6724
rect 32404 6808 32456 6860
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 34704 6808 34756 6860
rect 36360 6808 36412 6860
rect 33600 6740 33652 6792
rect 35440 6783 35492 6792
rect 35440 6749 35449 6783
rect 35449 6749 35483 6783
rect 35483 6749 35492 6783
rect 35440 6740 35492 6749
rect 35072 6672 35124 6724
rect 8576 6604 8628 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 11152 6604 11204 6656
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 15108 6604 15160 6656
rect 15476 6604 15528 6656
rect 16580 6604 16632 6656
rect 18236 6604 18288 6656
rect 18788 6604 18840 6656
rect 20536 6604 20588 6656
rect 20812 6604 20864 6656
rect 23848 6604 23900 6656
rect 25320 6604 25372 6656
rect 30012 6647 30064 6656
rect 30012 6613 30021 6647
rect 30021 6613 30055 6647
rect 30055 6613 30064 6647
rect 30012 6604 30064 6613
rect 31392 6604 31444 6656
rect 33048 6604 33100 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 3148 6400 3200 6452
rect 4344 6400 4396 6452
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 4252 6332 4304 6384
rect 4804 6375 4856 6384
rect 4804 6341 4813 6375
rect 4813 6341 4847 6375
rect 4847 6341 4856 6375
rect 4804 6332 4856 6341
rect 7012 6332 7064 6384
rect 8024 6400 8076 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 12072 6400 12124 6452
rect 13360 6400 13412 6452
rect 14372 6400 14424 6452
rect 15936 6443 15988 6452
rect 10324 6332 10376 6384
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 16856 6400 16908 6452
rect 20812 6400 20864 6452
rect 21732 6400 21784 6452
rect 25044 6400 25096 6452
rect 27160 6400 27212 6452
rect 28172 6443 28224 6452
rect 28172 6409 28181 6443
rect 28181 6409 28215 6443
rect 28215 6409 28224 6443
rect 28172 6400 28224 6409
rect 28632 6443 28684 6452
rect 28632 6409 28641 6443
rect 28641 6409 28675 6443
rect 28675 6409 28684 6443
rect 28632 6400 28684 6409
rect 30840 6400 30892 6452
rect 32588 6400 32640 6452
rect 34060 6400 34112 6452
rect 35900 6443 35952 6452
rect 35900 6409 35909 6443
rect 35909 6409 35943 6443
rect 35943 6409 35952 6443
rect 35900 6400 35952 6409
rect 36636 6443 36688 6452
rect 36636 6409 36645 6443
rect 36645 6409 36679 6443
rect 36679 6409 36688 6443
rect 36636 6400 36688 6409
rect 37096 6443 37148 6452
rect 37096 6409 37105 6443
rect 37105 6409 37139 6443
rect 37139 6409 37148 6443
rect 37096 6400 37148 6409
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 3792 6264 3844 6316
rect 2044 6196 2096 6248
rect 7196 6264 7248 6316
rect 3148 6128 3200 6180
rect 4252 6171 4304 6180
rect 4252 6137 4261 6171
rect 4261 6137 4295 6171
rect 4295 6137 4304 6171
rect 4252 6128 4304 6137
rect 4344 6171 4396 6180
rect 4344 6137 4353 6171
rect 4353 6137 4387 6171
rect 4387 6137 4396 6171
rect 4344 6128 4396 6137
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 7104 6239 7156 6248
rect 6920 6196 6972 6205
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 11152 6264 11204 6316
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 13360 6196 13412 6248
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 6092 6060 6144 6112
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9956 6060 10008 6112
rect 10784 6128 10836 6180
rect 12072 6128 12124 6180
rect 19248 6332 19300 6384
rect 14280 6264 14332 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 15752 6264 15804 6316
rect 17868 6264 17920 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 16672 6196 16724 6248
rect 21272 6264 21324 6316
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 23020 6239 23072 6248
rect 23020 6205 23029 6239
rect 23029 6205 23063 6239
rect 23063 6205 23072 6239
rect 23020 6196 23072 6205
rect 23572 6332 23624 6384
rect 32404 6332 32456 6384
rect 35532 6375 35584 6384
rect 35532 6341 35541 6375
rect 35541 6341 35575 6375
rect 35575 6341 35584 6375
rect 35532 6332 35584 6341
rect 23848 6239 23900 6248
rect 23848 6205 23857 6239
rect 23857 6205 23891 6239
rect 23891 6205 23900 6239
rect 23848 6196 23900 6205
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 25504 6196 25556 6248
rect 27436 6196 27488 6248
rect 29000 6264 29052 6316
rect 33232 6307 33284 6316
rect 31484 6239 31536 6248
rect 31484 6205 31493 6239
rect 31493 6205 31527 6239
rect 31527 6205 31536 6239
rect 31484 6196 31536 6205
rect 33232 6273 33241 6307
rect 33241 6273 33275 6307
rect 33275 6273 33284 6307
rect 33232 6264 33284 6273
rect 33692 6307 33744 6316
rect 33692 6273 33701 6307
rect 33701 6273 33735 6307
rect 33735 6273 33744 6307
rect 33692 6264 33744 6273
rect 34704 6264 34756 6316
rect 35440 6264 35492 6316
rect 36360 6196 36412 6248
rect 37096 6196 37148 6248
rect 38016 6239 38068 6248
rect 38016 6205 38025 6239
rect 38025 6205 38059 6239
rect 38059 6205 38068 6239
rect 38016 6196 38068 6205
rect 14372 6171 14424 6180
rect 14372 6137 14381 6171
rect 14381 6137 14415 6171
rect 14415 6137 14424 6171
rect 14372 6128 14424 6137
rect 15936 6128 15988 6180
rect 18144 6171 18196 6180
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 18236 6171 18288 6180
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 18236 6128 18288 6137
rect 20536 6128 20588 6180
rect 13176 6060 13228 6112
rect 14188 6060 14240 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 19800 6060 19852 6112
rect 22836 6128 22888 6180
rect 23940 6128 23992 6180
rect 24860 6128 24912 6180
rect 25596 6128 25648 6180
rect 27068 6128 27120 6180
rect 29736 6128 29788 6180
rect 30012 6171 30064 6180
rect 30012 6137 30021 6171
rect 30021 6137 30055 6171
rect 30055 6137 30064 6171
rect 30564 6171 30616 6180
rect 30012 6128 30064 6137
rect 30564 6137 30573 6171
rect 30573 6137 30607 6171
rect 30607 6137 30616 6171
rect 30564 6128 30616 6137
rect 32128 6171 32180 6180
rect 32128 6137 32137 6171
rect 32137 6137 32171 6171
rect 32171 6137 32180 6171
rect 32128 6128 32180 6137
rect 33416 6128 33468 6180
rect 34796 6128 34848 6180
rect 35072 6171 35124 6180
rect 35072 6137 35081 6171
rect 35081 6137 35115 6171
rect 35115 6137 35124 6171
rect 35072 6128 35124 6137
rect 35256 6128 35308 6180
rect 21732 6060 21784 6112
rect 22376 6103 22428 6112
rect 22376 6069 22385 6103
rect 22385 6069 22419 6103
rect 22419 6069 22428 6103
rect 22376 6060 22428 6069
rect 22928 6060 22980 6112
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 27252 6103 27304 6112
rect 27252 6069 27261 6103
rect 27261 6069 27295 6103
rect 27295 6069 27304 6103
rect 27252 6060 27304 6069
rect 30380 6060 30432 6112
rect 31208 6060 31260 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 1400 5856 1452 5908
rect 1768 5856 1820 5908
rect 2412 5856 2464 5908
rect 3148 5856 3200 5908
rect 3608 5899 3660 5908
rect 3608 5865 3617 5899
rect 3617 5865 3651 5899
rect 3651 5865 3660 5899
rect 3608 5856 3660 5865
rect 4160 5856 4212 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6920 5856 6972 5908
rect 5172 5788 5224 5840
rect 7104 5788 7156 5840
rect 1860 5720 1912 5772
rect 4988 5720 5040 5772
rect 5448 5720 5500 5772
rect 8392 5856 8444 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 12072 5856 12124 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 18144 5856 18196 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 22928 5856 22980 5908
rect 24952 5856 25004 5908
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 33232 5856 33284 5908
rect 7380 5788 7432 5840
rect 8668 5788 8720 5840
rect 10140 5788 10192 5840
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 10784 5788 10836 5797
rect 13176 5831 13228 5840
rect 13176 5797 13185 5831
rect 13185 5797 13219 5831
rect 13219 5797 13228 5831
rect 13176 5788 13228 5797
rect 15108 5788 15160 5840
rect 16948 5788 17000 5840
rect 17408 5788 17460 5840
rect 18052 5788 18104 5840
rect 20628 5831 20680 5840
rect 20628 5797 20637 5831
rect 20637 5797 20671 5831
rect 20671 5797 20680 5831
rect 20628 5788 20680 5797
rect 21180 5831 21232 5840
rect 21180 5797 21189 5831
rect 21189 5797 21223 5831
rect 21223 5797 21232 5831
rect 21180 5788 21232 5797
rect 21916 5788 21968 5840
rect 23296 5788 23348 5840
rect 25596 5788 25648 5840
rect 27160 5788 27212 5840
rect 29000 5788 29052 5840
rect 32496 5788 32548 5840
rect 34612 5831 34664 5840
rect 34612 5797 34621 5831
rect 34621 5797 34655 5831
rect 34655 5797 34664 5831
rect 34612 5788 34664 5797
rect 8024 5720 8076 5772
rect 8484 5720 8536 5772
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 6644 5652 6696 5704
rect 7196 5652 7248 5704
rect 2136 5627 2188 5636
rect 2136 5593 2145 5627
rect 2145 5593 2179 5627
rect 2179 5593 2188 5627
rect 2136 5584 2188 5593
rect 4252 5516 4304 5568
rect 6552 5516 6604 5568
rect 7472 5652 7524 5704
rect 8116 5652 8168 5704
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 10232 5652 10284 5704
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 14832 5652 14884 5704
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 13636 5627 13688 5636
rect 13636 5593 13645 5627
rect 13645 5593 13679 5627
rect 13679 5593 13688 5627
rect 18328 5652 18380 5704
rect 19708 5652 19760 5704
rect 20812 5720 20864 5772
rect 22744 5720 22796 5772
rect 23756 5720 23808 5772
rect 25136 5720 25188 5772
rect 27252 5720 27304 5772
rect 29276 5720 29328 5772
rect 32128 5720 32180 5772
rect 35532 5720 35584 5772
rect 36728 5720 36780 5772
rect 24676 5652 24728 5704
rect 33140 5652 33192 5704
rect 34152 5652 34204 5704
rect 34704 5652 34756 5704
rect 13636 5584 13688 5593
rect 18420 5584 18472 5636
rect 29736 5584 29788 5636
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 12992 5516 13044 5568
rect 13452 5516 13504 5568
rect 14188 5516 14240 5568
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 22192 5516 22244 5568
rect 24124 5559 24176 5568
rect 24124 5525 24133 5559
rect 24133 5525 24167 5559
rect 24167 5525 24176 5559
rect 24124 5516 24176 5525
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 25320 5516 25372 5568
rect 25504 5559 25556 5568
rect 25504 5525 25513 5559
rect 25513 5525 25547 5559
rect 25547 5525 25556 5559
rect 25504 5516 25556 5525
rect 27988 5559 28040 5568
rect 27988 5525 27997 5559
rect 27997 5525 28031 5559
rect 28031 5525 28040 5559
rect 27988 5516 28040 5525
rect 29920 5516 29972 5568
rect 31484 5559 31536 5568
rect 31484 5525 31493 5559
rect 31493 5525 31527 5559
rect 31527 5525 31536 5559
rect 31484 5516 31536 5525
rect 32220 5516 32272 5568
rect 33324 5516 33376 5568
rect 33600 5516 33652 5568
rect 35900 5516 35952 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 2872 5312 2924 5364
rect 5448 5355 5500 5364
rect 5448 5321 5457 5355
rect 5457 5321 5491 5355
rect 5491 5321 5500 5355
rect 5448 5312 5500 5321
rect 4988 5287 5040 5296
rect 4988 5253 4997 5287
rect 4997 5253 5031 5287
rect 5031 5253 5040 5287
rect 4988 5244 5040 5253
rect 5816 5244 5868 5296
rect 5172 5176 5224 5228
rect 2412 5151 2464 5160
rect 2412 5117 2421 5151
rect 2421 5117 2455 5151
rect 2455 5117 2464 5151
rect 2412 5108 2464 5117
rect 2872 5108 2924 5160
rect 7288 5312 7340 5364
rect 9128 5312 9180 5364
rect 10140 5312 10192 5364
rect 11612 5312 11664 5364
rect 13176 5312 13228 5364
rect 13728 5312 13780 5364
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 15108 5355 15160 5364
rect 15108 5321 15117 5355
rect 15117 5321 15151 5355
rect 15151 5321 15160 5355
rect 15108 5312 15160 5321
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 17960 5312 18012 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 20536 5312 20588 5364
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 21916 5355 21968 5364
rect 21916 5321 21925 5355
rect 21925 5321 21959 5355
rect 21959 5321 21968 5355
rect 23296 5355 23348 5364
rect 21916 5312 21968 5321
rect 23296 5321 23305 5355
rect 23305 5321 23339 5355
rect 23339 5321 23348 5355
rect 23296 5312 23348 5321
rect 25136 5312 25188 5364
rect 27252 5312 27304 5364
rect 29276 5312 29328 5364
rect 30012 5312 30064 5364
rect 34612 5312 34664 5364
rect 36544 5312 36596 5364
rect 36728 5355 36780 5364
rect 36728 5321 36737 5355
rect 36737 5321 36771 5355
rect 36771 5321 36780 5355
rect 36728 5312 36780 5321
rect 7196 5176 7248 5228
rect 8300 5244 8352 5296
rect 9956 5244 10008 5296
rect 15384 5244 15436 5296
rect 18236 5244 18288 5296
rect 20628 5244 20680 5296
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 13728 5176 13780 5228
rect 13912 5176 13964 5228
rect 14648 5176 14700 5228
rect 14924 5176 14976 5228
rect 15660 5176 15712 5228
rect 17592 5176 17644 5228
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 8116 5151 8168 5160
rect 1676 5040 1728 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 7196 5040 7248 5092
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 8300 5151 8352 5160
rect 8300 5117 8309 5151
rect 8309 5117 8343 5151
rect 8343 5117 8352 5151
rect 8300 5108 8352 5117
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 8024 5040 8076 5092
rect 9128 5040 9180 5092
rect 10232 5040 10284 5092
rect 12072 5108 12124 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 17684 5108 17736 5160
rect 17960 5108 18012 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 19708 5108 19760 5160
rect 22100 5176 22152 5228
rect 23204 5176 23256 5228
rect 24400 5176 24452 5228
rect 25320 5219 25372 5228
rect 25320 5185 25329 5219
rect 25329 5185 25363 5219
rect 25363 5185 25372 5219
rect 25320 5176 25372 5185
rect 29736 5244 29788 5296
rect 30564 5244 30616 5296
rect 36452 5287 36504 5296
rect 28172 5176 28224 5228
rect 29000 5219 29052 5228
rect 29000 5185 29009 5219
rect 29009 5185 29043 5219
rect 29043 5185 29052 5219
rect 29000 5176 29052 5185
rect 29552 5176 29604 5228
rect 36452 5253 36461 5287
rect 36461 5253 36495 5287
rect 36495 5253 36504 5287
rect 36452 5244 36504 5253
rect 27160 5151 27212 5160
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 13820 5040 13872 5092
rect 16488 5083 16540 5092
rect 16488 5049 16497 5083
rect 16497 5049 16531 5083
rect 16531 5049 16540 5083
rect 16488 5040 16540 5049
rect 16580 5083 16632 5092
rect 16580 5049 16589 5083
rect 16589 5049 16623 5083
rect 16623 5049 16632 5083
rect 16580 5040 16632 5049
rect 17224 5040 17276 5092
rect 27160 5117 27169 5151
rect 27169 5117 27203 5151
rect 27203 5117 27212 5151
rect 27160 5108 27212 5117
rect 21364 5040 21416 5092
rect 22100 5083 22152 5092
rect 22100 5049 22109 5083
rect 22109 5049 22143 5083
rect 22143 5049 22152 5083
rect 22100 5040 22152 5049
rect 22192 5083 22244 5092
rect 22192 5049 22201 5083
rect 22201 5049 22235 5083
rect 22235 5049 22244 5083
rect 22192 5040 22244 5049
rect 23848 5083 23900 5092
rect 23848 5049 23857 5083
rect 23857 5049 23891 5083
rect 23891 5049 23900 5083
rect 24400 5083 24452 5092
rect 23848 5040 23900 5049
rect 24400 5049 24409 5083
rect 24409 5049 24443 5083
rect 24443 5049 24452 5083
rect 25412 5083 25464 5092
rect 24400 5040 24452 5049
rect 25412 5049 25421 5083
rect 25421 5049 25455 5083
rect 25455 5049 25464 5083
rect 25412 5040 25464 5049
rect 27528 5040 27580 5092
rect 27988 5040 28040 5092
rect 31208 5151 31260 5160
rect 31208 5117 31217 5151
rect 31217 5117 31251 5151
rect 31251 5117 31260 5151
rect 31208 5108 31260 5117
rect 34612 5176 34664 5228
rect 34796 5176 34848 5228
rect 32588 5108 32640 5160
rect 29460 5040 29512 5092
rect 32496 5040 32548 5092
rect 33232 5083 33284 5092
rect 33232 5049 33241 5083
rect 33241 5049 33275 5083
rect 33275 5049 33284 5083
rect 33232 5040 33284 5049
rect 33324 5083 33376 5092
rect 33324 5049 33333 5083
rect 33333 5049 33367 5083
rect 33367 5049 33376 5083
rect 33324 5040 33376 5049
rect 31300 5015 31352 5024
rect 31300 4981 31309 5015
rect 31309 4981 31343 5015
rect 31343 4981 31352 5015
rect 31300 4972 31352 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2596 4632 2648 4684
rect 2872 4768 2924 4820
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 7012 4768 7064 4820
rect 7288 4768 7340 4820
rect 8668 4811 8720 4820
rect 2964 4743 3016 4752
rect 2964 4709 2973 4743
rect 2973 4709 3007 4743
rect 3007 4709 3016 4743
rect 2964 4700 3016 4709
rect 5448 4700 5500 4752
rect 6000 4700 6052 4752
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 5356 4632 5408 4684
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6920 4632 6972 4684
rect 7380 4632 7432 4684
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 9404 4811 9456 4820
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 9404 4768 9456 4777
rect 10232 4768 10284 4820
rect 8024 4700 8076 4752
rect 11612 4768 11664 4820
rect 11796 4768 11848 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 13084 4811 13136 4820
rect 13084 4777 13093 4811
rect 13093 4777 13127 4811
rect 13127 4777 13136 4811
rect 13084 4768 13136 4777
rect 10876 4700 10928 4752
rect 14832 4768 14884 4820
rect 16488 4811 16540 4820
rect 16488 4777 16497 4811
rect 16497 4777 16531 4811
rect 16531 4777 16540 4811
rect 16488 4768 16540 4777
rect 18512 4768 18564 4820
rect 18604 4768 18656 4820
rect 22100 4768 22152 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 23848 4811 23900 4820
rect 23848 4777 23857 4811
rect 23857 4777 23891 4811
rect 23891 4777 23900 4811
rect 23848 4768 23900 4777
rect 25320 4768 25372 4820
rect 27528 4768 27580 4820
rect 29460 4811 29512 4820
rect 29460 4777 29469 4811
rect 29469 4777 29503 4811
rect 29503 4777 29512 4811
rect 29460 4768 29512 4777
rect 31208 4811 31260 4820
rect 31208 4777 31217 4811
rect 31217 4777 31251 4811
rect 31251 4777 31260 4811
rect 31208 4768 31260 4777
rect 32128 4768 32180 4820
rect 33324 4768 33376 4820
rect 34152 4768 34204 4820
rect 13268 4700 13320 4752
rect 13912 4743 13964 4752
rect 13912 4709 13921 4743
rect 13921 4709 13955 4743
rect 13955 4709 13964 4743
rect 13912 4700 13964 4709
rect 16672 4700 16724 4752
rect 17408 4700 17460 4752
rect 22008 4700 22060 4752
rect 23756 4700 23808 4752
rect 24124 4743 24176 4752
rect 24124 4709 24133 4743
rect 24133 4709 24167 4743
rect 24167 4709 24176 4743
rect 24124 4700 24176 4709
rect 25412 4700 25464 4752
rect 27988 4700 28040 4752
rect 29920 4743 29972 4752
rect 29920 4709 29929 4743
rect 29929 4709 29963 4743
rect 29963 4709 29972 4743
rect 29920 4700 29972 4709
rect 30564 4700 30616 4752
rect 32864 4743 32916 4752
rect 32864 4709 32873 4743
rect 32873 4709 32907 4743
rect 32907 4709 32916 4743
rect 32864 4700 32916 4709
rect 12440 4632 12492 4684
rect 15476 4675 15528 4684
rect 15476 4641 15485 4675
rect 15485 4641 15519 4675
rect 15519 4641 15528 4675
rect 15476 4632 15528 4641
rect 15936 4632 15988 4684
rect 18788 4632 18840 4684
rect 19800 4675 19852 4684
rect 7472 4564 7524 4616
rect 10784 4564 10836 4616
rect 6460 4496 6512 4548
rect 8024 4496 8076 4548
rect 11244 4539 11296 4548
rect 11244 4505 11253 4539
rect 11253 4505 11287 4539
rect 11287 4505 11296 4539
rect 11244 4496 11296 4505
rect 13176 4496 13228 4548
rect 15660 4564 15712 4616
rect 17500 4564 17552 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 13636 4496 13688 4548
rect 8484 4428 8536 4480
rect 15844 4496 15896 4548
rect 19800 4641 19844 4675
rect 19844 4641 19852 4675
rect 21272 4675 21324 4684
rect 19800 4632 19852 4641
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 22192 4632 22244 4684
rect 23112 4632 23164 4684
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 24400 4607 24452 4616
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 27620 4632 27672 4684
rect 32588 4675 32640 4684
rect 27988 4607 28040 4616
rect 23020 4496 23072 4548
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 27988 4564 28040 4573
rect 28172 4564 28224 4616
rect 29000 4564 29052 4616
rect 30104 4564 30156 4616
rect 32036 4564 32088 4616
rect 32588 4641 32597 4675
rect 32597 4641 32631 4675
rect 32631 4641 32640 4675
rect 32588 4632 32640 4641
rect 33232 4632 33284 4684
rect 34612 4632 34664 4684
rect 14924 4428 14976 4480
rect 18788 4428 18840 4480
rect 38568 4428 38620 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 2596 4224 2648 4276
rect 2688 4224 2740 4276
rect 3056 4267 3108 4276
rect 3056 4233 3065 4267
rect 3065 4233 3099 4267
rect 3099 4233 3108 4267
rect 3056 4224 3108 4233
rect 4252 4224 4304 4276
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 5632 4224 5684 4276
rect 6368 4224 6420 4276
rect 7012 4267 7064 4276
rect 7012 4233 7021 4267
rect 7021 4233 7055 4267
rect 7055 4233 7064 4267
rect 7012 4224 7064 4233
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 11704 4224 11756 4276
rect 12440 4224 12492 4276
rect 8668 4088 8720 4140
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 6092 4020 6144 4072
rect 7012 4020 7064 4072
rect 7748 4020 7800 4072
rect 10784 4156 10836 4208
rect 12900 4156 12952 4208
rect 13268 4224 13320 4276
rect 17224 4224 17276 4276
rect 17500 4267 17552 4276
rect 17500 4233 17509 4267
rect 17509 4233 17543 4267
rect 17543 4233 17552 4267
rect 17500 4224 17552 4233
rect 18328 4224 18380 4276
rect 19800 4267 19852 4276
rect 19800 4233 19809 4267
rect 19809 4233 19843 4267
rect 19843 4233 19852 4267
rect 19800 4224 19852 4233
rect 22376 4224 22428 4276
rect 24032 4224 24084 4276
rect 26424 4267 26476 4276
rect 26424 4233 26433 4267
rect 26433 4233 26467 4267
rect 26467 4233 26476 4267
rect 26424 4224 26476 4233
rect 27620 4267 27672 4276
rect 27620 4233 27629 4267
rect 27629 4233 27663 4267
rect 27663 4233 27672 4267
rect 27620 4224 27672 4233
rect 27896 4267 27948 4276
rect 27896 4233 27905 4267
rect 27905 4233 27939 4267
rect 27939 4233 27948 4267
rect 27896 4224 27948 4233
rect 27988 4224 28040 4276
rect 29000 4267 29052 4276
rect 29000 4233 29009 4267
rect 29009 4233 29043 4267
rect 29043 4233 29052 4267
rect 29000 4224 29052 4233
rect 34612 4224 34664 4276
rect 14096 4156 14148 4208
rect 15292 4156 15344 4208
rect 15476 4156 15528 4208
rect 24676 4156 24728 4208
rect 25412 4156 25464 4208
rect 28080 4156 28132 4208
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 13360 4088 13412 4140
rect 15016 4088 15068 4140
rect 16304 4131 16356 4140
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 14004 4063 14056 4072
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 7196 3995 7248 4004
rect 7196 3961 7205 3995
rect 7205 3961 7239 3995
rect 7239 3961 7248 3995
rect 7196 3952 7248 3961
rect 9128 3952 9180 4004
rect 10508 3952 10560 4004
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 2412 3884 2464 3936
rect 8300 3884 8352 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 15292 4020 15344 4072
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17408 4088 17460 4140
rect 18788 4088 18840 4140
rect 21272 4131 21324 4140
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 19156 4020 19208 4072
rect 20720 4020 20772 4072
rect 22468 4020 22520 4072
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25412 4063 25464 4072
rect 25412 4029 25421 4063
rect 25421 4029 25455 4063
rect 25455 4029 25464 4063
rect 25412 4020 25464 4029
rect 30472 4088 30524 4140
rect 31392 4131 31444 4140
rect 26332 4020 26384 4072
rect 27528 4020 27580 4072
rect 29276 4063 29328 4072
rect 10600 3884 10652 3893
rect 12348 3884 12400 3936
rect 18604 3927 18656 3936
rect 18604 3893 18613 3927
rect 18613 3893 18647 3927
rect 18647 3893 18656 3927
rect 18604 3884 18656 3893
rect 23112 3884 23164 3936
rect 24032 3884 24084 3936
rect 24216 3927 24268 3936
rect 24216 3893 24225 3927
rect 24225 3893 24259 3927
rect 24259 3893 24268 3927
rect 24216 3884 24268 3893
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 29276 4029 29285 4063
rect 29285 4029 29319 4063
rect 29319 4029 29328 4063
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 29276 4020 29328 4029
rect 33600 4088 33652 4140
rect 30932 3952 30984 4004
rect 32220 4020 32272 4072
rect 32496 4063 32548 4072
rect 32496 4029 32505 4063
rect 32505 4029 32539 4063
rect 32539 4029 32548 4063
rect 32496 4020 32548 4029
rect 32588 4020 32640 4072
rect 30472 3884 30524 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 2872 3680 2924 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 6552 3723 6604 3732
rect 6552 3689 6561 3723
rect 6561 3689 6595 3723
rect 6595 3689 6604 3723
rect 6552 3680 6604 3689
rect 6920 3723 6972 3732
rect 6920 3689 6929 3723
rect 6929 3689 6963 3723
rect 6963 3689 6972 3723
rect 6920 3680 6972 3689
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 10692 3680 10744 3732
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 12808 3680 12860 3732
rect 13176 3680 13228 3732
rect 13452 3723 13504 3732
rect 13452 3689 13461 3723
rect 13461 3689 13495 3723
rect 13495 3689 13504 3723
rect 13452 3680 13504 3689
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 15752 3680 15804 3732
rect 16028 3723 16080 3732
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 16488 3680 16540 3732
rect 18880 3680 18932 3732
rect 19156 3723 19208 3732
rect 19156 3689 19165 3723
rect 19165 3689 19199 3723
rect 19199 3689 19208 3723
rect 19156 3680 19208 3689
rect 23020 3680 23072 3732
rect 24124 3680 24176 3732
rect 24676 3680 24728 3732
rect 27988 3723 28040 3732
rect 27988 3689 27997 3723
rect 27997 3689 28031 3723
rect 28031 3689 28040 3723
rect 27988 3680 28040 3689
rect 29920 3680 29972 3732
rect 32036 3680 32088 3732
rect 32496 3680 32548 3732
rect 3608 3612 3660 3664
rect 7748 3655 7800 3664
rect 7748 3621 7757 3655
rect 7757 3621 7791 3655
rect 7791 3621 7800 3655
rect 7748 3612 7800 3621
rect 8484 3612 8536 3664
rect 24216 3612 24268 3664
rect 28816 3612 28868 3664
rect 35440 3612 35492 3664
rect 2412 3544 2464 3596
rect 5908 3544 5960 3596
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 10784 3587 10836 3596
rect 10784 3553 10793 3587
rect 10793 3553 10827 3587
rect 10827 3553 10836 3587
rect 10784 3544 10836 3553
rect 12256 3544 12308 3596
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 15476 3587 15528 3596
rect 12348 3544 12400 3553
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 15568 3544 15620 3596
rect 16764 3587 16816 3596
rect 16764 3553 16808 3587
rect 16808 3553 16816 3587
rect 16764 3544 16816 3553
rect 28080 3544 28132 3596
rect 30748 3544 30800 3596
rect 30932 3587 30984 3596
rect 30932 3553 30941 3587
rect 30941 3553 30975 3587
rect 30975 3553 30984 3587
rect 30932 3544 30984 3553
rect 7380 3408 7432 3460
rect 8024 3451 8076 3460
rect 8024 3417 8033 3451
rect 8033 3417 8067 3451
rect 8067 3417 8076 3451
rect 8024 3408 8076 3417
rect 7288 3340 7340 3392
rect 8116 3340 8168 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2412 3136 2464 3188
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 7472 3136 7524 3188
rect 8024 3136 8076 3188
rect 8484 3136 8536 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10784 3136 10836 3188
rect 12256 3136 12308 3188
rect 13084 3136 13136 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 17684 3136 17736 3188
rect 30748 3179 30800 3188
rect 30748 3145 30757 3179
rect 30757 3145 30791 3179
rect 30791 3145 30800 3179
rect 30748 3136 30800 3145
rect 11060 3068 11112 3120
rect 16764 3111 16816 3120
rect 16764 3077 16773 3111
rect 16773 3077 16807 3111
rect 16807 3077 16816 3111
rect 16764 3068 16816 3077
rect 30932 3068 30984 3120
rect 10508 3000 10560 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 12808 2932 12860 2984
rect 7288 2864 7340 2916
rect 7472 2864 7524 2916
rect 8208 2864 8260 2916
rect 6828 2796 6880 2848
rect 10416 2796 10468 2848
rect 12348 2864 12400 2916
rect 14096 2932 14148 2984
rect 21272 3000 21324 3052
rect 15292 2932 15344 2984
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 7380 2592 7432 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 11888 2592 11940 2644
rect 11244 2456 11296 2508
rect 14924 2592 14976 2644
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 29644 2320 29696 2372
rect 11888 2252 11940 2304
rect 12900 2252 12952 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 2504 280 2556 332
rect 7012 280 7064 332
rect 15660 76 15712 128
rect 20628 76 20680 128
<< metal2 >>
rect 1214 15586 1270 16000
rect 3698 15586 3754 16000
rect 6182 15586 6238 16000
rect 8666 15586 8722 16000
rect 1214 15558 1624 15586
rect 1214 15520 1270 15558
rect 110 14376 166 14385
rect 110 14311 166 14320
rect 124 13190 152 14311
rect 112 13184 164 13190
rect 18 13152 74 13161
rect 112 13126 164 13132
rect 18 13087 74 13096
rect 32 12374 60 13087
rect 20 12368 72 12374
rect 20 12310 72 12316
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 112 10464 164 10470
rect 112 10406 164 10412
rect 124 9761 152 10406
rect 110 9752 166 9761
rect 110 9687 166 9696
rect 110 8664 166 8673
rect 110 8599 166 8608
rect 124 8401 152 8599
rect 110 8392 166 8401
rect 110 8327 166 8336
rect 1412 6866 1440 11086
rect 1596 10742 1624 15558
rect 3436 15558 3754 15586
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 2056 11218 2084 11766
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2240 11676 2268 12038
rect 2332 11830 2360 12242
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2792 11762 2820 12718
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11830 2912 12174
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2320 11688 2372 11694
rect 2240 11648 2320 11676
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1584 10736 1636 10742
rect 1688 10713 1716 10950
rect 1584 10678 1636 10684
rect 1674 10704 1730 10713
rect 1596 10452 1624 10678
rect 1674 10639 1730 10648
rect 1688 10606 1716 10639
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1780 10470 1808 11154
rect 2056 10810 2084 11154
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10606 2176 11630
rect 2240 11218 2268 11648
rect 2320 11630 2372 11636
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 1768 10464 1820 10470
rect 1596 10424 1716 10452
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1596 8634 1624 10231
rect 1688 10130 1716 10424
rect 1768 10406 1820 10412
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9586 1716 10066
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1688 9178 1716 9522
rect 1780 9382 1808 10406
rect 2148 9654 2176 10542
rect 2240 10198 2268 11154
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1582 6896 1638 6905
rect 1400 6860 1452 6866
rect 1780 6882 1808 9318
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1964 8090 1992 9046
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1872 7002 1900 7958
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1780 6854 1900 6882
rect 1582 6831 1638 6840
rect 1400 6802 1452 6808
rect 1412 5914 1440 6802
rect 1596 6458 1624 6831
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1780 5914 1808 6598
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1872 5778 1900 6854
rect 2044 6248 2096 6254
rect 2042 6216 2044 6225
rect 2096 6216 2098 6225
rect 2042 6151 2098 6160
rect 2056 6118 2084 6151
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1596 4282 1624 4655
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1398 82 1454 480
rect 1688 82 1716 5034
rect 1872 5030 1900 5714
rect 2148 5642 2176 9590
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2332 7954 2360 8978
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 7857 2360 7890
rect 2318 7848 2374 7857
rect 2318 7783 2320 7792
rect 2372 7783 2374 7792
rect 2320 7754 2372 7760
rect 2332 7723 2360 7754
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 6662 2268 7278
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2240 5030 2268 6598
rect 2424 6338 2452 8230
rect 2516 8022 2544 11086
rect 2884 11014 2912 11494
rect 3160 11121 3188 12582
rect 3436 12306 3464 15558
rect 3698 15520 3754 15558
rect 6104 15558 6238 15586
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3146 11112 3202 11121
rect 3068 11070 3146 11098
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10606 2912 10950
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2976 10266 3004 10678
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2976 9722 3004 10202
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2516 6458 2544 6870
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2424 6310 2544 6338
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2424 5681 2452 5850
rect 2410 5672 2466 5681
rect 2410 5607 2466 5616
rect 2424 5166 2452 5607
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 1872 1193 1900 4966
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3777 2452 3878
rect 2410 3768 2466 3777
rect 2410 3703 2466 3712
rect 2424 3602 2452 3703
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2424 3194 2452 3538
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 1858 1184 1914 1193
rect 1858 1119 1914 1128
rect 2516 338 2544 6310
rect 2608 5273 2636 9318
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8090 2728 8366
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 3068 8022 3096 11070
rect 3146 11047 3202 11056
rect 3528 10674 3556 11494
rect 3712 11354 3740 11766
rect 3804 11694 3832 12038
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4068 11552 4120 11558
rect 3804 11512 4068 11540
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 9042 3556 9386
rect 3804 9110 3832 11512
rect 4068 11494 4120 11500
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3988 9178 4016 10678
rect 4080 10470 4108 11154
rect 4264 11082 4292 11290
rect 4448 11218 4476 11630
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4264 10266 4292 11018
rect 4448 10810 4476 11154
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4632 10674 4660 11562
rect 5000 11558 5028 12242
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 10266 4844 10610
rect 4908 10538 4936 10950
rect 5000 10742 5028 11494
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 5276 10674 5304 11494
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10266 4936 10474
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9382 4752 10066
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9586 4936 9998
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3160 8498 3188 8910
rect 3528 8634 3556 8978
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7546 3004 7890
rect 3068 7546 3096 7958
rect 3528 7954 3556 8570
rect 3896 8566 3924 9046
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3976 8832 4028 8838
rect 4172 8820 4200 8910
rect 4028 8792 4200 8820
rect 3976 8774 4028 8780
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 8022 3648 8230
rect 3896 8090 3924 8502
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 2964 7540 3016 7546
rect 2884 7500 2964 7528
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6322 2728 6598
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2594 5264 2650 5273
rect 2594 5199 2650 5208
rect 2608 4690 2636 5199
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 4282 2636 4626
rect 2700 4282 2728 6258
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2792 5137 2820 5743
rect 2884 5370 2912 7500
rect 2964 7482 3016 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2884 5166 2912 5306
rect 2872 5160 2924 5166
rect 2778 5128 2834 5137
rect 2872 5102 2924 5108
rect 2778 5063 2834 5072
rect 2884 4826 2912 5102
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2884 3738 2912 4762
rect 2976 4758 3004 7278
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6458 3188 7142
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3054 6216 3110 6225
rect 3160 6186 3188 6394
rect 3054 6151 3110 6160
rect 3148 6180 3200 6186
rect 2964 4752 3016 4758
rect 2964 4694 3016 4700
rect 3068 4282 3096 6151
rect 3148 6122 3200 6128
rect 3160 5914 3188 6122
rect 3620 5914 3648 6734
rect 3804 6662 3832 6938
rect 3988 6730 4016 8774
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7002 4200 7822
rect 4264 7546 4292 7958
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 7274 4384 8230
rect 4448 8090 4476 8366
rect 4724 8362 4752 9318
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4816 8022 4844 9046
rect 5184 8838 5212 9454
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 4804 8016 4856 8022
rect 5184 7993 5212 8774
rect 4804 7958 4856 7964
rect 5170 7984 5226 7993
rect 5170 7919 5226 7928
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6322 3832 6598
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 4172 5914 4200 6734
rect 4264 6390 4292 6870
rect 4356 6644 4384 7210
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4448 6798 4476 6938
rect 4908 6934 4936 7142
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4356 6616 4476 6644
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4356 6186 4384 6394
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 3620 3670 3648 5850
rect 4264 5574 4292 6122
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3974 5128 4030 5137
rect 3974 5063 4030 5072
rect 3988 4146 4016 5063
rect 4264 4282 4292 5510
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 2504 332 2556 338
rect 2504 274 2556 280
rect 1398 54 1716 82
rect 4250 82 4306 480
rect 4448 82 4476 6616
rect 4816 6390 4844 6666
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5846 5212 6054
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5000 5302 5028 5714
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5184 5234 5212 5782
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5368 4690 5396 8774
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5552 7886 5580 8502
rect 5736 8362 5764 8978
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6458 5672 6802
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5644 5914 5672 6394
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5460 5370 5488 5714
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5460 4758 5488 5306
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4908 4282 4936 4626
rect 5644 4282 5672 5850
rect 5828 5302 5856 11494
rect 6104 7954 6132 15558
rect 6182 15520 6238 15558
rect 8404 15558 8722 15586
rect 7194 14920 7250 14929
rect 7194 14855 7250 14864
rect 7208 12986 7236 14855
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 6564 11626 6592 12242
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6748 11218 6776 12038
rect 7484 11665 7512 12242
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7656 11688 7708 11694
rect 7470 11656 7526 11665
rect 7656 11630 7708 11636
rect 7470 11591 7526 11600
rect 7484 11558 7512 11591
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7668 11354 7696 11630
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 8128 11286 8156 12038
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6748 10742 6776 11154
rect 6932 10810 6960 11154
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 8022 10840 8078 10849
rect 6920 10804 6972 10810
rect 8022 10775 8078 10784
rect 6920 10746 6972 10752
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6932 9518 6960 10746
rect 8036 10742 8064 10775
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7024 9382 7052 10406
rect 7760 10266 7788 10542
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7944 10266 7972 10474
rect 8128 10266 8156 11222
rect 8312 10810 8340 11562
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7932 10260 7984 10266
rect 8116 10260 8168 10266
rect 7984 10220 8064 10248
rect 7932 10202 7984 10208
rect 7116 9382 7144 10202
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9518 7236 9862
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7208 9042 7236 9454
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 7196 9036 7248 9042
rect 7392 9024 7420 9386
rect 7484 9178 7512 9998
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7472 9036 7524 9042
rect 7392 8996 7472 9024
rect 7196 8978 7248 8984
rect 7472 8978 7524 8984
rect 6196 8294 6224 8978
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7024 8401 7052 8570
rect 7010 8392 7066 8401
rect 7208 8362 7236 8978
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7010 8327 7066 8336
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6104 7478 6132 7890
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6196 7002 6224 8230
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 6118 6132 6802
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5552 3369 5580 4014
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5920 3602 5948 3946
rect 6012 3738 6040 4694
rect 6104 4690 6132 6054
rect 6196 4826 6224 6938
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6104 4078 6132 4626
rect 6380 4282 6408 6734
rect 6472 4554 6500 7414
rect 6656 5710 6684 8230
rect 7208 8090 7236 8298
rect 7300 8294 7328 8910
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6564 3738 6592 5510
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 6380 3194 6408 3538
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6840 2854 6868 8026
rect 7484 7954 7512 8978
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8036 8634 8064 10220
rect 8116 10202 8168 10208
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8401 7696 8434
rect 7654 8392 7710 8401
rect 8036 8362 8064 8570
rect 7654 8327 7710 8336
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 6934 6960 7822
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7206 7236 7754
rect 7484 7750 7512 7890
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6932 6254 6960 6870
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6390 7052 6598
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5914 6960 6190
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 4826 7052 6326
rect 7208 6322 7236 7142
rect 7484 6662 7512 7686
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 7932 7472 7984 7478
rect 8036 7460 8064 7686
rect 7984 7432 8064 7460
rect 7932 7414 7984 7420
rect 8128 7410 8156 7822
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 7002 7696 7210
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 5846 7144 6190
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 5234 7236 5646
rect 7300 5370 7328 6054
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 3738 6960 4626
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7024 4078 7052 4218
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7208 4010 7236 5034
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7300 4154 7328 4762
rect 7392 4690 7420 5782
rect 7484 5710 7512 6598
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8036 6458 8064 6802
rect 8128 6798 8156 7346
rect 8220 7342 8248 9522
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7585 8340 7686
rect 8298 7576 8354 7585
rect 8298 7511 8354 7520
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8036 5098 8064 5714
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5166 8156 5646
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4758 8064 5034
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7300 4126 7420 4154
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7208 3738 7236 3946
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7392 3466 7420 4126
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7300 2922 7328 3334
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 7010 2680 7066 2689
rect 7392 2650 7420 3402
rect 7484 3194 7512 4558
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8036 4282 8064 4490
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7760 3670 7788 4014
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 8036 3466 8064 4218
rect 8114 3496 8170 3505
rect 8024 3460 8076 3466
rect 8114 3431 8170 3440
rect 8024 3402 8076 3408
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8036 3194 8064 3402
rect 8128 3398 8156 3431
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8220 2922 8248 6054
rect 8404 5914 8432 15558
rect 8666 15520 8722 15558
rect 11150 15632 11206 16000
rect 11150 15580 11152 15632
rect 11204 15580 11206 15632
rect 13634 15586 13690 16000
rect 11150 15520 11206 15580
rect 13372 15558 13690 15586
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11762 8616 12174
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8496 9178 8524 11086
rect 8680 10470 8708 12582
rect 8956 11898 8984 12582
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8956 11558 8984 11834
rect 10428 11762 10456 12718
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10612 11898 10640 12106
rect 10600 11892 10652 11898
rect 10652 11852 10732 11880
rect 10600 11834 10652 11840
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9232 11354 9260 11698
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 10428 11286 10456 11698
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 8956 10742 8984 11222
rect 9876 10810 9904 11222
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8956 10130 8984 10678
rect 9876 10470 9904 10746
rect 10152 10742 10180 11086
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 10152 10266 10180 10678
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8496 8498 8524 9114
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8588 8378 8616 9454
rect 9048 9382 9076 10066
rect 10244 9722 10272 10542
rect 10612 10470 10640 10610
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 8496 8350 8616 8378
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8496 5778 8524 8350
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8588 7546 8616 8230
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6730 8708 7278
rect 8772 6934 8800 7686
rect 8864 7274 8892 7822
rect 9048 7546 9076 9318
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9140 8362 9168 8570
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8312 5166 8340 5238
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8496 4486 8524 5714
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 2961 8340 3878
rect 8588 3720 8616 6598
rect 8680 6118 8708 6666
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5846 8708 6054
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 4826 8708 5646
rect 9140 5370 9168 8298
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7478 9352 7686
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9220 7404 9272 7410
rect 9588 7404 9640 7410
rect 9220 7346 9272 7352
rect 9416 7364 9588 7392
rect 9232 7313 9260 7346
rect 9218 7304 9274 7313
rect 9218 7239 9274 7248
rect 9416 6798 9444 7364
rect 9588 7346 9640 7352
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6458 9444 6734
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 5914 9536 6938
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9140 5098 9168 5306
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8680 4146 8708 4762
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9140 4010 9168 5034
rect 9416 4826 9444 5102
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8588 3692 8708 3720
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8496 3194 8524 3606
rect 8680 3233 8708 3692
rect 8666 3224 8722 3233
rect 8484 3188 8536 3194
rect 9784 3194 9812 9318
rect 9968 6984 9996 9590
rect 10704 9518 10732 11852
rect 10980 11558 11008 12242
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10980 11014 11008 11494
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 9926 11008 10950
rect 11072 10266 11100 12174
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11164 11121 11192 11630
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11150 11112 11206 11121
rect 11150 11047 11206 11056
rect 11164 11014 11192 11047
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11532 10674 11560 11562
rect 11900 11150 11928 13262
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12442 12388 13126
rect 13372 12986 13400 15558
rect 13634 15520 13690 15558
rect 15476 15564 15528 15570
rect 16210 15564 16266 16000
rect 16210 15520 16212 15564
rect 15476 15506 15528 15512
rect 16264 15520 16266 15564
rect 18694 15586 18750 16000
rect 19156 15632 19208 15638
rect 18694 15558 18828 15586
rect 19156 15574 19208 15580
rect 21178 15586 21234 16000
rect 23662 15586 23718 16000
rect 26146 15586 26202 16000
rect 18694 15520 18750 15558
rect 16212 15506 16264 15512
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12084 11762 12112 12242
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12544 11626 12572 12038
rect 13096 11830 13124 12242
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12544 11354 12572 11562
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10266 11376 10406
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9518 11008 9862
rect 11348 9586 11376 10202
rect 11900 10130 11928 11086
rect 11992 10538 12020 11222
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 10266 12020 10474
rect 12544 10266 12572 10610
rect 12636 10266 12664 11562
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10704 9178 10732 9454
rect 11348 9382 11376 9522
rect 11532 9382 11560 9998
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10888 8974 10916 9318
rect 10980 9110 11008 9318
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8634 10916 8910
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10980 8566 11008 9046
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10060 8022 10088 8298
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10966 7848 11022 7857
rect 10152 7002 10180 7822
rect 10140 6996 10192 7002
rect 9968 6956 10088 6984
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9968 6118 9996 6802
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5574 9996 6054
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5302 9996 5510
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 8666 3159 8722 3168
rect 9772 3188 9824 3194
rect 8484 3130 8536 3136
rect 9772 3130 9824 3136
rect 8298 2952 8354 2961
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 8208 2916 8260 2922
rect 8298 2887 8354 2896
rect 8208 2858 8260 2864
rect 7010 2615 7066 2624
rect 7380 2644 7432 2650
rect 7024 338 7052 2615
rect 7380 2586 7432 2592
rect 7484 2281 7512 2858
rect 7470 2272 7526 2281
rect 7470 2207 7526 2216
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 7012 332 7064 338
rect 7012 274 7064 280
rect 4250 54 4476 82
rect 7024 82 7052 274
rect 7102 82 7158 480
rect 7024 54 7158 82
rect 1398 0 1454 54
rect 4250 0 4306 54
rect 7102 0 7158 54
rect 9954 82 10010 480
rect 10060 82 10088 6956
rect 10140 6938 10192 6944
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 5846 10180 6598
rect 10336 6390 10364 7822
rect 11164 7834 11192 8298
rect 11022 7806 11192 7834
rect 10966 7783 11022 7792
rect 10980 7750 11008 7783
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 6934 10916 7278
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10796 5846 10824 6122
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10152 5370 10180 5782
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10244 5098 10272 5646
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4826 10272 5034
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10796 4622 10824 5782
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10784 4616 10836 4622
rect 10704 4576 10784 4604
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10520 3058 10548 3946
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10704 3738 10732 4576
rect 10784 4558 10836 4564
rect 10784 4208 10836 4214
rect 10784 4154 10836 4156
rect 10888 4154 10916 4694
rect 10784 4150 10916 4154
rect 10796 4126 10916 4150
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10796 3602 10824 4126
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10796 3194 10824 3538
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11072 3126 11100 7686
rect 11164 7342 11192 7806
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11256 6866 11284 7482
rect 11532 7410 11560 9318
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11808 8634 11836 8978
rect 12176 8634 12204 9386
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 8022 12112 8502
rect 12636 8090 12664 8842
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 12254 7984 12310 7993
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11624 6934 11652 7890
rect 11808 7410 11836 7890
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6322 11192 6598
rect 11256 6322 11284 6802
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11164 5914 11192 6258
rect 11256 6225 11284 6258
rect 11242 6216 11298 6225
rect 11242 6151 11298 6160
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11612 5772 11664 5778
rect 11716 5760 11744 7142
rect 11808 6798 11836 7346
rect 12084 7206 12112 7958
rect 12254 7919 12310 7928
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 6934 12112 7142
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 12084 6458 12112 6870
rect 12176 6662 12204 7278
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12084 6186 12112 6394
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12084 5914 12112 6122
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11796 5772 11848 5778
rect 11716 5732 11796 5760
rect 11612 5714 11664 5720
rect 11796 5714 11848 5720
rect 11624 5370 11652 5714
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11624 4826 11652 5306
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 11256 4146 11284 4490
rect 11716 4282 11744 4966
rect 11808 4826 11836 5714
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10428 2650 10456 2790
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 11256 2514 11284 4082
rect 11716 3777 11744 4218
rect 11702 3768 11758 3777
rect 11702 3703 11758 3712
rect 11900 2650 11928 5510
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4826 12112 5102
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12176 3738 12204 6598
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12268 3602 12296 7919
rect 12728 4826 12756 8298
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 4282 12480 4626
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12728 4078 12756 4762
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3602 12388 3878
rect 12820 3738 12848 11766
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13188 11082 13216 11562
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13004 9722 13032 10134
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13280 8906 13308 12786
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 10849 13400 12718
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13358 10840 13414 10849
rect 13358 10775 13414 10784
rect 13372 9518 13400 10775
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13372 8430 13400 9114
rect 13464 8634 13492 12038
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13556 10810 13584 11222
rect 13636 11144 13688 11150
rect 13740 11132 13768 11766
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 13688 11104 13768 11132
rect 13636 11086 13688 11092
rect 13634 10840 13690 10849
rect 13544 10804 13596 10810
rect 13634 10775 13690 10784
rect 13544 10746 13596 10752
rect 13648 10606 13676 10775
rect 13740 10742 13768 11104
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9654 13768 9862
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 8022 13584 8366
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7274 12940 7822
rect 13740 7478 13768 9590
rect 14200 9586 14228 10610
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14096 9444 14148 9450
rect 14096 9386 14148 9392
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 4214 12940 7210
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 5574 13032 6734
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5846 13216 6054
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12268 3194 12296 3538
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12360 2922 12388 3538
rect 12820 2990 12848 3674
rect 13004 3058 13032 5510
rect 13096 4826 13124 5646
rect 13188 5370 13216 5782
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13096 3194 13124 4762
rect 13280 4758 13308 6598
rect 13372 6458 13400 7142
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13188 3738 13216 4490
rect 13280 4282 13308 4694
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13372 4146 13400 6190
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13464 3738 13492 5510
rect 13648 5234 13676 5578
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13740 5234 13768 5306
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13648 4554 13676 5170
rect 13832 5098 13860 7686
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13924 4758 13952 5170
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 14016 4078 14044 9318
rect 14108 5273 14136 9386
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14660 9178 14688 9318
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14200 8566 14228 8978
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6322 14320 6802
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14384 6186 14412 6394
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5914 14228 6054
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14200 5574 14228 5850
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14094 5264 14150 5273
rect 14660 5234 14688 6258
rect 14094 5199 14150 5208
rect 14648 5228 14700 5234
rect 14108 4214 14136 5199
rect 14648 5170 14700 5176
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14752 4468 14780 10406
rect 14936 8401 14964 11630
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14922 8392 14978 8401
rect 14922 8327 14978 8336
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14844 5370 14872 5646
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14844 4826 14872 5306
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 5137 14964 5170
rect 14922 5128 14978 5137
rect 14922 5063 14978 5072
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14924 4480 14976 4486
rect 14752 4440 14924 4468
rect 14924 4422 14976 4428
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14016 3738 14044 4014
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 14108 2689 14136 2926
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14094 2680 14150 2689
rect 11888 2644 11940 2650
rect 14289 2672 14585 2692
rect 14936 2650 14964 4422
rect 15028 4146 15056 11494
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15304 10742 15332 11154
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15212 8838 15240 9998
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15120 8022 15148 8366
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15212 7410 15240 8774
rect 15304 8362 15332 8910
rect 15396 8498 15424 9454
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15304 8090 15332 8298
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15488 7546 15516 15506
rect 16224 15475 16252 15506
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12714 15884 13126
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15580 11694 15608 12378
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15764 7954 15792 12582
rect 15856 11898 15884 12650
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16132 11558 16160 12174
rect 16224 11898 16252 12310
rect 16684 12170 16712 12786
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10538 15884 10950
rect 16132 10810 16160 11494
rect 16224 11286 16252 11834
rect 16500 11626 16528 12106
rect 16684 11830 16712 12106
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 16304 11620 16356 11626
rect 16304 11562 16356 11568
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16224 10810 16252 11222
rect 16316 11218 16344 11562
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16316 10606 16344 11154
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15856 10266 15884 10474
rect 16316 10266 16344 10542
rect 16592 10266 16620 11086
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 15856 9722 15884 10202
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 16684 9518 16712 9862
rect 17236 9586 17264 9998
rect 17604 9722 17632 10202
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16028 9444 16080 9450
rect 15948 9404 16028 9432
rect 15948 9110 15976 9404
rect 16028 9386 16080 9392
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 15948 8362 15976 9046
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8498 16528 8774
rect 17512 8634 17540 9046
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 8634 17632 8910
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7546 15792 7890
rect 15476 7540 15528 7546
rect 15752 7540 15804 7546
rect 15528 7500 15608 7528
rect 15476 7482 15528 7488
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15120 6662 15148 7278
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15120 5370 15148 5782
rect 15488 5681 15516 6598
rect 15474 5672 15530 5681
rect 15474 5607 15530 5616
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 15028 3641 15056 4082
rect 15304 4078 15332 4150
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15014 3632 15070 3641
rect 15014 3567 15070 3576
rect 15304 2990 15332 4014
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 14094 2615 14150 2624
rect 14924 2644 14976 2650
rect 11888 2586 11940 2592
rect 14924 2586 14976 2592
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 11900 105 11928 2246
rect 9954 54 10088 82
rect 11886 96 11942 105
rect 9954 0 10010 54
rect 11886 31 11942 40
rect 12806 82 12862 480
rect 12912 82 12940 2246
rect 15396 1873 15424 5238
rect 15488 4690 15516 5607
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4214 15516 4626
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15488 3602 15516 4150
rect 15580 3602 15608 7500
rect 15752 7482 15804 7488
rect 15948 6916 15976 8298
rect 16500 8022 16528 8434
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16670 7440 16726 7449
rect 16670 7375 16726 7384
rect 16684 7342 16712 7375
rect 16868 7342 16896 7890
rect 17144 7410 17172 8366
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16868 7002 16896 7278
rect 17328 7206 17356 7890
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16028 6928 16080 6934
rect 15948 6888 16028 6916
rect 15948 6458 15976 6888
rect 16028 6870 16080 6876
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 5234 15700 5646
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 4622 15700 5170
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15764 3738 15792 6258
rect 15948 6186 15976 6394
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16316 5574 16344 6734
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 4554 15884 5102
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15948 4154 15976 4626
rect 15948 4126 16068 4154
rect 16316 4146 16344 5510
rect 16592 5098 16620 6598
rect 16868 6458 16896 6938
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16684 5574 16712 6190
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5846 16988 6054
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16500 4826 16528 5034
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16040 4078 16068 4126
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16040 3738 16068 4014
rect 16500 3738 16528 4762
rect 16684 4758 16712 5510
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 17236 4282 17264 5034
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 15488 3194 15516 3538
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 16776 3126 16804 3538
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 17328 2961 17356 7142
rect 17696 6866 17724 11630
rect 18248 11286 18276 12582
rect 18800 12442 18828 15558
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 19168 11354 19196 15574
rect 21178 15558 21312 15586
rect 21178 15520 21234 15558
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 11558 19288 11698
rect 19536 11694 19564 12242
rect 19812 12102 19840 12582
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18248 10810 18276 11222
rect 18236 10804 18288 10810
rect 18236 10746 18288 10752
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18156 10266 18184 10474
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18248 10130 18276 10746
rect 18708 10742 18736 11290
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10810 19104 11086
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9654 18460 9862
rect 18800 9722 18828 10202
rect 19260 10062 19288 11494
rect 19812 11393 19840 11494
rect 19798 11384 19854 11393
rect 19798 11319 19854 11328
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19536 10742 19564 11018
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18432 9450 18460 9590
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18156 8906 18184 9386
rect 18524 8974 18552 9522
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 19076 8838 19104 9998
rect 19352 9654 19380 10066
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19352 9382 19380 9590
rect 19996 9586 20024 9998
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18616 8430 18644 8774
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 8022 18644 8230
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 17774 7576 17830 7585
rect 17774 7511 17830 7520
rect 18052 7540 18104 7546
rect 17788 7478 17816 7511
rect 18052 7482 18104 7488
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17958 7440 18014 7449
rect 17958 7375 18014 7384
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6322 17908 6802
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17420 5370 17448 5782
rect 17972 5370 18000 7375
rect 18064 5846 18092 7482
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6186 18276 6598
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18156 5914 18184 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17420 4758 17448 5306
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 4146 17448 4694
rect 17604 4622 17632 5170
rect 17972 5166 18000 5306
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17512 4282 17540 4558
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17696 3194 17724 5102
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17314 2952 17370 2961
rect 17314 2887 17370 2896
rect 15382 1864 15438 1873
rect 15382 1799 15438 1808
rect 12806 54 12940 82
rect 15658 128 15714 480
rect 15658 76 15660 128
rect 15712 76 15714 128
rect 12806 0 12862 54
rect 15658 0 15714 76
rect 18248 82 18276 5238
rect 18340 4282 18368 5646
rect 18432 5642 18460 6258
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18524 5166 18552 7686
rect 18616 7410 18644 7958
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18708 6934 18736 7822
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18800 6662 18828 7278
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4826 18552 5102
rect 18616 4826 18644 5850
rect 18800 5234 18828 6598
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18786 4720 18842 4729
rect 18786 4655 18788 4664
rect 18840 4655 18842 4664
rect 18788 4626 18840 4632
rect 18800 4486 18828 4626
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18800 4146 18828 4422
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 2553 18644 3878
rect 18892 3738 18920 7754
rect 19076 7546 19104 8774
rect 19444 8498 19472 9046
rect 20088 8974 20116 13126
rect 20456 12782 20484 13262
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 11762 20484 12718
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20444 11756 20496 11762
rect 20496 11716 20576 11744
rect 20444 11698 20496 11704
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20456 10674 20484 11562
rect 20548 11354 20576 11716
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20456 10266 20484 10610
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20732 10130 20760 12650
rect 20824 12646 20852 13330
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 10849 20852 12582
rect 21284 12374 21312 15558
rect 23662 15558 23796 15586
rect 23662 15520 23718 15558
rect 23768 12986 23796 15558
rect 25792 15558 26202 15586
rect 25792 12986 25820 15558
rect 26146 15520 26202 15558
rect 27988 15564 28040 15570
rect 28722 15564 28778 16000
rect 28722 15520 28724 15564
rect 27988 15506 28040 15512
rect 28776 15520 28778 15564
rect 31206 15586 31262 16000
rect 33690 15586 33746 16000
rect 36174 15586 36230 16000
rect 31206 15558 31340 15586
rect 31206 15520 31262 15558
rect 28724 15506 28776 15512
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 21284 11898 21312 12174
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20810 10840 20866 10849
rect 20956 10832 21252 10852
rect 20810 10775 20866 10784
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20824 10033 20852 10775
rect 21468 10606 21496 12718
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 21916 12164 21968 12170
rect 21916 12106 21968 12112
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21560 11014 21588 11562
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21560 10810 21588 10950
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21284 10266 21312 10474
rect 21652 10470 21680 11222
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 20810 10024 20866 10033
rect 20810 9959 20866 9968
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21284 9450 21312 10202
rect 21652 9722 21680 10406
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 20088 8022 20116 8910
rect 21284 8838 21312 9386
rect 21468 9178 21496 9522
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 8022 20300 8230
rect 20076 8016 20128 8022
rect 20076 7958 20128 7964
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7546 20300 7958
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20364 7002 20392 7822
rect 20456 7818 20484 8298
rect 20548 8022 20576 8298
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 7410 21312 8774
rect 21376 8634 21404 8774
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21744 8362 21772 12038
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21836 10810 21864 11086
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21928 10248 21956 12106
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22020 11150 22048 11562
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21836 10220 21956 10248
rect 21836 8974 21864 10220
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21928 9722 21956 10066
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21836 8634 21864 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21928 8566 21956 9046
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19260 5778 19288 6326
rect 19812 6118 19840 6802
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6186 20576 6598
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19260 5370 19288 5714
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19720 5370 19748 5646
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19720 5166 19748 5306
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19812 4690 19840 6054
rect 20548 5370 20576 6122
rect 20640 5846 20668 6734
rect 20824 6662 20852 7210
rect 21284 7002 21312 7346
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6458 20852 6598
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20812 6452 20864 6458
rect 21284 6440 21312 6938
rect 21376 6934 21404 8298
rect 21744 7954 21772 8298
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21928 8022 21956 8230
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21836 7274 21864 7822
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21744 7002 21772 7142
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 20812 6394 20864 6400
rect 21192 6412 21312 6440
rect 21192 5846 21220 6412
rect 21376 6322 21404 6870
rect 21744 6458 21772 6938
rect 21836 6730 21864 7210
rect 22020 7206 22048 7822
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20824 5370 20852 5714
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 19800 4684 19852 4690
rect 19800 4626 19852 4632
rect 19812 4282 19840 4626
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19168 3738 19196 4014
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18602 2544 18658 2553
rect 18602 2479 18658 2488
rect 18510 82 18566 480
rect 20640 134 20668 5238
rect 21284 4690 21312 6258
rect 21744 6118 21772 6394
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 21928 5370 21956 5782
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4146 21312 4626
rect 21376 4154 21404 5034
rect 22020 4758 22048 7142
rect 22112 5234 22140 11562
rect 22296 11558 22324 12242
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 10713 22324 11494
rect 22282 10704 22338 10713
rect 22282 10639 22338 10648
rect 22296 9489 22324 10639
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22282 9480 22338 9489
rect 22282 9415 22338 9424
rect 22388 7426 22416 10542
rect 22836 10192 22888 10198
rect 22836 10134 22888 10140
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9722 22784 9998
rect 22848 9722 22876 10134
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8566 22600 8774
rect 22940 8634 22968 12038
rect 23032 11626 23060 12242
rect 23020 11620 23072 11626
rect 23072 11580 23152 11608
rect 23020 11562 23072 11568
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23032 10062 23060 11086
rect 23124 10985 23152 11580
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23110 10976 23166 10985
rect 23110 10911 23166 10920
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22480 7546 22508 8026
rect 22572 7868 22600 8502
rect 22652 7880 22704 7886
rect 22572 7840 22652 7868
rect 22652 7822 22704 7828
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22388 7398 22508 7426
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22388 6118 22416 6734
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22204 5098 22232 5510
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 22112 4826 22140 5034
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22204 4690 22232 5034
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22388 4282 22416 6054
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 21272 4140 21324 4146
rect 21376 4126 21496 4154
rect 21272 4082 21324 4088
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 3233 20760 4014
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20718 3224 20774 3233
rect 20956 3216 21252 3236
rect 20718 3159 20774 3168
rect 21284 3058 21312 4082
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 18248 54 18566 82
rect 20628 128 20680 134
rect 20628 70 20680 76
rect 21362 82 21418 480
rect 21468 82 21496 4126
rect 22480 4078 22508 7398
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22756 5778 22784 6938
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22848 6186 22876 6802
rect 23124 6769 23152 9318
rect 23216 8090 23244 11494
rect 23308 11218 23336 12378
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24136 11665 24164 11698
rect 24122 11656 24178 11665
rect 24122 11591 24178 11600
rect 24214 11384 24270 11393
rect 24214 11319 24270 11328
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23584 10674 23612 10950
rect 23952 10713 23980 11154
rect 23938 10704 23994 10713
rect 23572 10668 23624 10674
rect 23938 10639 23994 10648
rect 23572 10610 23624 10616
rect 23584 10545 23612 10610
rect 23952 10606 23980 10639
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24136 10266 24164 10542
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24136 9926 24164 10202
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 23400 9602 23428 9862
rect 23662 9752 23718 9761
rect 23662 9687 23718 9696
rect 23676 9654 23704 9687
rect 23664 9648 23716 9654
rect 23400 9574 23520 9602
rect 23664 9590 23716 9596
rect 23492 9160 23520 9574
rect 24228 9178 24256 11319
rect 24412 9654 24440 12718
rect 24504 11898 24532 12786
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24504 11694 24532 11834
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24688 11676 24716 12038
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24768 11688 24820 11694
rect 24688 11648 24768 11676
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10266 24624 10542
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24412 9518 24440 9590
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24216 9172 24268 9178
rect 23492 9132 23612 9160
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23492 8566 23520 8978
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23216 7546 23244 8026
rect 23492 7993 23520 8502
rect 23478 7984 23534 7993
rect 23478 7919 23534 7928
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23584 7449 23612 9132
rect 24216 9114 24268 9120
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24044 8498 24072 8910
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23768 8022 23796 8298
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 24044 7818 24072 8434
rect 24032 7812 24084 7818
rect 24032 7754 24084 7760
rect 23570 7440 23626 7449
rect 23570 7375 23626 7384
rect 23110 6760 23166 6769
rect 23110 6695 23166 6704
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5914 22968 6054
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 23032 4554 23060 6190
rect 23124 4690 23152 6695
rect 23584 6390 23612 7375
rect 24136 7206 24164 8774
rect 24596 8430 24624 9522
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24412 8022 24440 8230
rect 24400 8016 24452 8022
rect 24400 7958 24452 7964
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23860 6254 23888 6598
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23952 6186 23980 7142
rect 24412 7002 24440 7958
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 24136 6254 24164 6734
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23308 5370 23336 5782
rect 23768 5778 23796 6054
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23216 4826 23244 5170
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23768 4758 23796 5714
rect 24688 5710 24716 11648
rect 24768 11630 24820 11636
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24780 10470 24808 11154
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24780 9450 24808 9930
rect 24872 9586 24900 10474
rect 24964 9722 24992 10474
rect 25044 10192 25096 10198
rect 25044 10134 25096 10140
rect 25056 9722 25084 10134
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24768 9444 24820 9450
rect 24768 9386 24820 9392
rect 24872 9178 24900 9522
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 9178 25084 9318
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25056 8362 25084 9114
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23860 4826 23888 5034
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 24136 4758 24164 5510
rect 24412 5234 24440 5510
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23020 4548 23072 4554
rect 23020 4490 23072 4496
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 23032 3738 23060 4490
rect 23124 3942 23152 4626
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24044 4282 24072 4558
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 18510 0 18566 54
rect 21362 54 21496 82
rect 24044 82 24072 3878
rect 24136 3738 24164 4694
rect 24412 4622 24440 5034
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24688 4214 24716 5646
rect 24676 4208 24728 4214
rect 24676 4150 24728 4156
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24228 3670 24256 3878
rect 24688 3738 24716 4150
rect 24872 4078 24900 6122
rect 24964 5914 24992 6734
rect 25056 6458 25084 6870
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 25148 5778 25176 11766
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25240 10674 25268 10746
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25240 10062 25268 10610
rect 25332 10577 25360 12038
rect 26054 11792 26110 11801
rect 26054 11727 26110 11736
rect 26068 11694 26096 11727
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25318 10568 25374 10577
rect 25318 10503 25374 10512
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25332 6662 25360 10406
rect 25424 8498 25452 11562
rect 26238 11384 26294 11393
rect 26238 11319 26294 11328
rect 26252 11286 26280 11319
rect 26240 11280 26292 11286
rect 26240 11222 26292 11228
rect 26252 11082 26280 11222
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10538 25820 10950
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 9178 25636 10406
rect 25872 9988 25924 9994
rect 25872 9930 25924 9936
rect 25884 9178 25912 9930
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 26344 9042 26372 12310
rect 26436 11286 26464 12582
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26424 11280 26476 11286
rect 26424 11222 26476 11228
rect 26436 10266 26464 11222
rect 26528 10266 26556 12038
rect 26698 11792 26754 11801
rect 26698 11727 26754 11736
rect 26712 11694 26740 11727
rect 26700 11688 26752 11694
rect 26700 11630 26752 11636
rect 26608 11620 26660 11626
rect 26608 11562 26660 11568
rect 26976 11620 27028 11626
rect 26976 11562 27028 11568
rect 26620 11393 26648 11562
rect 26606 11384 26662 11393
rect 26606 11319 26662 11328
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26620 9586 26648 11086
rect 26712 10470 26740 11222
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26896 10810 26924 11086
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26712 10198 26740 10406
rect 26700 10192 26752 10198
rect 26700 10134 26752 10140
rect 26712 9654 26740 10134
rect 26896 9761 26924 10746
rect 26882 9752 26938 9761
rect 26882 9687 26938 9696
rect 26700 9648 26752 9654
rect 26700 9590 26752 9596
rect 26608 9580 26660 9586
rect 26608 9522 26660 9528
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26344 8634 26372 8978
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25424 8090 25452 8434
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26240 8288 26292 8294
rect 26240 8230 26292 8236
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 26252 8022 26280 8230
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 26332 7880 26384 7886
rect 26332 7822 26384 7828
rect 26344 7478 26372 7822
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25504 6248 25556 6254
rect 25504 6190 25556 6196
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 25148 5370 25176 5714
rect 25516 5574 25544 6190
rect 25608 6186 25636 7142
rect 26344 7002 26372 7414
rect 26332 6996 26384 7002
rect 26332 6938 26384 6944
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25608 5846 25636 6122
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25148 4729 25176 5306
rect 25332 5234 25360 5510
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 25332 4826 25360 5170
rect 25412 5092 25464 5098
rect 25412 5034 25464 5040
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 25424 4758 25452 5034
rect 25412 4752 25464 4758
rect 25134 4720 25190 4729
rect 25412 4694 25464 4700
rect 25134 4655 25190 4664
rect 25412 4208 25464 4214
rect 25412 4150 25464 4156
rect 25424 4078 25452 4150
rect 25516 4146 25544 5510
rect 26436 4282 26464 8366
rect 26528 8362 26556 9318
rect 26620 9024 26648 9522
rect 26712 9178 26740 9590
rect 26988 9178 27016 11562
rect 27448 11558 27476 12242
rect 28000 11830 28028 15506
rect 28736 15475 28764 15506
rect 31312 12714 31340 15558
rect 33336 15558 33746 15586
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 31300 12708 31352 12714
rect 31300 12650 31352 12656
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29104 12374 29132 12582
rect 29092 12368 29144 12374
rect 29092 12310 29144 12316
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 28092 11558 28120 12242
rect 29000 12096 29052 12102
rect 29000 12038 29052 12044
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27528 11552 27580 11558
rect 27528 11494 27580 11500
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27356 10266 27384 10610
rect 27448 10577 27476 11494
rect 27434 10568 27490 10577
rect 27434 10503 27490 10512
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26976 9172 27028 9178
rect 27028 9132 27108 9160
rect 26976 9114 27028 9120
rect 26700 9036 26752 9042
rect 26620 8996 26700 9024
rect 26700 8978 26752 8984
rect 26976 8832 27028 8838
rect 26976 8774 27028 8780
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 26804 7546 26832 7958
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26988 7410 27016 8774
rect 27080 8498 27108 9132
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26436 4154 26464 4218
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 26344 4126 26464 4154
rect 26344 4078 26372 4126
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 25412 4072 25464 4078
rect 25412 4014 25464 4020
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26620 3942 26648 7278
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26712 6934 26740 7142
rect 26700 6928 26752 6934
rect 26700 6870 26752 6876
rect 26712 5914 26740 6870
rect 27080 6186 27108 8230
rect 27264 7886 27292 8910
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27172 6458 27200 7142
rect 27264 6934 27292 7822
rect 27252 6928 27304 6934
rect 27252 6870 27304 6876
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27068 6180 27120 6186
rect 27120 6140 27200 6168
rect 27068 6122 27120 6128
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 27172 5846 27200 6140
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27160 5840 27212 5846
rect 27160 5782 27212 5788
rect 27172 5166 27200 5782
rect 27264 5778 27292 6054
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 27264 5370 27292 5714
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24214 82 24270 480
rect 24044 54 24270 82
rect 21362 0 21418 54
rect 24214 0 24270 54
rect 27066 82 27122 480
rect 27356 82 27384 9454
rect 27540 9110 27568 11494
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 27988 11348 28040 11354
rect 27988 11290 28040 11296
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 28000 10062 28028 11290
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 28000 9654 28028 9998
rect 27988 9648 28040 9654
rect 27988 9590 28040 9596
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27528 9104 27580 9110
rect 27528 9046 27580 9052
rect 27988 9104 28040 9110
rect 27988 9046 28040 9052
rect 27540 8634 27568 9046
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 28000 8294 28028 9046
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28000 8090 28028 8230
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 27448 6254 27476 7142
rect 27540 7002 27568 7346
rect 28092 7313 28120 11494
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28184 10470 28212 11154
rect 29012 11150 29040 12038
rect 31312 11898 31340 12650
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 30116 11218 30144 11834
rect 31312 11694 31340 11834
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31116 11552 31168 11558
rect 31116 11494 31168 11500
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30104 11212 30156 11218
rect 30104 11154 30156 11160
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28184 8974 28212 10406
rect 28264 10192 28316 10198
rect 28264 10134 28316 10140
rect 28276 9722 28304 10134
rect 28460 10062 28488 10610
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 29012 9722 29040 11086
rect 29828 11008 29880 11014
rect 29828 10950 29880 10956
rect 29840 10674 29868 10950
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 29012 8634 29040 9658
rect 29840 9586 29868 10610
rect 30116 10266 30144 11154
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29288 9178 29316 9454
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29012 8090 29040 8570
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 28078 7304 28134 7313
rect 28078 7239 28134 7248
rect 28920 7206 28948 7890
rect 29104 7546 29132 8366
rect 29932 8022 29960 8910
rect 30012 8424 30064 8430
rect 30012 8366 30064 8372
rect 30024 8090 30052 8366
rect 30012 8084 30064 8090
rect 30012 8026 30064 8032
rect 29920 8016 29972 8022
rect 29920 7958 29972 7964
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29104 7342 29132 7482
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28184 6458 28212 6734
rect 28644 6458 28672 6802
rect 28920 6730 28948 7142
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 28908 6724 28960 6730
rect 28908 6666 28960 6672
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28632 6452 28684 6458
rect 28632 6394 28684 6400
rect 29012 6322 29040 6802
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 27988 5568 28040 5574
rect 27988 5510 28040 5516
rect 28000 5098 28028 5510
rect 29012 5234 29040 5782
rect 29288 5778 29316 6734
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29288 5370 29316 5714
rect 29276 5364 29328 5370
rect 29276 5306 29328 5312
rect 29564 5234 29592 7142
rect 29748 6866 29776 7278
rect 30116 6934 30144 10202
rect 30392 10130 30420 11290
rect 30840 11280 30892 11286
rect 30840 11222 30892 11228
rect 30852 11121 30880 11222
rect 31024 11144 31076 11150
rect 30838 11112 30894 11121
rect 31024 11086 31076 11092
rect 30838 11047 30894 11056
rect 31036 10810 31064 11086
rect 31128 10810 31156 11494
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 30668 10266 30696 10406
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30392 9178 30420 10066
rect 30668 9450 30696 10202
rect 31208 9920 31260 9926
rect 31208 9862 31260 9868
rect 31220 9722 31248 9862
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 30656 9444 30708 9450
rect 30656 9386 30708 9392
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30668 9110 30696 9386
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30840 8424 30892 8430
rect 30840 8366 30892 8372
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31404 8378 31432 11018
rect 31772 10674 31800 11494
rect 32140 11218 32168 11698
rect 32784 11558 32812 12786
rect 32772 11552 32824 11558
rect 32772 11494 32824 11500
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 32140 10742 32168 11154
rect 32128 10736 32180 10742
rect 32128 10678 32180 10684
rect 32402 10704 32458 10713
rect 31760 10668 31812 10674
rect 32402 10639 32458 10648
rect 31760 10610 31812 10616
rect 32416 10606 32444 10639
rect 32404 10600 32456 10606
rect 32404 10542 32456 10548
rect 31668 10532 31720 10538
rect 31668 10474 31720 10480
rect 32496 10532 32548 10538
rect 32496 10474 32548 10480
rect 31680 10266 31708 10474
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31484 9512 31536 9518
rect 31484 9454 31536 9460
rect 32402 9480 32458 9489
rect 31496 8838 31524 9454
rect 31576 9444 31628 9450
rect 32402 9415 32458 9424
rect 31576 9386 31628 9392
rect 31484 8832 31536 8838
rect 31484 8774 31536 8780
rect 31496 8498 31524 8774
rect 31484 8492 31536 8498
rect 31484 8434 31536 8440
rect 30852 7954 30880 8366
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30484 7546 30512 7890
rect 30472 7540 30524 7546
rect 30472 7482 30524 7488
rect 30104 6928 30156 6934
rect 30104 6870 30156 6876
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 30024 6186 30052 6598
rect 29736 6180 29788 6186
rect 29736 6122 29788 6128
rect 30012 6180 30064 6186
rect 30012 6122 30064 6128
rect 29748 5642 29776 6122
rect 29736 5636 29788 5642
rect 29736 5578 29788 5584
rect 29748 5302 29776 5578
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 29736 5296 29788 5302
rect 29736 5238 29788 5244
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 27540 4826 27568 5034
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 28000 4758 28028 5034
rect 27988 4752 28040 4758
rect 27908 4712 27988 4740
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27632 4282 27660 4626
rect 27908 4282 27936 4712
rect 27988 4694 28040 4700
rect 28184 4622 28212 5170
rect 29460 5092 29512 5098
rect 29460 5034 29512 5040
rect 29472 4826 29500 5034
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29932 4758 29960 5510
rect 30024 5370 30052 6122
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 29920 4752 29972 4758
rect 29920 4694 29972 4700
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 28000 4282 28028 4558
rect 29012 4282 29040 4558
rect 27620 4276 27672 4282
rect 27620 4218 27672 4224
rect 27896 4276 27948 4282
rect 27896 4218 27948 4224
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 27632 4185 27660 4218
rect 27618 4176 27674 4185
rect 27618 4111 27674 4120
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27540 2553 27568 4014
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28000 3738 28028 4218
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 27988 3732 28040 3738
rect 27988 3674 28040 3680
rect 28092 3602 28120 4150
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 28814 3768 28870 3777
rect 28814 3703 28870 3712
rect 28828 3670 28856 3703
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28828 2650 28856 3606
rect 29288 3505 29316 4014
rect 29932 3738 29960 4694
rect 30116 4622 30144 6870
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30392 6118 30420 6802
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 30484 4146 30512 7482
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30564 6180 30616 6186
rect 30564 6122 30616 6128
rect 30576 5302 30604 6122
rect 30564 5296 30616 5302
rect 30564 5238 30616 5244
rect 30576 4758 30604 5238
rect 30564 4752 30616 4758
rect 30564 4694 30616 4700
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30472 3936 30524 3942
rect 30668 3924 30696 7346
rect 30852 6798 30880 7890
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 31128 7002 31156 7278
rect 31116 6996 31168 7002
rect 31116 6938 31168 6944
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30852 6458 30880 6734
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 31208 6112 31260 6118
rect 31208 6054 31260 6060
rect 31220 5166 31248 6054
rect 31208 5160 31260 5166
rect 31208 5102 31260 5108
rect 31220 4826 31248 5102
rect 31312 5030 31340 8366
rect 31404 8350 31524 8378
rect 31588 8362 31616 9386
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32324 8634 32352 9318
rect 32416 8820 32444 9415
rect 32508 9382 32536 10474
rect 32496 9376 32548 9382
rect 32496 9318 32548 9324
rect 32508 9042 32536 9318
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32496 8832 32548 8838
rect 32416 8792 32496 8820
rect 32496 8774 32548 8780
rect 32508 8634 32536 8774
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32784 8401 32812 11494
rect 33336 11354 33364 15558
rect 33690 15520 33746 15558
rect 35912 15558 36230 15586
rect 35714 14784 35770 14793
rect 35714 14719 35770 14728
rect 35622 13696 35678 13705
rect 35622 13631 35678 13640
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35636 12986 35664 13631
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 33876 12776 33928 12782
rect 33876 12718 33928 12724
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 33612 11898 33640 12242
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 33612 11558 33640 11834
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 32864 10804 32916 10810
rect 32864 10746 32916 10752
rect 32876 9586 32904 10746
rect 32968 10062 32996 10950
rect 33888 10826 33916 12718
rect 35348 12300 35400 12306
rect 35348 12242 35400 12248
rect 34704 12096 34756 12102
rect 34704 12038 34756 12044
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 33968 11688 34020 11694
rect 33968 11630 34020 11636
rect 33980 10985 34008 11630
rect 34152 11552 34204 11558
rect 34152 11494 34204 11500
rect 34164 11286 34192 11494
rect 34152 11280 34204 11286
rect 34152 11222 34204 11228
rect 34612 11280 34664 11286
rect 34612 11222 34664 11228
rect 33966 10976 34022 10985
rect 33966 10911 34022 10920
rect 33796 10798 33916 10826
rect 33980 10810 34008 10911
rect 33968 10804 34020 10810
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 33416 10532 33468 10538
rect 33416 10474 33468 10480
rect 33140 10464 33192 10470
rect 33192 10424 33272 10452
rect 33140 10406 33192 10412
rect 32956 10056 33008 10062
rect 32956 9998 33008 10004
rect 32864 9580 32916 9586
rect 32864 9522 32916 9528
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 32956 8492 33008 8498
rect 32956 8434 33008 8440
rect 32770 8392 32826 8401
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31300 5024 31352 5030
rect 31300 4966 31352 4972
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31404 4146 31432 6598
rect 31496 6254 31524 8350
rect 31576 8356 31628 8362
rect 32770 8327 32826 8336
rect 31576 8298 31628 8304
rect 32968 8090 32996 8434
rect 33060 8294 33088 8910
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33048 8288 33100 8294
rect 33048 8230 33100 8236
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 33060 8022 33088 8230
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 32864 7336 32916 7342
rect 32864 7278 32916 7284
rect 32404 6860 32456 6866
rect 32404 6802 32456 6808
rect 32588 6860 32640 6866
rect 32588 6802 32640 6808
rect 32416 6390 32444 6802
rect 32600 6458 32628 6802
rect 32588 6452 32640 6458
rect 32588 6394 32640 6400
rect 32404 6384 32456 6390
rect 32404 6326 32456 6332
rect 31484 6248 31536 6254
rect 31484 6190 31536 6196
rect 31496 5574 31524 6190
rect 32128 6180 32180 6186
rect 32128 6122 32180 6128
rect 32140 5778 32168 6122
rect 32496 5840 32548 5846
rect 32496 5782 32548 5788
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 31484 5568 31536 5574
rect 31484 5510 31536 5516
rect 32140 4826 32168 5714
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 32128 4820 32180 4826
rect 32128 4762 32180 4768
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 30932 4004 30984 4010
rect 30932 3946 30984 3952
rect 30524 3896 30696 3924
rect 30472 3878 30524 3884
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 30944 3602 30972 3946
rect 32048 3738 32076 4558
rect 32232 4078 32260 5510
rect 32508 5098 32536 5782
rect 32600 5166 32628 6394
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 32600 4690 32628 5102
rect 32876 4758 32904 7278
rect 33060 6662 33088 7822
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33152 5710 33180 8774
rect 33244 6322 33272 10424
rect 33428 10198 33456 10474
rect 33520 10470 33548 10678
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33416 10192 33468 10198
rect 33416 10134 33468 10140
rect 33416 8832 33468 8838
rect 33416 8774 33468 8780
rect 33428 8362 33456 8774
rect 33324 8356 33376 8362
rect 33324 8298 33376 8304
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33336 8090 33364 8298
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33336 7206 33364 8026
rect 33428 7478 33456 8298
rect 33416 7472 33468 7478
rect 33416 7414 33468 7420
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 33428 7002 33456 7414
rect 33416 6996 33468 7002
rect 33416 6938 33468 6944
rect 33232 6316 33284 6322
rect 33232 6258 33284 6264
rect 33244 5914 33272 6258
rect 33428 6186 33456 6938
rect 33416 6180 33468 6186
rect 33416 6122 33468 6128
rect 33232 5908 33284 5914
rect 33232 5850 33284 5856
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33324 5568 33376 5574
rect 33324 5510 33376 5516
rect 33336 5098 33364 5510
rect 33232 5092 33284 5098
rect 33232 5034 33284 5040
rect 33324 5092 33376 5098
rect 33324 5034 33376 5040
rect 32864 4752 32916 4758
rect 32864 4694 32916 4700
rect 33244 4690 33272 5034
rect 33336 4826 33364 5034
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 32588 4684 32640 4690
rect 32588 4626 32640 4632
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 32600 4078 32628 4626
rect 32220 4072 32272 4078
rect 32220 4014 32272 4020
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32508 3738 32536 4014
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 29274 3496 29330 3505
rect 29274 3431 29330 3440
rect 30760 3194 30788 3538
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30944 3126 30972 3538
rect 30932 3120 30984 3126
rect 30932 3062 30984 3068
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 27526 2544 27582 2553
rect 27526 2479 27582 2488
rect 33520 2417 33548 10406
rect 33692 9444 33744 9450
rect 33692 9386 33744 9392
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 33612 8634 33640 8774
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 33612 5574 33640 6734
rect 33704 6322 33732 9386
rect 33796 7410 33824 10798
rect 33968 10746 34020 10752
rect 34164 10266 34192 11222
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34624 10538 34652 11222
rect 34612 10532 34664 10538
rect 34612 10474 34664 10480
rect 34716 10266 34744 12038
rect 35164 11688 35216 11694
rect 35164 11630 35216 11636
rect 34980 11076 35032 11082
rect 34980 11018 35032 11024
rect 34992 10674 35020 11018
rect 35072 11008 35124 11014
rect 35072 10950 35124 10956
rect 34980 10668 35032 10674
rect 34980 10610 35032 10616
rect 34152 10260 34204 10266
rect 34152 10202 34204 10208
rect 34704 10260 34756 10266
rect 34704 10202 34756 10208
rect 34612 10192 34664 10198
rect 34612 10134 34664 10140
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34624 9722 34652 10134
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 34716 9432 34744 10202
rect 34992 10062 35020 10610
rect 35084 10538 35112 10950
rect 35176 10742 35204 11630
rect 35360 11558 35388 12242
rect 35728 11898 35756 14719
rect 35912 12918 35940 15558
rect 36174 15520 36230 15558
rect 38658 15586 38714 16000
rect 38658 15558 38792 15586
rect 38658 15520 38714 15558
rect 35900 12912 35952 12918
rect 35900 12854 35952 12860
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 37094 12064 37150 12073
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 35164 10736 35216 10742
rect 35164 10678 35216 10684
rect 35072 10532 35124 10538
rect 35072 10474 35124 10480
rect 34888 10056 34940 10062
rect 34888 9998 34940 10004
rect 34980 10056 35032 10062
rect 34980 9998 35032 10004
rect 34796 9444 34848 9450
rect 34716 9404 34796 9432
rect 34796 9386 34848 9392
rect 34428 9376 34480 9382
rect 34428 9318 34480 9324
rect 34520 9376 34572 9382
rect 34520 9318 34572 9324
rect 34440 9042 34468 9318
rect 34532 9178 34560 9318
rect 34520 9172 34572 9178
rect 34520 9114 34572 9120
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 34428 9036 34480 9042
rect 34428 8978 34480 8984
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33888 6934 33916 8910
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34624 8566 34652 9046
rect 34900 8566 34928 9998
rect 34992 9586 35020 9998
rect 35084 9654 35112 10474
rect 35176 10198 35204 10678
rect 35256 10464 35308 10470
rect 35256 10406 35308 10412
rect 35164 10192 35216 10198
rect 35164 10134 35216 10140
rect 35072 9648 35124 9654
rect 35072 9590 35124 9596
rect 34980 9580 35032 9586
rect 34980 9522 35032 9528
rect 34980 9172 35032 9178
rect 34980 9114 35032 9120
rect 34612 8560 34664 8566
rect 34612 8502 34664 8508
rect 34888 8560 34940 8566
rect 34888 8502 34940 8508
rect 34992 8498 35020 9114
rect 35268 8634 35296 10406
rect 35360 8838 35388 11494
rect 35992 11212 36044 11218
rect 35992 11154 36044 11160
rect 35808 11008 35860 11014
rect 35808 10950 35860 10956
rect 35820 9178 35848 10950
rect 36004 10538 36032 11154
rect 36450 10568 36506 10577
rect 35992 10532 36044 10538
rect 35992 10474 36044 10480
rect 36084 10532 36136 10538
rect 36450 10503 36506 10512
rect 36084 10474 36136 10480
rect 36004 10441 36032 10474
rect 35990 10432 36046 10441
rect 35990 10367 36046 10376
rect 36004 10033 36032 10367
rect 36096 10198 36124 10474
rect 36084 10192 36136 10198
rect 36084 10134 36136 10140
rect 36176 10192 36228 10198
rect 36176 10134 36228 10140
rect 35990 10024 36046 10033
rect 35990 9959 36046 9968
rect 36188 9722 36216 10134
rect 36176 9716 36228 9722
rect 36176 9658 36228 9664
rect 36188 9178 36216 9658
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 36176 9172 36228 9178
rect 36176 9114 36228 9120
rect 35900 9104 35952 9110
rect 35900 9046 35952 9052
rect 35348 8832 35400 8838
rect 35348 8774 35400 8780
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 33968 8356 34020 8362
rect 33968 8298 34020 8304
rect 33980 7886 34008 8298
rect 35072 8016 35124 8022
rect 35072 7958 35124 7964
rect 33968 7880 34020 7886
rect 33968 7822 34020 7828
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 7546 34192 7686
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 34072 7002 34100 7142
rect 34060 6996 34112 7002
rect 34060 6938 34112 6944
rect 33876 6928 33928 6934
rect 33876 6870 33928 6876
rect 34072 6458 34100 6938
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34060 6452 34112 6458
rect 34060 6394 34112 6400
rect 33692 6316 33744 6322
rect 33692 6258 33744 6264
rect 34624 5846 34652 7142
rect 35084 7002 35112 7958
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35268 7410 35296 7686
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 35072 6996 35124 7002
rect 35072 6938 35124 6944
rect 34704 6860 34756 6866
rect 34704 6802 34756 6808
rect 34716 6322 34744 6802
rect 35072 6724 35124 6730
rect 35072 6666 35124 6672
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33600 5568 33652 5574
rect 33600 5510 33652 5516
rect 33612 4146 33640 5510
rect 34164 4826 34192 5646
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34624 5370 34652 5782
rect 34716 5710 34744 6258
rect 35084 6186 35112 6666
rect 35268 6186 35296 7346
rect 34796 6180 34848 6186
rect 34796 6122 34848 6128
rect 35072 6180 35124 6186
rect 35072 6122 35124 6128
rect 35256 6180 35308 6186
rect 35256 6122 35308 6128
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34808 5234 34836 6122
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 34624 4690 34652 5170
rect 34612 4684 34664 4690
rect 34612 4626 34664 4632
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34624 4282 34652 4626
rect 34612 4276 34664 4282
rect 34612 4218 34664 4224
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 35360 3233 35388 8774
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35728 7886 35756 8434
rect 35912 8294 35940 9046
rect 36188 8362 36216 9114
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8634 36308 8910
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36176 8356 36228 8362
rect 36176 8298 36228 8304
rect 35900 8288 35952 8294
rect 35900 8230 35952 8236
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35532 7812 35584 7818
rect 35532 7754 35584 7760
rect 35544 7392 35572 7754
rect 35624 7404 35676 7410
rect 35544 7364 35624 7392
rect 35440 6792 35492 6798
rect 35440 6734 35492 6740
rect 35452 6322 35480 6734
rect 35544 6390 35572 7364
rect 35624 7346 35676 7352
rect 35728 7274 35756 7822
rect 35716 7268 35768 7274
rect 35716 7210 35768 7216
rect 35912 6934 35940 8230
rect 36268 7948 36320 7954
rect 36268 7890 36320 7896
rect 36280 7206 36308 7890
rect 36360 7268 36412 7274
rect 36360 7210 36412 7216
rect 36268 7200 36320 7206
rect 36268 7142 36320 7148
rect 35900 6928 35952 6934
rect 35900 6870 35952 6876
rect 35912 6458 35940 6870
rect 36280 6769 36308 7142
rect 36372 6866 36400 7210
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 36266 6760 36322 6769
rect 36266 6695 36322 6704
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35452 3670 35480 6258
rect 35544 5778 35572 6326
rect 36360 6248 36412 6254
rect 36464 6225 36492 10503
rect 36556 9586 36584 12038
rect 37094 11999 37150 12008
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36636 9444 36688 9450
rect 36636 9386 36688 9392
rect 36648 9178 36676 9386
rect 36636 9172 36688 9178
rect 36636 9114 36688 9120
rect 36636 9036 36688 9042
rect 36636 8978 36688 8984
rect 36648 8362 36676 8978
rect 36544 8356 36596 8362
rect 36544 8298 36596 8304
rect 36636 8356 36688 8362
rect 36636 8298 36688 8304
rect 36360 6190 36412 6196
rect 36450 6216 36506 6225
rect 35532 5772 35584 5778
rect 35532 5714 35584 5720
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35440 3664 35492 3670
rect 35440 3606 35492 3612
rect 35346 3224 35402 3233
rect 35346 3159 35402 3168
rect 33506 2408 33562 2417
rect 29644 2372 29696 2378
rect 33506 2343 33562 2352
rect 29644 2314 29696 2320
rect 27066 54 27384 82
rect 29656 82 29684 2314
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 32494 1864 32550 1873
rect 32494 1799 32550 1808
rect 29918 82 29974 480
rect 29656 54 29974 82
rect 32508 82 32536 1799
rect 32770 82 32826 480
rect 32508 54 32826 82
rect 27066 0 27122 54
rect 29918 0 29974 54
rect 32770 0 32826 54
rect 35622 82 35678 480
rect 35912 82 35940 5510
rect 36372 4185 36400 6190
rect 36450 6151 36506 6160
rect 36464 5302 36492 6151
rect 36556 5370 36584 8298
rect 36636 7472 36688 7478
rect 36636 7414 36688 7420
rect 36648 7274 36676 7414
rect 36636 7268 36688 7274
rect 36636 7210 36688 7216
rect 36634 6760 36690 6769
rect 36634 6695 36690 6704
rect 36648 6458 36676 6695
rect 37108 6458 37136 11999
rect 38764 11121 38792 15558
rect 39578 11248 39634 11257
rect 39578 11183 39634 11192
rect 38750 11112 38806 11121
rect 38750 11047 38806 11056
rect 39592 10810 39620 11183
rect 39580 10804 39632 10810
rect 39580 10746 39632 10752
rect 37924 10668 37976 10674
rect 37924 10610 37976 10616
rect 37936 10577 37964 10610
rect 37922 10568 37978 10577
rect 37922 10503 37978 10512
rect 37188 9444 37240 9450
rect 37188 9386 37240 9392
rect 37200 8566 37228 9386
rect 37188 8560 37240 8566
rect 37188 8502 37240 8508
rect 38014 8392 38070 8401
rect 38014 8327 38070 8336
rect 37738 8256 37794 8265
rect 37738 8191 37794 8200
rect 37752 8090 37780 8191
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 36636 6452 36688 6458
rect 36636 6394 36688 6400
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 37108 6254 37136 6394
rect 38028 6254 38056 8327
rect 37096 6248 37148 6254
rect 37096 6190 37148 6196
rect 38016 6248 38068 6254
rect 38016 6190 38068 6196
rect 36728 5772 36780 5778
rect 36728 5714 36780 5720
rect 36740 5370 36768 5714
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36728 5364 36780 5370
rect 36728 5306 36780 5312
rect 36452 5296 36504 5302
rect 36452 5238 36504 5244
rect 38568 4480 38620 4486
rect 38568 4422 38620 4428
rect 36358 4176 36414 4185
rect 36358 4111 36414 4120
rect 35622 54 35940 82
rect 38474 82 38530 480
rect 38580 82 38608 4422
rect 38474 54 38608 82
rect 35622 0 35678 54
rect 38474 0 38530 54
<< via2 >>
rect 110 14320 166 14376
rect 18 13096 74 13152
rect 110 9696 166 9752
rect 110 8608 166 8664
rect 110 8336 166 8392
rect 1674 10648 1730 10704
rect 1582 10240 1638 10296
rect 1582 6840 1638 6896
rect 2042 6196 2044 6216
rect 2044 6196 2096 6216
rect 2096 6196 2098 6216
rect 2042 6160 2098 6196
rect 1582 4664 1638 4720
rect 2318 7812 2374 7848
rect 2318 7792 2320 7812
rect 2320 7792 2372 7812
rect 2372 7792 2374 7812
rect 2410 5616 2466 5672
rect 2410 3712 2466 3768
rect 1858 1128 1914 1184
rect 3146 11056 3202 11112
rect 2594 5208 2650 5264
rect 2778 5752 2834 5808
rect 2778 5072 2834 5128
rect 3054 6160 3110 6216
rect 5170 7928 5226 7984
rect 3974 5072 4030 5128
rect 7194 14864 7250 14920
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 7470 11600 7526 11656
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 8022 10784 8078 10840
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7010 8336 7066 8392
rect 5538 3304 5594 3360
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7654 8336 7710 8392
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 8298 7520 8354 7576
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7010 2624 7066 2680
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 8114 3440 8170 3496
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 9218 7248 9274 7304
rect 8666 3168 8722 3224
rect 11150 11056 11206 11112
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 8298 2896 8354 2952
rect 7470 2216 7526 2272
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 10966 7792 11022 7848
rect 11242 6160 11298 6216
rect 12254 7928 12310 7984
rect 11702 3712 11758 3768
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 13358 10784 13414 10840
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 13634 10784 13690 10840
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14094 5208 14150 5264
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14922 8336 14978 8392
rect 14922 5072 14978 5128
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 14094 2624 14150 2680
rect 15474 5616 15530 5672
rect 15014 3576 15070 3632
rect 11886 40 11942 96
rect 16670 7384 16726 7440
rect 19798 11328 19854 11384
rect 17774 7520 17830 7576
rect 17958 7384 18014 7440
rect 17314 2896 17370 2952
rect 15382 1808 15438 1864
rect 18786 4684 18842 4720
rect 18786 4664 18788 4684
rect 18788 4664 18840 4684
rect 18840 4664 18842 4684
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20810 10784 20866 10840
rect 20810 9968 20866 10024
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 18602 2488 18658 2544
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 22282 10648 22338 10704
rect 22282 9424 22338 9480
rect 23110 10920 23166 10976
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20718 3168 20774 3224
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 24122 11600 24178 11656
rect 24214 11328 24270 11384
rect 23938 10648 23994 10704
rect 23662 9696 23718 9752
rect 23478 7928 23534 7984
rect 23570 7384 23626 7440
rect 23110 6704 23166 6760
rect 26054 11736 26110 11792
rect 25318 10512 25374 10568
rect 26238 11328 26294 11384
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 26698 11736 26754 11792
rect 26606 11328 26662 11384
rect 26882 9696 26938 9752
rect 25134 4664 25190 4720
rect 27434 10512 27490 10568
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 28078 7248 28134 7304
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 30838 11056 30894 11112
rect 32402 10648 32458 10704
rect 32402 9424 32458 9480
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 27618 4120 27674 4176
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 28814 3712 28870 3768
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 35714 14728 35770 14784
rect 35622 13640 35678 13696
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 33966 10920 34022 10976
rect 32770 8336 32826 8392
rect 29274 3440 29330 3496
rect 27526 2488 27582 2544
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 36450 10512 36506 10568
rect 35990 10376 36046 10432
rect 35990 9968 36046 10024
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 36266 6704 36322 6760
rect 37094 12008 37150 12064
rect 35346 3168 35402 3224
rect 33506 2352 33562 2408
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 32494 1808 32550 1864
rect 36450 6160 36506 6216
rect 36634 6704 36690 6760
rect 39578 11192 39634 11248
rect 38750 11056 38806 11112
rect 37922 10512 37978 10568
rect 38014 8336 38070 8392
rect 37738 8200 37794 8256
rect 36358 4120 36414 4176
<< metal3 >>
rect 0 15376 480 15496
rect 62 14922 122 15376
rect 39520 15240 40000 15360
rect 7189 14922 7255 14925
rect 62 14920 7255 14922
rect 62 14864 7194 14920
rect 7250 14864 7255 14920
rect 62 14862 7255 14864
rect 7189 14859 7255 14862
rect 35709 14786 35775 14789
rect 39622 14786 39682 15240
rect 35709 14784 39682 14786
rect 35709 14728 35714 14784
rect 35770 14728 39682 14784
rect 35709 14726 39682 14728
rect 35709 14723 35775 14726
rect 0 14376 480 14408
rect 0 14320 110 14376
rect 166 14320 480 14376
rect 0 14288 480 14320
rect 39520 13880 40000 14000
rect 35617 13698 35683 13701
rect 39622 13698 39682 13880
rect 35617 13696 39682 13698
rect 35617 13640 35622 13696
rect 35678 13640 39682 13696
rect 35617 13638 39682 13640
rect 35617 13635 35683 13638
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 0 13152 480 13184
rect 0 13096 18 13152
rect 74 13096 480 13152
rect 0 13064 480 13096
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 39520 12520 40000 12640
rect 27610 12479 27930 12480
rect 0 11976 480 12096
rect 37089 12066 37155 12069
rect 39622 12066 39682 12520
rect 37089 12064 39682 12066
rect 37089 12008 37094 12064
rect 37150 12008 39682 12064
rect 37089 12006 39682 12008
rect 37089 12003 37155 12006
rect 7610 12000 7930 12001
rect 62 11522 122 11976
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 26049 11794 26115 11797
rect 26693 11794 26759 11797
rect 26049 11792 26759 11794
rect 26049 11736 26054 11792
rect 26110 11736 26698 11792
rect 26754 11736 26759 11792
rect 26049 11734 26759 11736
rect 26049 11731 26115 11734
rect 26693 11731 26759 11734
rect 7465 11658 7531 11661
rect 24117 11658 24183 11661
rect 7465 11656 24183 11658
rect 7465 11600 7470 11656
rect 7526 11600 24122 11656
rect 24178 11600 24183 11656
rect 7465 11598 24183 11600
rect 7465 11595 7531 11598
rect 24117 11595 24183 11598
rect 9622 11522 9628 11524
rect 62 11462 9628 11522
rect 9622 11460 9628 11462
rect 9692 11460 9698 11524
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 19793 11386 19859 11389
rect 24209 11386 24275 11389
rect 26233 11386 26299 11389
rect 26601 11386 26667 11389
rect 19793 11384 26667 11386
rect 19793 11328 19798 11384
rect 19854 11328 24214 11384
rect 24270 11328 26238 11384
rect 26294 11328 26606 11384
rect 26662 11328 26667 11384
rect 19793 11326 26667 11328
rect 19793 11323 19859 11326
rect 24209 11323 24275 11326
rect 26233 11323 26299 11326
rect 26601 11323 26667 11326
rect 39520 11250 40000 11280
rect 39492 11248 40000 11250
rect 39492 11192 39578 11248
rect 39634 11192 40000 11248
rect 39492 11190 40000 11192
rect 39520 11160 40000 11190
rect 3141 11114 3207 11117
rect 11145 11114 11211 11117
rect 3141 11112 11211 11114
rect 3141 11056 3146 11112
rect 3202 11056 11150 11112
rect 11206 11056 11211 11112
rect 3141 11054 11211 11056
rect 3141 11051 3207 11054
rect 11145 11051 11211 11054
rect 30833 11114 30899 11117
rect 38745 11114 38811 11117
rect 30833 11112 38811 11114
rect 30833 11056 30838 11112
rect 30894 11056 38750 11112
rect 38806 11056 38811 11112
rect 30833 11054 38811 11056
rect 30833 11051 30899 11054
rect 38745 11051 38811 11054
rect 23105 10978 23171 10981
rect 33961 10978 34027 10981
rect 23105 10976 34027 10978
rect 23105 10920 23110 10976
rect 23166 10920 33966 10976
rect 34022 10920 34027 10976
rect 23105 10918 34027 10920
rect 23105 10915 23171 10918
rect 33961 10915 34027 10918
rect 7610 10912 7930 10913
rect 0 10752 480 10872
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 8017 10842 8083 10845
rect 13353 10842 13419 10845
rect 8017 10840 13419 10842
rect 8017 10784 8022 10840
rect 8078 10784 13358 10840
rect 13414 10784 13419 10840
rect 8017 10782 13419 10784
rect 8017 10779 8083 10782
rect 13353 10779 13419 10782
rect 13629 10842 13695 10845
rect 20805 10842 20871 10845
rect 13629 10840 20871 10842
rect 13629 10784 13634 10840
rect 13690 10784 20810 10840
rect 20866 10784 20871 10840
rect 13629 10782 20871 10784
rect 13629 10779 13695 10782
rect 20805 10779 20871 10782
rect 62 10298 122 10752
rect 1669 10706 1735 10709
rect 22277 10706 22343 10709
rect 1669 10704 22343 10706
rect 1669 10648 1674 10704
rect 1730 10648 22282 10704
rect 22338 10648 22343 10704
rect 1669 10646 22343 10648
rect 1669 10643 1735 10646
rect 22277 10643 22343 10646
rect 23933 10706 23999 10709
rect 32397 10706 32463 10709
rect 23933 10704 32463 10706
rect 23933 10648 23938 10704
rect 23994 10648 32402 10704
rect 32458 10648 32463 10704
rect 23933 10646 32463 10648
rect 23933 10643 23999 10646
rect 32397 10643 32463 10646
rect 23422 10508 23428 10572
rect 23492 10570 23498 10572
rect 25313 10570 25379 10573
rect 23492 10568 25379 10570
rect 23492 10512 25318 10568
rect 25374 10512 25379 10568
rect 23492 10510 25379 10512
rect 23492 10508 23498 10510
rect 25313 10507 25379 10510
rect 27429 10570 27495 10573
rect 36445 10570 36511 10573
rect 37917 10570 37983 10573
rect 27429 10568 37983 10570
rect 27429 10512 27434 10568
rect 27490 10512 36450 10568
rect 36506 10512 37922 10568
rect 37978 10512 37983 10568
rect 27429 10510 37983 10512
rect 27429 10507 27495 10510
rect 36445 10507 36511 10510
rect 37917 10507 37983 10510
rect 35985 10434 36051 10437
rect 35985 10432 39682 10434
rect 35985 10376 35990 10432
rect 36046 10376 39682 10432
rect 35985 10374 39682 10376
rect 35985 10371 36051 10374
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 1577 10298 1643 10301
rect 62 10296 1643 10298
rect 62 10240 1582 10296
rect 1638 10240 1643 10296
rect 62 10238 1643 10240
rect 1577 10235 1643 10238
rect 20805 10026 20871 10029
rect 35985 10026 36051 10029
rect 20805 10024 36051 10026
rect 20805 9968 20810 10024
rect 20866 9968 35990 10024
rect 36046 9968 36051 10024
rect 20805 9966 36051 9968
rect 20805 9963 20871 9966
rect 35985 9963 36051 9966
rect 39622 9920 39682 10374
rect 7610 9824 7930 9825
rect 0 9752 480 9784
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 39520 9800 40000 9920
rect 34277 9759 34597 9760
rect 0 9696 110 9752
rect 166 9696 480 9752
rect 0 9664 480 9696
rect 23657 9754 23723 9757
rect 26877 9754 26943 9757
rect 23657 9752 26943 9754
rect 23657 9696 23662 9752
rect 23718 9696 26882 9752
rect 26938 9696 26943 9752
rect 23657 9694 26943 9696
rect 23657 9691 23723 9694
rect 26877 9691 26943 9694
rect 22277 9482 22343 9485
rect 32397 9482 32463 9485
rect 22277 9480 32463 9482
rect 22277 9424 22282 9480
rect 22338 9424 32402 9480
rect 32458 9424 32463 9480
rect 22277 9422 32463 9424
rect 22277 9419 22343 9422
rect 32397 9419 32463 9422
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 7610 8736 7930 8737
rect 0 8664 480 8696
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8608 110 8664
rect 166 8608 480 8664
rect 0 8576 480 8608
rect 39520 8576 40000 8696
rect 105 8394 171 8397
rect 7005 8394 7071 8397
rect 105 8392 7071 8394
rect 105 8336 110 8392
rect 166 8336 7010 8392
rect 7066 8336 7071 8392
rect 105 8334 7071 8336
rect 105 8331 171 8334
rect 7005 8331 7071 8334
rect 7649 8394 7715 8397
rect 14917 8394 14983 8397
rect 7649 8392 14983 8394
rect 7649 8336 7654 8392
rect 7710 8336 14922 8392
rect 14978 8336 14983 8392
rect 7649 8334 14983 8336
rect 7649 8331 7715 8334
rect 14917 8331 14983 8334
rect 32765 8394 32831 8397
rect 38009 8394 38075 8397
rect 32765 8392 38075 8394
rect 32765 8336 32770 8392
rect 32826 8336 38014 8392
rect 38070 8336 38075 8392
rect 32765 8334 38075 8336
rect 32765 8331 32831 8334
rect 38009 8331 38075 8334
rect 37733 8258 37799 8261
rect 39622 8258 39682 8576
rect 37733 8256 39682 8258
rect 37733 8200 37738 8256
rect 37794 8200 39682 8256
rect 37733 8198 39682 8200
rect 37733 8195 37799 8198
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 5165 7986 5231 7989
rect 12249 7986 12315 7989
rect 23473 7986 23539 7989
rect 5165 7984 23539 7986
rect 5165 7928 5170 7984
rect 5226 7928 12254 7984
rect 12310 7928 23478 7984
rect 23534 7928 23539 7984
rect 5165 7926 23539 7928
rect 5165 7923 5231 7926
rect 12249 7923 12315 7926
rect 23473 7923 23539 7926
rect 2313 7850 2379 7853
rect 10961 7850 11027 7853
rect 2313 7848 11027 7850
rect 2313 7792 2318 7848
rect 2374 7792 10966 7848
rect 11022 7792 11027 7848
rect 2313 7790 11027 7792
rect 2313 7787 2379 7790
rect 10961 7787 11027 7790
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 8293 7578 8359 7581
rect 17769 7578 17835 7581
rect 8293 7576 17835 7578
rect 8293 7520 8298 7576
rect 8354 7520 17774 7576
rect 17830 7520 17835 7576
rect 8293 7518 17835 7520
rect 8293 7515 8359 7518
rect 17769 7515 17835 7518
rect 0 7352 480 7472
rect 16665 7442 16731 7445
rect 17953 7442 18019 7445
rect 23565 7442 23631 7445
rect 16665 7440 23631 7442
rect 16665 7384 16670 7440
rect 16726 7384 17958 7440
rect 18014 7384 23570 7440
rect 23626 7384 23631 7440
rect 16665 7382 23631 7384
rect 16665 7379 16731 7382
rect 17953 7379 18019 7382
rect 23565 7379 23631 7382
rect 62 6898 122 7352
rect 9213 7306 9279 7309
rect 28073 7306 28139 7309
rect 9213 7304 28139 7306
rect 9213 7248 9218 7304
rect 9274 7248 28078 7304
rect 28134 7248 28139 7304
rect 9213 7246 28139 7248
rect 9213 7243 9279 7246
rect 28073 7243 28139 7246
rect 39520 7216 40000 7336
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 1577 6898 1643 6901
rect 62 6896 1643 6898
rect 62 6840 1582 6896
rect 1638 6840 1643 6896
rect 62 6838 1643 6840
rect 1577 6835 1643 6838
rect 23105 6762 23171 6765
rect 36261 6762 36327 6765
rect 23105 6760 36327 6762
rect 23105 6704 23110 6760
rect 23166 6704 36266 6760
rect 36322 6704 36327 6760
rect 23105 6702 36327 6704
rect 23105 6699 23171 6702
rect 36261 6699 36327 6702
rect 36629 6762 36695 6765
rect 39622 6762 39682 7216
rect 36629 6760 39682 6762
rect 36629 6704 36634 6760
rect 36690 6704 39682 6760
rect 36629 6702 39682 6704
rect 36629 6699 36695 6702
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 0 6264 480 6384
rect 62 5810 122 6264
rect 2037 6218 2103 6221
rect 3049 6218 3115 6221
rect 11237 6218 11303 6221
rect 2037 6216 11303 6218
rect 2037 6160 2042 6216
rect 2098 6160 3054 6216
rect 3110 6160 11242 6216
rect 11298 6160 11303 6216
rect 2037 6158 11303 6160
rect 2037 6155 2103 6158
rect 3049 6155 3115 6158
rect 11237 6155 11303 6158
rect 36445 6218 36511 6221
rect 39614 6218 39620 6220
rect 36445 6216 39620 6218
rect 36445 6160 36450 6216
rect 36506 6160 39620 6216
rect 36445 6158 39620 6160
rect 36445 6155 36511 6158
rect 39614 6156 39620 6158
rect 39684 6156 39690 6220
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 39520 5948 40000 5976
rect 39520 5946 39620 5948
rect 39492 5886 39620 5946
rect 39520 5884 39620 5886
rect 39684 5884 40000 5948
rect 39520 5856 40000 5884
rect 2773 5810 2839 5813
rect 62 5808 2839 5810
rect 62 5752 2778 5808
rect 2834 5752 2839 5808
rect 62 5750 2839 5752
rect 2773 5747 2839 5750
rect 2405 5674 2471 5677
rect 15469 5674 15535 5677
rect 2405 5672 15535 5674
rect 2405 5616 2410 5672
rect 2466 5616 15474 5672
rect 15530 5616 15535 5672
rect 2405 5614 15535 5616
rect 2405 5611 2471 5614
rect 15469 5611 15535 5614
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 2589 5266 2655 5269
rect 14089 5266 14155 5269
rect 2589 5264 14155 5266
rect 2589 5208 2594 5264
rect 2650 5208 14094 5264
rect 14150 5208 14155 5264
rect 2589 5206 14155 5208
rect 2589 5203 2655 5206
rect 14089 5203 14155 5206
rect 0 5040 480 5160
rect 2773 5130 2839 5133
rect 3969 5130 4035 5133
rect 14917 5130 14983 5133
rect 2773 5128 14983 5130
rect 2773 5072 2778 5128
rect 2834 5072 3974 5128
rect 4030 5072 14922 5128
rect 14978 5072 14983 5128
rect 2773 5070 14983 5072
rect 2773 5067 2839 5070
rect 3969 5067 4035 5070
rect 14917 5067 14983 5070
rect 62 4722 122 5040
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 1577 4722 1643 4725
rect 62 4720 1643 4722
rect 62 4664 1582 4720
rect 1638 4664 1643 4720
rect 62 4662 1643 4664
rect 1577 4659 1643 4662
rect 18781 4722 18847 4725
rect 25129 4722 25195 4725
rect 18781 4720 25195 4722
rect 18781 4664 18786 4720
rect 18842 4664 25134 4720
rect 25190 4664 25195 4720
rect 18781 4662 25195 4664
rect 18781 4659 18847 4662
rect 25129 4659 25195 4662
rect 39520 4496 40000 4616
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 27613 4178 27679 4181
rect 36353 4178 36419 4181
rect 27613 4176 36419 4178
rect 27613 4120 27618 4176
rect 27674 4120 36358 4176
rect 36414 4120 36419 4176
rect 27613 4118 36419 4120
rect 27613 4115 27679 4118
rect 36353 4115 36419 4118
rect 0 3952 480 4072
rect 62 3634 122 3952
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 2405 3770 2471 3773
rect 11697 3770 11763 3773
rect 2405 3768 11763 3770
rect 2405 3712 2410 3768
rect 2466 3712 11702 3768
rect 11758 3712 11763 3768
rect 2405 3710 11763 3712
rect 2405 3707 2471 3710
rect 11697 3707 11763 3710
rect 28809 3770 28875 3773
rect 39622 3770 39682 4496
rect 28809 3768 39682 3770
rect 28809 3712 28814 3768
rect 28870 3712 39682 3768
rect 28809 3710 39682 3712
rect 28809 3707 28875 3710
rect 15009 3634 15075 3637
rect 62 3632 15075 3634
rect 62 3576 15014 3632
rect 15070 3576 15075 3632
rect 62 3574 15075 3576
rect 15009 3571 15075 3574
rect 8109 3498 8175 3501
rect 29269 3498 29335 3501
rect 8109 3496 29335 3498
rect 8109 3440 8114 3496
rect 8170 3440 29274 3496
rect 29330 3440 29335 3496
rect 8109 3438 29335 3440
rect 8109 3435 8175 3438
rect 29269 3435 29335 3438
rect 5533 3362 5599 3365
rect 62 3360 5599 3362
rect 62 3304 5538 3360
rect 5594 3304 5599 3360
rect 62 3302 5599 3304
rect 62 2848 122 3302
rect 5533 3299 5599 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 8661 3226 8727 3229
rect 20713 3226 20779 3229
rect 8661 3224 20779 3226
rect 8661 3168 8666 3224
rect 8722 3168 20718 3224
rect 20774 3168 20779 3224
rect 8661 3166 20779 3168
rect 8661 3163 8727 3166
rect 20713 3163 20779 3166
rect 35341 3226 35407 3229
rect 39520 3226 40000 3256
rect 35341 3224 40000 3226
rect 35341 3168 35346 3224
rect 35402 3168 40000 3224
rect 35341 3166 40000 3168
rect 35341 3163 35407 3166
rect 39520 3136 40000 3166
rect 8293 2954 8359 2957
rect 17309 2954 17375 2957
rect 8293 2952 17375 2954
rect 8293 2896 8298 2952
rect 8354 2896 17314 2952
rect 17370 2896 17375 2952
rect 8293 2894 17375 2896
rect 8293 2891 8359 2894
rect 17309 2891 17375 2894
rect 0 2728 480 2848
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 7005 2682 7071 2685
rect 14089 2682 14155 2685
rect 7005 2680 14155 2682
rect 7005 2624 7010 2680
rect 7066 2624 14094 2680
rect 14150 2624 14155 2680
rect 7005 2622 14155 2624
rect 7005 2619 7071 2622
rect 14089 2619 14155 2622
rect 18597 2546 18663 2549
rect 27521 2546 27587 2549
rect 18597 2544 27587 2546
rect 18597 2488 18602 2544
rect 18658 2488 27526 2544
rect 27582 2488 27587 2544
rect 18597 2486 27587 2488
rect 18597 2483 18663 2486
rect 27521 2483 27587 2486
rect 33501 2410 33567 2413
rect 33501 2408 39682 2410
rect 33501 2352 33506 2408
rect 33562 2352 39682 2408
rect 33501 2350 39682 2352
rect 33501 2347 33567 2350
rect 7465 2274 7531 2277
rect 62 2272 7531 2274
rect 62 2216 7470 2272
rect 7526 2216 7531 2272
rect 62 2214 7531 2216
rect 62 1760 122 2214
rect 7465 2211 7531 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 39622 1896 39682 2350
rect 15377 1866 15443 1869
rect 32489 1866 32555 1869
rect 15377 1864 32555 1866
rect 15377 1808 15382 1864
rect 15438 1808 32494 1864
rect 32550 1808 32555 1864
rect 15377 1806 32555 1808
rect 15377 1803 15443 1806
rect 32489 1803 32555 1806
rect 39520 1776 40000 1896
rect 0 1640 480 1760
rect 1853 1186 1919 1189
rect 62 1184 1919 1186
rect 62 1128 1858 1184
rect 1914 1128 1919 1184
rect 62 1126 1919 1128
rect 62 672 122 1126
rect 1853 1123 1919 1126
rect 0 552 480 672
rect 39520 552 40000 672
rect 11881 98 11947 101
rect 39622 98 39682 552
rect 11881 96 39682 98
rect 11881 40 11886 96
rect 11942 40 39682 96
rect 11881 38 39682 40
rect 11881 35 11947 38
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 9628 11460 9692 11524
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 23428 10508 23492 10572
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 39620 6156 39684 6220
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 39620 5884 39684 5948
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 9630 10658 9690 11459
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 39619 6220 39685 6221
rect 39619 6156 39620 6220
rect 39684 6156 39685 6220
rect 39619 6155 39685 6156
rect 39622 5949 39682 6155
rect 39619 5948 39685 5949
rect 39619 5884 39620 5948
rect 39684 5884 39685 5948
rect 39619 5883 39685 5884
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 9542 10422 9778 10658
rect 23342 10572 23578 10658
rect 23342 10508 23428 10572
rect 23428 10508 23492 10572
rect 23492 10508 23578 10572
rect 23342 10422 23578 10508
<< metal5 >>
rect 9500 10658 23620 10700
rect 9500 10422 9542 10658
rect 9778 10422 23342 10658
rect 23578 10422 23620 10658
rect 9500 10380 23620 10422
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_37
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_49
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 774 592
use scs8hd_buf_1  _112_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_71 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__D
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_83
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 1142 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_86
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _191_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use scs8hd_buf_1  _174_
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_112
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_nor2_4  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _198_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_155
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_165
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 28152 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_298
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_320
timestamp 1586364061
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_324
timestamp 1586364061
transform 1 0 30912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_336
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_348
timestamp 1586364061
transform 1 0 33120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_360
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_14
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__C
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_8  _155_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_1  FILLER_2_99
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_109
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 15916 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_159
timestamp 1586364061
transform 1 0 15732 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_250
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_261
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_293
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 1142 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29716 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_2_313
timestamp 1586364061
transform 1 0 29900 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_317
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_327
timestamp 1586364061
transform 1 0 31188 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 32292 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 32660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_341
timestamp 1586364061
transform 1 0 32476 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_345
timestamp 1586364061
transform 1 0 32844 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_357
timestamp 1586364061
transform 1 0 33948 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_369
timestamp 1586364061
transform 1 0 35052 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_381
timestamp 1586364061
transform 1 0 36156 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_393
timestamp 1586364061
transform 1 0 37260 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_18
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use scs8hd_or2_4  _139_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _123_
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_166
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_224
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_228
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_248
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_268
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_272
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_285
timestamp 1586364061
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_289
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_296
timestamp 1586364061
transform 1 0 28336 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_300
timestamp 1586364061
transform 1 0 28704 0 1 3808
box -38 -48 314 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 29716 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_309
timestamp 1586364061
transform 1 0 29532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_313
timestamp 1586364061
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_317
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 31648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 32200 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 32016 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_334
timestamp 1586364061
transform 1 0 31832 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_347
timestamp 1586364061
transform 1 0 33028 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_365
timestamp 1586364061
transform 1 0 34684 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_371
timestamp 1586364061
transform 1 0 35236 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_383
timestamp 1586364061
transform 1 0 36340 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_395
timestamp 1586364061
transform 1 0 37444 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_21
timestamp 1586364061
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_1  _166_
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_or2_4  _076_
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 682 592
use scs8hd_decap_8  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 774 592
use scs8hd_or3_4  _111_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__C
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_99
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_6  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_233
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23368 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_244
timestamp 1586364061
transform 1 0 23552 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_264
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_268
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_283
timestamp 1586364061
transform 1 0 27140 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_287
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_290
timestamp 1586364061
transform 1 0 27784 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27876 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 29440 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_310
timestamp 1586364061
transform 1 0 29624 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 31188 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_320
timestamp 1586364061
transform 1 0 30544 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_326
timestamp 1586364061
transform 1 0 31096 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_329
timestamp 1586364061
transform 1 0 31372 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_333
timestamp 1586364061
transform 1 0 31740 0 -1 4896
box -38 -48 130 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 33672 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_346
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_350
timestamp 1586364061
transform 1 0 33304 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_357
timestamp 1586364061
transform 1 0 33948 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34684 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34408 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_364
timestamp 1586364061
transform 1 0 34592 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_368
timestamp 1586364061
transform 1 0 34960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_380
timestamp 1586364061
transform 1 0 36064 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_392
timestamp 1586364061
transform 1 0 37168 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_396
timestamp 1586364061
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 406 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_nor3_4  _152_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_120
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_144
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_261
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_277
timestamp 1586364061
transform 1 0 26588 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_280
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_284
timestamp 1586364061
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_297
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_301
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29440 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 31188 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 31004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_323
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_336
timestamp 1586364061
transform 1 0 32016 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_341
timestamp 1586364061
transform 1 0 32476 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_345
timestamp 1586364061
transform 1 0 32844 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_357
timestamp 1586364061
transform 1 0 33948 0 1 4896
box -38 -48 406 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_361
timestamp 1586364061
transform 1 0 34316 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_370
timestamp 1586364061
transform 1 0 35144 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_385
timestamp 1586364061
transform 1 0 36524 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_389
timestamp 1586364061
transform 1 0 36892 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_401
timestamp 1586364061
transform 1 0 37996 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_25
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_39
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_35
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _073_
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_inv_8  _096_
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 866 592
use scs8hd_or3_4  _121_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__C
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use scs8hd_nor3_4  _151_
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__C
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 130 592
use scs8hd_or2_4  _173_
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_121
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_192
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_196
timestamp 1586364061
transform 1 0 19136 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_6  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_206
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 27140 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 27048 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_280
timestamp 1586364061
transform 1 0 26864 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_279
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_292
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_300
timestamp 1586364061
transform 1 0 28704 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_304
timestamp 1586364061
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 29624 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_305
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_325
timestamp 1586364061
transform 1 0 31004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_321
timestamp 1586364061
transform 1 0 30636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_323
timestamp 1586364061
transform 1 0 30820 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_319
timestamp 1586364061
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_331
timestamp 1586364061
transform 1 0 31556 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 31372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 31188 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 31372 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 32292 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 32384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 32752 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_335
timestamp 1586364061
transform 1 0 31924 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_338
timestamp 1586364061
transform 1 0 32200 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33120 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 34132 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_350
timestamp 1586364061
transform 1 0 33304 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_356
timestamp 1586364061
transform 1 0 33856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_346
timestamp 1586364061
transform 1 0 32936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_357
timestamp 1586364061
transform 1 0 33948 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_360
timestamp 1586364061
transform 1 0 34224 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_371
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_361
timestamp 1586364061
transform 1 0 34316 0 1 5984
box -38 -48 314 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35972 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_382
timestamp 1586364061
transform 1 0 36248 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 36984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_388
timestamp 1586364061
transform 1 0 36800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_392
timestamp 1586364061
transform 1 0 37168 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_399
timestamp 1586364061
transform 1 0 37812 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_nand2_4  _097_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _131_
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__D
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _156_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_195
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_230
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_285
timestamp 1586364061
transform 1 0 27324 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_289
timestamp 1586364061
transform 1 0 27692 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 28520 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_297
timestamp 1586364061
transform 1 0 28428 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 30084 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 29532 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_307
timestamp 1586364061
transform 1 0 29348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_311
timestamp 1586364061
transform 1 0 29716 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_332
timestamp 1586364061
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33120 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_346
timestamp 1586364061
transform 1 0 32936 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_350
timestamp 1586364061
transform 1 0 33304 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35236 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_365
timestamp 1586364061
transform 1 0 34684 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_369
timestamp 1586364061
transform 1 0 35052 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_384
timestamp 1586364061
transform 1 0 36432 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_388
timestamp 1586364061
transform 1 0 36800 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_396
timestamp 1586364061
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__C
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_67
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _077_
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__D
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _142_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_9_206
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_277
timestamp 1586364061
transform 1 0 26588 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_294
timestamp 1586364061
transform 1 0 28152 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_298
timestamp 1586364061
transform 1 0 28520 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_315
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 31096 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 30912 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_321
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_337
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_343
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 36248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_63
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _141_
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_109
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_or2_4  _113_
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _124_
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_180
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_241
timestamp 1586364061
transform 1 0 23276 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_273
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 28888 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_291
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_299
timestamp 1586364061
transform 1 0 28612 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 29900 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_311
timestamp 1586364061
transform 1 0 29716 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_315
timestamp 1586364061
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_328
timestamp 1586364061
transform 1 0 31280 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32844 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 33028 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_10_358
timestamp 1586364061
transform 1 0 34040 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_363
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_376
timestamp 1586364061
transform 1 0 35696 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_388
timestamp 1586364061
transform 1 0 36800 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_139
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_218
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_278
timestamp 1586364061
transform 1 0 26680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 29808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 29624 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 31372 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_321
timestamp 1586364061
transform 1 0 30636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_325
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_340
timestamp 1586364061
transform 1 0 32384 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_344
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_393
timestamp 1586364061
transform 1 0 37260 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_397
timestamp 1586364061
transform 1 0 37628 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_405
timestamp 1586364061
transform 1 0 38364 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_or2_4  _165_
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use scs8hd_nor3_4  _150_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_103
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_192
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_223
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_233
timestamp 1586364061
transform 1 0 22540 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27692 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27416 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_279
timestamp 1586364061
transform 1 0 26772 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_284
timestamp 1586364061
transform 1 0 27232 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_298
timestamp 1586364061
transform 1 0 28520 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 29900 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 29256 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_308
timestamp 1586364061
transform 1 0 29440 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31096 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31464 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_332
timestamp 1586364061
transform 1 0 31648 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_341
timestamp 1586364061
transform 1 0 32476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_345
timestamp 1586364061
transform 1 0 32844 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 35328 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_364
timestamp 1586364061
transform 1 0 34592 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_383
timestamp 1586364061
transform 1 0 36340 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_387
timestamp 1586364061
transform 1 0 36708 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_391
timestamp 1586364061
transform 1 0 37076 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_14
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_17
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_25
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_21
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_nor3_4  _149_
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_81
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_85
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_146
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_228
timestamp 1586364061
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_249
timestamp 1586364061
transform 1 0 24012 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_250
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_257
timestamp 1586364061
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_288
timestamp 1586364061
transform 1 0 27600 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_285
timestamp 1586364061
transform 1 0 27324 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_289
timestamp 1586364061
transform 1 0 27692 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_292
timestamp 1586364061
transform 1 0 27968 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_295
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_299
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_302
timestamp 1586364061
transform 1 0 28888 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 30084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_315
timestamp 1586364061
transform 1 0 30084 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_314
timestamp 1586364061
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 31004 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_319
timestamp 1586364061
transform 1 0 30452 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_328
timestamp 1586364061
transform 1 0 31280 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32844 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_333
timestamp 1586364061
transform 1 0 31740 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_355
timestamp 1586364061
transform 1 0 33764 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_359
timestamp 1586364061
transform 1 0 34132 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_354
timestamp 1586364061
transform 1 0 33672 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_358
timestamp 1586364061
transform 1 0 34040 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_371
timestamp 1586364061
transform 1 0 35236 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_381
timestamp 1586364061
transform 1 0 36156 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_375
timestamp 1586364061
transform 1 0 35604 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_397
timestamp 1586364061
transform 1 0 37628 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_170
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_249
timestamp 1586364061
transform 1 0 24012 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_280
timestamp 1586364061
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29808 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 31004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_323
timestamp 1586364061
transform 1 0 30820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_327
timestamp 1586364061
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_340
timestamp 1586364061
transform 1 0 32384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_344
timestamp 1586364061
transform 1 0 32752 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_351
timestamp 1586364061
transform 1 0 33396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_355
timestamp 1586364061
transform 1 0 33764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_359
timestamp 1586364061
transform 1 0 34132 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_380
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_387
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_398
timestamp 1586364061
transform 1 0 37720 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_402
timestamp 1586364061
transform 1 0 38088 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_406
timestamp 1586364061
transform 1 0 38456 0 1 10336
box -38 -48 130 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 590 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_111
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_115
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_221
timestamp 1586364061
transform 1 0 21436 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_233
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_252
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_264
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_269
timestamp 1586364061
transform 1 0 25852 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_285
timestamp 1586364061
transform 1 0 27324 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_293
timestamp 1586364061
transform 1 0 28060 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_297
timestamp 1586364061
transform 1 0 28428 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 30084 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_309
timestamp 1586364061
transform 1 0 29532 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_314
timestamp 1586364061
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_341
timestamp 1586364061
transform 1 0 32476 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33304 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_353
timestamp 1586364061
transform 1 0 33580 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_370
timestamp 1586364061
transform 1 0 35144 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35880 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_374
timestamp 1586364061
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_381
timestamp 1586364061
transform 1 0 36156 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_393
timestamp 1586364061
transform 1 0 37260 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_or3_4  _084_
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _069_
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use scs8hd_inv_8  _154_
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_194
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_211
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_248
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_252
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 26220 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_265
timestamp 1586364061
transform 1 0 25484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 27784 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27232 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_282
timestamp 1586364061
transform 1 0 27048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_286
timestamp 1586364061
transform 1 0 27416 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 28244 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_297
timestamp 1586364061
transform 1 0 28428 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30728 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_325
timestamp 1586364061
transform 1 0 31004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_329
timestamp 1586364061
transform 1 0 31372 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 31740 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_336
timestamp 1586364061
transform 1 0 32016 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_348
timestamp 1586364061
transform 1 0 33120 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_352
timestamp 1586364061
transform 1 0 33488 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35328 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_371
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_375
timestamp 1586364061
transform 1 0 35604 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_183
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 20976 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23000 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_241
timestamp 1586364061
transform 1 0 23276 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 25116 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_253
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_258
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_265
timestamp 1586364061
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_273
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_279
timestamp 1586364061
transform 1 0 26772 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 27968 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_291
timestamp 1586364061
transform 1 0 27876 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_295
timestamp 1586364061
transform 1 0 28244 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_307
timestamp 1586364061
transform 1 0 29348 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_319
timestamp 1586364061
transform 1 0 30452 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_331
timestamp 1586364061
transform 1 0 31556 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_335
timestamp 1586364061
transform 1 0 31924 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_353
timestamp 1586364061
transform 1 0 33580 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_357
timestamp 1586364061
transform 1 0 33948 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34684 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_368
timestamp 1586364061
transform 1 0 34960 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_380
timestamp 1586364061
transform 1 0 36064 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_392
timestamp 1586364061
transform 1 0 37168 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_396
timestamp 1586364061
transform 1 0 37536 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  _085_
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _153_
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_91
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 590 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_185
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_221
timestamp 1586364061
transform 1 0 21436 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_233
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_245
timestamp 1586364061
transform 1 0 23644 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26128 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_264
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_268
timestamp 1586364061
transform 1 0 25760 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26588 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_279
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_291
timestamp 1586364061
transform 1 0 27876 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_303
timestamp 1586364061
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 29808 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_310
timestamp 1586364061
transform 1 0 29624 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_314
timestamp 1586364061
transform 1 0 29992 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_326
timestamp 1586364061
transform 1 0 31096 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_338
timestamp 1586364061
transform 1 0 32200 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_350
timestamp 1586364061
transform 1 0 33304 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_362
timestamp 1586364061
transform 1 0 34408 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 552 480 672 6 address[0]
port 0 nsew default input
rlabel metal2 s 1214 15520 1270 16000 6 address[1]
port 1 nsew default input
rlabel metal2 s 3698 15520 3754 16000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 1640 480 1760 6 address[3]
port 3 nsew default input
rlabel metal2 s 6182 15520 6238 16000 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 2728 480 2848 6 address[5]
port 5 nsew default input
rlabel metal2 s 8666 15520 8722 16000 6 address[6]
port 6 nsew default input
rlabel metal2 s 11150 15520 11206 16000 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 13634 15520 13690 16000 6 bottom_grid_pin_4_
port 8 nsew default tristate
rlabel metal3 s 39520 552 40000 672 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal3 s 39520 1776 40000 1896 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal2 s 16210 15520 16266 16000 6 chanx_left_in[1]
port 11 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[2]
port 12 nsew default input
rlabel metal2 s 18694 15520 18750 16000 6 chanx_left_in[3]
port 13 nsew default input
rlabel metal3 s 39520 3136 40000 3256 6 chanx_left_in[4]
port 14 nsew default input
rlabel metal2 s 21178 15520 21234 16000 6 chanx_left_in[5]
port 15 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chanx_left_in[6]
port 16 nsew default input
rlabel metal3 s 39520 4496 40000 4616 6 chanx_left_in[7]
port 17 nsew default input
rlabel metal3 s 39520 5856 40000 5976 6 chanx_left_in[8]
port 18 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chanx_left_out[0]
port 19 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[1]
port 20 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 chanx_left_out[2]
port 21 nsew default tristate
rlabel metal2 s 23662 15520 23718 16000 6 chanx_left_out[3]
port 22 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chanx_left_out[4]
port 23 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chanx_left_out[5]
port 24 nsew default tristate
rlabel metal3 s 39520 7216 40000 7336 6 chanx_left_out[6]
port 25 nsew default tristate
rlabel metal3 s 39520 8576 40000 8696 6 chanx_left_out[7]
port 26 nsew default tristate
rlabel metal2 s 26146 15520 26202 16000 6 chanx_left_out[8]
port 27 nsew default tristate
rlabel metal3 s 39520 9800 40000 9920 6 chanx_right_in[0]
port 28 nsew default input
rlabel metal2 s 21362 0 21418 480 6 chanx_right_in[1]
port 29 nsew default input
rlabel metal2 s 28722 15520 28778 16000 6 chanx_right_in[2]
port 30 nsew default input
rlabel metal2 s 31206 15520 31262 16000 6 chanx_right_in[3]
port 31 nsew default input
rlabel metal3 s 39520 11160 40000 11280 6 chanx_right_in[4]
port 32 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_right_in[5]
port 33 nsew default input
rlabel metal3 s 39520 12520 40000 12640 6 chanx_right_in[6]
port 34 nsew default input
rlabel metal2 s 24214 0 24270 480 6 chanx_right_in[7]
port 35 nsew default input
rlabel metal2 s 27066 0 27122 480 6 chanx_right_in[8]
port 36 nsew default input
rlabel metal2 s 33690 15520 33746 16000 6 chanx_right_out[0]
port 37 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 39520 13880 40000 14000 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal2 s 36174 15520 36230 16000 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 0 10752 480 10872 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal2 s 29918 0 29974 480 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal2 s 4250 0 4306 480 6 data_in
port 46 nsew default input
rlabel metal2 s 1398 0 1454 480 6 enable
port 47 nsew default input
rlabel metal3 s 39520 15240 40000 15360 6 top_grid_pin_0_
port 48 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 top_grid_pin_10_
port 49 nsew default tristate
rlabel metal2 s 38658 15520 38714 16000 6 top_grid_pin_12_
port 50 nsew default tristate
rlabel metal2 s 38474 0 38530 480 6 top_grid_pin_14_
port 51 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 top_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 32770 0 32826 480 6 top_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 top_grid_pin_6_
port 54 nsew default tristate
rlabel metal2 s 35622 0 35678 480 6 top_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< end >>
