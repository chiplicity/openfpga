* NGSPICE file created from sb_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_0__1_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk right_bottom_grid_pin_34_ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_
+ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_
+ right_bottom_grid_pin_41_ top_left_grid_pin_1_ VPWR VGND
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X _067_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_114_ chany_bottom_in[10] chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _104_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_20.mux_l1_in_1_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_113_ _113_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l3_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S mux_right_track_10.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_112_ chany_bottom_in[12] chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_10.mux_l2_in_1_ _061_/HI chany_bottom_in[9] mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_17.mux_l3_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_7 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l3_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_10.mux_l2_in_0_ right_bottom_grid_pin_35_ mux_right_track_10.mux_l1_in_0_/X
+ mux_right_track_10.mux_l2_in_0_/S mux_right_track_10.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_111_ chany_bottom_in[13] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_8 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_12.mux_l2_in_1_/S
+ mux_right_track_12.mux_l3_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ _045_/HI chany_bottom_in[8] mux_right_track_8.mux_l2_in_1_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l2_in_1_ _046_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[12] chany_bottom_in[2] mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X _117_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ chany_bottom_in[14] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_8.mux_l3_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X _125_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l2_in_1_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_10.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_34_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S mux_right_track_22.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_0.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_22.mux_l1_in_1_ _035_/HI chany_bottom_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_1_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l3_in_0_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l3_in_0_/X _080_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_10.mux_l3_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_22.mux_l1_in_0_ right_bottom_grid_pin_41_ chany_top_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_1_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_34.mux_l2_in_0_ _041_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _081_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l2_in_1_ _055_/HI chanx_right_in[14] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l2_in_0_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_099_ chany_top_in[5] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l2_in_1_ _059_/HI mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _069_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _072_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_18.mux_l1_in_1_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.mux_l1_in_0_ chany_bottom_in[1] right_bottom_grid_pin_39_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_098_ chany_top_in[6] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_0_/S mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[7] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[2] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_1_ _047_/HI chany_bottom_in[17] mux_top_track_16.mux_l2_in_0_/S
+ mux_top_track_16.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_097_ _097_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_1_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_1_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _101_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_096_ chany_top_in[8] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_4.mux_l1_in_2_/S mux_top_track_4.mux_l2_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_079_ _079_/A chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_3_ _043_/HI chany_bottom_in[5] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[8] chanx_right_in[19] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_095_ chany_top_in[9] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_078_ _078_/A chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_4.mux_l1_in_3_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[5] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_3_/S mux_right_track_4.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_094_ chany_top_in[10] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_077_ _077_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_1_ _064_/HI chany_bottom_in[13] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_4.mux_l1_in_3_/S mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l2_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_3_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ _093_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
X_076_ _076_/A chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ chany_top_in[13] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_3_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_28.mux_l2_in_0_ _038_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_30.mux_l2_in_0_ _039_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_20.mux_l2_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l2_in_1_ _058_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_092_ chany_top_in[12] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[17] mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_075_ _075_/A chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_28.mux_l1_in_0_ chany_bottom_in[11] right_bottom_grid_pin_36_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_30.mux_l1_in_0_ chany_bottom_in[7] right_bottom_grid_pin_37_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ chany_top_in[13] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_074_ _074_/A chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[3] mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_109_ _109_/A chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ ccff_tail mux_bottom_track_33.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l2_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_090_ chany_top_in[14] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_33.mux_l1_in_1_ _057_/HI chanx_right_in[13] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_2_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_073_ _073_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_125_ _125_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ chany_bottom_in[16] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_14.mux_l2_in_1_/S
+ mux_right_track_14.mux_l3_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_2_/S clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_24.mux_l2_in_1_ _049_/HI chany_bottom_in[18] mux_top_track_24.mux_l2_in_1_/S
+ mux_top_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[6] chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_072_ _072_/A chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 _065_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ _124_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S mux_right_track_12.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_107_ chany_bottom_in[17] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_12.mux_l2_in_1_ _062_/HI chany_bottom_in[10] mux_right_track_12.mux_l2_in_1_/S
+ mux_right_track_12.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_1_ _060_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l2_in_1_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[2] right_bottom_grid_pin_40_ mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_24.mux_l2_in_0_ chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_1_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_071_ _071_/A chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_123_ _123_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_106_ chany_bottom_in[18] chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_12.mux_l2_in_0_ right_bottom_grid_pin_36_ mux_right_track_12.mux_l1_in_0_/X
+ mux_right_track_12.mux_l2_in_1_/S mux_right_track_12.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_12.mux_l3_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_38_ right_bottom_grid_pin_36_
+ mux_right_track_0.mux_l1_in_2_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ _036_/HI chany_bottom_in[19] mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ _048_/HI chany_bottom_in[13] mux_top_track_2.mux_l2_in_1_/S
+ mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_070_ _070_/A chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ chany_bottom_in[2] chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[6] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_105_ _105_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_12.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[2] mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _124_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_24.mux_l2_in_0_ chany_bottom_in[18] mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_1_ chany_bottom_in[4] chanx_right_in[16] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_121_ _121_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_104_ _104_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ _053_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l3_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[19] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_0.mux_l1_in_1_/S mux_top_track_0.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[18] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_0_ chanx_right_in[9] chanx_right_in[2] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_120_ chany_bottom_in[4] chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_36.mux_l2_in_0_ _042_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_103_ _103_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[5] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X _068_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_track_0.mux_l1_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X _071_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_102_ chany_top_in[2] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_36.mux_l1_in_0_ chany_bottom_in[0] right_bottom_grid_pin_40_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_2_/S mux_right_track_0.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_101_ _101_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_32.mux_l3_in_0_/S mux_right_track_0.mux_l1_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l2_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_100_ chany_top_in[4] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S mux_top_track_32.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_6.mux_l1_in_3_ _044_/HI chany_bottom_in[6] mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_32.mux_l2_in_1_ _050_/HI chany_bottom_in[10] mux_top_track_32.mux_l2_in_0_/S
+ mux_top_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_6.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l3_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_32.mux_l2_in_0_ chanx_right_in[14] mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_0_/S mux_top_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_22.mux_l2_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/S clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S mux_right_track_18.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_089_ _089_/A chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S mux_right_track_20.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_18.mux_l1_in_1_ _065_/HI chany_bottom_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l2_in_0_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_20.mux_l1_in_1_ _034_/HI chany_bottom_in[16] mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_1_ _052_/HI mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_32.mux_l1_in_0_ chanx_right_in[7] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_088_ chany_top_in[16] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_18.mux_l1_in_0_ right_bottom_grid_pin_39_ chany_top_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_6.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_0_ right_bottom_grid_pin_40_ chany_top_in[16] mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_36.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l1_in_1_/S clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_32.mux_l2_in_0_ _040_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _121_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[11] mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X _070_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_087_ chany_top_in[17] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[4] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_1_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_32.mux_l2_in_0_/S mux_top_track_32.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[3] right_bottom_grid_pin_38_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ chany_top_in[18] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_069_ _069_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l3_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l2_in_0_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _085_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_068_ _068_/A chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_14.mux_l3_in_0_/S
+ mux_right_track_16.mux_l1_in_1_/S clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_24.mux_l3_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l1_in_3_ _033_/HI chany_bottom_in[4] mux_right_track_2.mux_l1_in_2_/S
+ mux_right_track_2.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_084_ _084_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_067_ _067_/A chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_119_ chany_bottom_in[5] chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S mux_right_track_14.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_14.mux_l2_in_1_ _063_/HI chany_bottom_in[12] mux_right_track_14.mux_l2_in_1_/S
+ mux_right_track_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_083_ _083_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_2.mux_l1_in_2_/S mux_right_track_2.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_066_ right_bottom_grid_pin_41_ chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_118_ chany_bottom_in[6] chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_33.mux_l1_in_1_/S
+ ccff_tail clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_14.mux_l2_in_0_ right_bottom_grid_pin_37_ mux_right_track_14.mux_l1_in_0_/X
+ mux_right_track_14.mux_l2_in_1_/S mux_right_track_14.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ _082_/A chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_4.mux_l2_in_1_ _051_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_2.mux_l1_in_2_/S mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/S clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_117_ _117_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_4.mux_l1_in_2_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_2 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_33.mux_l1_in_1_/S clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_24.mux_l2_in_1_/S mux_top_track_24.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_14.mux_l1_in_0_ chany_top_in[19] chany_top_in[12] mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_081_ _081_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _084_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_2_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_0.mux_l3_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_26.mux_l2_in_0_ _037_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _123_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.mux_l2_in_1_ _054_/HI chanx_right_in[15] mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ chanx_right_in[17] chanx_right_in[10] mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_116_ chany_bottom_in[8] chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_8.mux_l1_in_1_/S mux_top_track_8.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ _056_/HI chanx_right_in[18] mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_2_/S mux_right_track_2.mux_l2_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l3_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_080_ _080_/A chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_2_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_115_ chany_bottom_in[9] chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[15] right_bottom_grid_pin_35_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_4 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_16.mux_l3_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

