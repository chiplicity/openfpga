* NGSPICE file created from sb_0__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

.subckt sb_0__0_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] prog_clk right_bottom_grid_pin_11_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ top_left_grid_pin_1_ VPWR VGND
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.mux_l1_in_0__S mux_right_track_18.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_66_ chanx_right_in[14] chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_49_ chany_top_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_65_ chanx_right_in[15] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_48_ chany_top_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_10.mux_l2_in_0__A1 mux_right_track_10.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A mux_right_track_28.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_64_ chanx_right_in[16] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_14.mux_l1_in_0__S mux_right_track_14.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A mux_top_track_0.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0__S mux_right_track_6.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0__A1 mux_right_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_63_ chanx_right_in[17] chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ _46_/A chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.mux_l2_in_0_ _28_/HI mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_62_ chanx_right_in[18] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_45_ _45_/A chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_10.mux_l1_in_0__S mux_right_track_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l2_in_0_/X _79_/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[4] mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l2_in_0_ _22_/HI mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ _23_/HI mux_top_track_0.mux_l1_in_0_/X mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_30.mux_l1_in_0__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_61_ chanx_right_in[19] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_44_ _44_/A chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l2_in_0_/X _54_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A mux_right_track_14.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[3] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__42__A _42_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l2_in_1__S mux_right_track_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_60_ chanx_right_in[0] chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_18.mux_l1_in_0_/S
+ mux_right_track_18.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_34.mux_l2_in_0_ _39_/HI mux_right_track_34.mux_l1_in_0_/X ccff_tail
+ mux_right_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l2_in_0_/X _55_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_43_ _43_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__50__A _50_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_34.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _43_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_33_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__45__A _45_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_28.mux_l1_in_0__S mux_right_track_28.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _46_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_18.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__53__A _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_42_ _42_/A chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.mux_l1_in_0_ right_bottom_grid_pin_11_ chany_top_in[16] mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__48__A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 _38_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__61__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A mux_right_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__56__A _56_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_41_ chany_top_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__64__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__59__A _59_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_30.mux_l2_in_0__S mux_right_track_30.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__72__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__67__A _67_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.mux_l1_in_0__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_40_ chany_top_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__75__A _75_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__78__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l3_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.mux_l2_in_1_ _20_/HI right_bottom_grid_pin_9_ mux_right_track_4.mux_l2_in_1_/S
+ mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_0.mux_l2_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_36_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 right_bottom_grid_pin_7_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_0_/S mux_right_track_4.mux_l2_in_1_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l2_in_0_ _31_/HI mux_right_track_16.mux_l1_in_0_/X mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ right_bottom_grid_pin_5_ mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__S mux_right_track_12.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_9_ chany_top_in[7] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[1] mux_right_track_4.mux_l1_in_0_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_28.mux_l2_in_0_ _36_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _57_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_30.mux_l2_in_0_ _37_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 _20_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_79_ _79_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _51_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ right_bottom_grid_pin_5_ chany_top_in[13] mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_30.mux_l1_in_0_ right_bottom_grid_pin_7_ chany_top_in[14] mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_78_ chanx_right_in[2] chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ _77_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__A1 mux_right_track_12.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 _22_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l1_in_0__S mux_right_track_34.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_76_ chanx_right_in[4] chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A mux_right_track_10.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_26.mux_l2_in_0__S mux_right_track_26.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ _59_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A mux_top_track_8.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_1_ _27_/HI right_bottom_grid_pin_9_ mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_75_ _75_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.mux_l2_in_0_ _24_/HI mux_top_track_24.mux_l1_in_0_/X mux_top_track_24.mux_l2_in_0_/S
+ mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__40__A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_58_ _58_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_30.mux_l1_in_0__S mux_right_track_30.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_12.mux_l2_in_0_ _29_/HI mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_0_ right_bottom_grid_pin_5_ mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__43__A _43_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_74_ chanx_right_in[6] chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _67_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_57_ _57_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__51__A _51_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_1_ mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__46__A _46_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _59_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.mux_l1_in_0_ right_bottom_grid_pin_5_ chany_top_in[5] mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[19] mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l2_in_0_ _34_/HI mux_right_track_24.mux_l1_in_0_/X mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__54__A _54_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_73_ chanx_right_in[7] chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__49__A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_56_ _56_/A chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A0 _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_39_ _39_/HI _39_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__62__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__57__A _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l2_in_0_/X _53_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__70__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ chanx_right_in[8] chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_26.mux_l2_in_0__A0 _35_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l3_in_0__S mux_right_track_6.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__65__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_55_ _55_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_1_ chany_top_in[11] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A mux_right_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.mux_l2_in_0__A1 mux_right_track_18.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ _38_/HI _38_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__73__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__S mux_right_track_12.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__68__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X _42_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_34.mux_l2_in_0__A0 _39_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_71_ chanx_right_in[9] chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_track_0.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_26.mux_l2_in_0__A1 mux_right_track_26.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_54_ _54_/A chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X _45_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__76__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ _37_/HI _37_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l2_in_0__A1 mux_right_track_34.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__79__A _79_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_70_ chanx_right_in[10] chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_53_ _53_/A chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l3_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_36_ _36_/HI _36_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 right_bottom_grid_pin_9_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_24.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_52_ _52_/A chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_6.mux_l1_in_0_/S mux_right_track_6.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_35_ _35_/HI _35_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_51_ _51_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_34_ _34_/HI _34_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ _21_/HI right_bottom_grid_pin_11_ mux_right_track_6.mux_l2_in_0_/S
+ mux_right_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 _23_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A mux_right_track_26.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_50_ _50_/A chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_26.mux_l1_in_0__S mux_right_track_26.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_18.mux_l2_in_0_ _32_/HI mux_right_track_18.mux_l1_in_0_/X mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ right_bottom_grid_pin_7_ mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A mux_top_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_18.mux_l2_in_0__S mux_right_track_18.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A0 _21_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.mux_l1_in_0_ right_bottom_grid_pin_11_ chany_top_in[8] mux_right_track_18.mux_l1_in_0_/S
+ mux_right_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_6.mux_l3_in_0__A0 mux_right_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[2] mux_right_track_6.mux_l1_in_0_/S
+ mux_right_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_0_ _26_/HI mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_32.mux_l2_in_0_ _38_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _56_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X _75_/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A mux_top_track_4.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X _44_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l2_in_0_/X _47_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_6.mux_l3_in_0__A1 mux_right_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _50_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[5] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_32.mux_l1_in_0_ right_bottom_grid_pin_9_ chany_top_in[15] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0__S mux_right_track_14.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A mux_right_track_12.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0__A1 mux_right_track_14.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__41__A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0__S mux_right_track_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_30.mux_l2_in_0__A0 _37_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__44__A _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A mux_right_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_30.mux_l2_in_0__A1 mux_right_track_30.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__52__A _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0__S mux_right_track_10.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__47__A _47_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 right_bottom_grid_pin_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__60__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__55__A _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l2_in_1_ _33_/HI right_bottom_grid_pin_11_ mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A mux_right_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_34.mux_l1_in_0__A0 right_bottom_grid_pin_11_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__63__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_34.mux_l1_in_0_/S
+ ccff_tail prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__58__A _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__71__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_14.mux_l2_in_0_ _30_/HI mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_0_ right_bottom_grid_pin_7_ mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__66__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 right_bottom_grid_pin_5_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_69_ chanx_right_in[11] chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_34.mux_l1_in_0__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/S prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__74__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.mux_l2_in_0__S mux_right_track_28.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__69__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l3_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _58_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_14.mux_l1_in_0_ right_bottom_grid_pin_7_ chany_top_in[6] mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__77__A _77_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[0] mux_right_track_2.mux_l1_in_0_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l2_in_0_ _25_/HI mux_top_track_4.mux_l1_in_0_/X mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ _35_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_68_ chanx_right_in[12] chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l2_in_0_/X _77_/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_28.mux_l2_in_0__A0 _36_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_0_/S mux_right_track_2.mux_l2_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l2_in_0_/X _52_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_67_ _67_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 right_bottom_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.mux_l2_in_0__A1 mux_right_track_28.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_26.mux_l1_in_0_ right_bottom_grid_pin_3_ chany_top_in[12] mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_4.mux_l2_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_8.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

