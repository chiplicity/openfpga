* NGSPICE file created from sb_0__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_0__0_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] prog_clk right_bottom_grid_pin_1_
+ right_top_grid_pin_42_ right_top_grid_pin_43_ right_top_grid_pin_44_ right_top_grid_pin_45_
+ right_top_grid_pin_46_ right_top_grid_pin_47_ right_top_grid_pin_48_ right_top_grid_pin_49_
+ top_left_grid_pin_1_ vpwr vgnd
XFILLER_26_74 vgnd vpwr scs8hd_decap_12
XFILLER_13_166 vgnd vpwr scs8hd_decap_12
XFILLER_3_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l1_in_0__S mux_right_track_18.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_247 vpwr vgnd scs8hd_fill_2
XFILLER_10_147 vgnd vpwr scs8hd_decap_12
XFILLER_12_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_236 vgnd vpwr scs8hd_decap_8
XFILLER_18_225 vgnd vpwr scs8hd_fill_1
X_66_ chanx_right_in[10] chany_top_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_24_239 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_18.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_16.mux_l2_in_0_/S mux_right_track_18.mux_l1_in_0_/S
+ mem_right_track_18.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_272 vgnd vpwr scs8hd_decap_3
XFILLER_15_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_44 vgnd vpwr scs8hd_decap_12
X_49_ _49_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_20_253 vpwr vgnd scs8hd_fill_2
XFILLER_18_86 vgnd vpwr scs8hd_decap_12
XFILLER_34_74 vgnd vpwr scs8hd_decap_12
XFILLER_37_161 vpwr vgnd scs8hd_fill_2
XFILLER_20_98 vgnd vpwr scs8hd_decap_12
XFILLER_19_150 vgnd vpwr scs8hd_decap_3
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_175 vgnd vpwr scs8hd_decap_8
XFILLER_34_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_15_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_156 vgnd vpwr scs8hd_decap_8
XFILLER_40_123 vgnd vpwr scs8hd_decap_12
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_263 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_145 vpwr vgnd scs8hd_fill_2
XFILLER_31_167 vpwr vgnd scs8hd_fill_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_223 vpwr vgnd scs8hd_fill_2
XFILLER_22_167 vgnd vpwr scs8hd_decap_12
XFILLER_22_156 vgnd vpwr scs8hd_decap_8
XFILLER_22_123 vgnd vpwr scs8hd_decap_3
Xmem_right_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_86 vgnd vpwr scs8hd_decap_12
XFILLER_9_105 vgnd vpwr scs8hd_decap_12
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_178 vgnd vpwr scs8hd_decap_12
XFILLER_3_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_171 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_10_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 _24_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_218 vpwr vgnd scs8hd_fill_2
XFILLER_18_259 vgnd vpwr scs8hd_decap_12
XFILLER_41_251 vgnd vpwr scs8hd_decap_8
XFILLER_5_141 vgnd vpwr scs8hd_decap_12
X_65_ chanx_right_in[11] chany_top_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_23_251 vpwr vgnd scs8hd_fill_2
XFILLER_23_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D mux_right_track_18.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_12
X_48_ _48_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_20_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_98 vgnd vpwr scs8hd_decap_12
XFILLER_34_86 vgnd vpwr scs8hd_decap_12
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_107 vgnd vpwr scs8hd_decap_12
XFILLER_37_184 vpwr vgnd scs8hd_fill_2
XFILLER_20_22 vgnd vpwr scs8hd_decap_12
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XFILLER_28_162 vgnd vpwr scs8hd_decap_12
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XFILLER_40_135 vpwr vgnd scs8hd_fill_2
XFILLER_15_44 vgnd vpwr scs8hd_decap_12
XFILLER_31_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XFILLER_16_110 vgnd vpwr scs8hd_decap_12
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_0_/S
+ mem_right_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_98 vgnd vpwr scs8hd_decap_12
XFILLER_9_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.scs8hd_buf_4_0__A mux_right_track_12.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_27_205 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_20.mux_l2_in_0__S mux_right_track_20.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0__A1 mux_right_track_10.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_208 vpwr vgnd scs8hd_fill_2
XFILLER_41_263 vpwr vgnd scs8hd_fill_2
X_64_ chanx_right_in[12] chany_top_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A0 mux_right_track_6.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__S mux_right_track_14.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_123 vgnd vpwr scs8hd_decap_12
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_68 vgnd vpwr scs8hd_decap_12
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
X_47_ _47_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_34_98 vgnd vpwr scs8hd_fill_1
XFILLER_11_255 vgnd vpwr scs8hd_decap_12
XFILLER_7_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_119 vgnd vpwr scs8hd_decap_3
XFILLER_37_196 vgnd vpwr scs8hd_decap_4
XFILLER_1_80 vgnd vpwr scs8hd_decap_12
XFILLER_20_34 vgnd vpwr scs8hd_decap_12
XFILLER_29_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_251 vpwr vgnd scs8hd_fill_2
Xmem_right_track_26.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_26.mux_l1_in_0_/S ccff_tail
+ mem_right_track_26.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_19_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D mux_right_track_0.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_122 vpwr vgnd scs8hd_fill_2
XFILLER_15_56 vgnd vpwr scs8hd_decap_12
XFILLER_31_44 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_103 vpwr vgnd scs8hd_fill_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_129 vgnd vpwr scs8hd_decap_12
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_184 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.scs8hd_buf_4_0_ mux_right_track_12.mux_l2_in_0_/X _49_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_27_228 vgnd vpwr scs8hd_decap_4
XFILLER_35_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_228 vpwr vgnd scs8hd_fill_2
XFILLER_18_217 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l1_in_0__S mux_right_track_6.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0__A1 mux_right_track_6.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_63_ _63_/A chany_top_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_23_264 vgnd vpwr scs8hd_decap_8
XFILLER_23_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_253 vpwr vgnd scs8hd_fill_2
XFILLER_14_220 vgnd vpwr scs8hd_decap_12
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
X_46_ _46_/A chanx_right_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_20_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_267 vgnd vpwr scs8hd_decap_8
XFILLER_7_227 vgnd vpwr scs8hd_decap_12
XFILLER_7_205 vgnd vpwr scs8hd_decap_4
Xmux_right_track_10.mux_l2_in_0_ _24_/HI mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
X_29_ _29_/HI _29_/LO vgnd vpwr scs8hd_conb_1
XFILLER_4_208 vgnd vpwr scs8hd_decap_12
XFILLER_29_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_46 vgnd vpwr scs8hd_decap_12
XFILLER_6_59 vpwr vgnd scs8hd_fill_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_263 vgnd vpwr scs8hd_decap_12
Xmem_right_track_26.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_24.mux_l2_in_0_/S mux_right_track_26.mux_l1_in_0_/S
+ mem_right_track_26.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_34_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D mux_right_track_20.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_68 vgnd vpwr scs8hd_decap_12
XFILLER_31_56 vgnd vpwr scs8hd_decap_12
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XFILLER_16_123 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_20.scs8hd_buf_4_0_ mux_right_track_20.mux_l2_in_0_/X _45_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_39_215 vgnd vpwr scs8hd_decap_4
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_80 vgnd vpwr scs8hd_decap_12
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_27 vgnd vpwr scs8hd_decap_4
XFILLER_36_229 vgnd vpwr scs8hd_decap_4
XFILLER_8_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D mux_right_track_2.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_37_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_166 vgnd vpwr scs8hd_decap_12
X_62_ chanx_right_in[14] chany_top_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_17_251 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
X_45_ _45_/A chanx_right_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_20_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D mux_right_track_20.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0__S mux_right_track_10.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_202 vgnd vpwr scs8hd_decap_12
XFILLER_7_239 vgnd vpwr scs8hd_decap_12
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
X_28_ _28_/HI _28_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_132 vpwr vgnd scs8hd_fill_2
XFILLER_37_154 vgnd vpwr scs8hd_decap_4
XFILLER_1_93 vgnd vpwr scs8hd_decap_12
XFILLER_20_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_176 vgnd vpwr scs8hd_decap_6
XFILLER_28_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_19_154 vpwr vgnd scs8hd_fill_2
XFILLER_25_157 vgnd vpwr scs8hd_decap_12
XFILLER_31_68 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_ right_top_grid_pin_43_ chany_top_in[4] mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_149 vpwr vgnd scs8hd_fill_2
XFILLER_16_135 vgnd vpwr scs8hd_decap_12
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ _19_/HI mux_top_track_0.mux_l1_in_0_/X mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_22.mux_l2_in_0_ _31_/HI mux_right_track_22.mux_l1_in_0_/X mux_right_track_22.mux_l2_in_0_/S
+ mux_right_track_22.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_238 vpwr vgnd scs8hd_fill_2
XFILLER_39_227 vgnd vpwr scs8hd_decap_8
XFILLER_30_171 vgnd vpwr scs8hd_fill_1
XFILLER_15_190 vgnd vpwr scs8hd_decap_12
XFILLER_30_193 vgnd vpwr scs8hd_decap_4
XFILLER_13_105 vgnd vpwr scs8hd_decap_12
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_12_171 vgnd vpwr scs8hd_decap_12
XFILLER_12_59 vpwr vgnd scs8hd_fill_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_ _18_/HI right_bottom_grid_pin_1_ mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_56 vgnd vpwr scs8hd_decap_12
XFILLER_26_274 vgnd vpwr scs8hd_decap_3
XFILLER_26_241 vgnd vpwr scs8hd_decap_3
XFILLER_5_178 vgnd vpwr scs8hd_decap_12
X_61_ chanx_right_in[15] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_222 vpwr vgnd scs8hd_fill_2
XFILLER_2_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_80 vgnd vpwr scs8hd_decap_12
X_44_ _44_/A chanx_right_out[11] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_20.scs8hd_buf_4_0__A mux_right_track_20.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D mux_right_track_6.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
X_27_ _27_/HI _27_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_188 vpwr vgnd scs8hd_fill_2
XFILLER_29_68 vgnd vpwr scs8hd_decap_12
XFILLER_28_188 vpwr vgnd scs8hd_fill_2
XFILLER_6_39 vgnd vpwr scs8hd_decap_12
XFILLER_3_276 vgnd vpwr scs8hd_fill_1
XFILLER_34_114 vgnd vpwr scs8hd_decap_8
XFILLER_19_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_106 vgnd vpwr scs8hd_fill_1
XFILLER_25_169 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_147 vgnd vpwr scs8hd_decap_12
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_206 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_93 vgnd vpwr scs8hd_decap_12
XFILLER_13_117 vgnd vpwr scs8hd_decap_12
XFILLER_29_261 vpwr vgnd scs8hd_fill_2
XFILLER_8_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_264 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[3] mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D mux_right_track_8.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_68 vgnd vpwr scs8hd_decap_12
XFILLER_26_220 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_41_267 vgnd vpwr scs8hd_decap_8
XANTENNA__42__A _42_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_22.mux_l1_in_0_ right_top_grid_pin_49_ chany_top_in[10] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_6.mux_l2_in_1__S mux_right_track_6.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_60_ chanx_right_in[16] chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_32_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 _27_/HI vgnd vpwr scs8hd_diode_2
XFILLER_23_234 vgnd vpwr scs8hd_decap_3
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.scs8hd_buf_4_0__A mux_right_track_6.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_245 vgnd vpwr scs8hd_decap_8
XANTENNA__37__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
X_43_ _43_/A chanx_right_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_259 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D mux_right_track_26.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_26_ _26_/HI _26_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_101 vpwr vgnd scs8hd_fill_2
XFILLER_37_145 vpwr vgnd scs8hd_fill_2
XFILLER_28_123 vgnd vpwr scs8hd_decap_12
XANTENNA__50__A _50_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_126 vgnd vpwr scs8hd_decap_12
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 _32_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_126 vgnd vpwr scs8hd_decap_12
XFILLER_15_27 vgnd vpwr scs8hd_decap_4
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_107 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XFILLER_16_159 vgnd vpwr scs8hd_decap_12
XANTENNA__45__A _45_/A vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_129 vgnd vpwr scs8hd_decap_8
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_59 vpwr vgnd scs8hd_fill_2
XFILLER_21_140 vpwr vgnd scs8hd_fill_2
XFILLER_13_129 vgnd vpwr scs8hd_decap_12
XFILLER_21_173 vpwr vgnd scs8hd_fill_2
XFILLER_29_240 vpwr vgnd scs8hd_fill_2
XFILLER_12_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_35_210 vpwr vgnd scs8hd_fill_2
XFILLER_35_276 vgnd vpwr scs8hd_fill_1
XFILLER_12_39 vgnd vpwr scs8hd_decap_12
XFILLER_41_202 vgnd vpwr scs8hd_decap_12
XFILLER_26_254 vpwr vgnd scs8hd_fill_2
XFILLER_26_232 vgnd vpwr scs8hd_fill_1
XFILLER_32_268 vgnd vpwr scs8hd_decap_8
XFILLER_27_80 vgnd vpwr scs8hd_decap_12
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
Xmux_right_track_4.scs8hd_buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _53_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_4_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vgnd vpwr scs8hd_decap_4
XANTENNA__53__A _53_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_183 vgnd vpwr scs8hd_decap_12
X_42_ _42_/A chanx_right_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_227 vgnd vpwr scs8hd_decap_12
XANTENNA__48__A _48_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_271 vgnd vpwr scs8hd_decap_6
XFILLER_6_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_124 vpwr vgnd scs8hd_fill_2
X_25_ _25_/HI _25_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XFILLER_34_138 vgnd vpwr scs8hd_decap_4
XFILLER_35_80 vgnd vpwr scs8hd_decap_12
XFILLER_25_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_33_160 vpwr vgnd scs8hd_fill_2
XFILLER_40_119 vgnd vpwr scs8hd_decap_3
XFILLER_25_149 vpwr vgnd scs8hd_fill_2
XFILLER_25_138 vpwr vgnd scs8hd_fill_2
XFILLER_31_27 vgnd vpwr scs8hd_decap_4
Xmem_right_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_16.mux_l1_in_0_/S mux_right_track_16.mux_l2_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__61__A chanx_right_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_21_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_163 vgnd vpwr scs8hd_decap_8
XFILLER_26_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 _20_/HI vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA__56__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_196 vgnd vpwr scs8hd_decap_12
XFILLER_8_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_266 vgnd vpwr scs8hd_decap_8
XFILLER_26_200 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.scs8hd_buf_4_0__A mux_top_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_18.scs8hd_buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _46_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_32_214 vgnd vpwr scs8hd_fill_1
XFILLER_32_236 vgnd vpwr scs8hd_decap_8
XFILLER_4_74 vgnd vpwr scs8hd_decap_12
XFILLER_23_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 _22_/HI vgnd vpwr scs8hd_diode_2
X_41_ chany_top_in[13] chanx_right_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_1_195 vgnd vpwr scs8hd_decap_12
XFILLER_1_162 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_4
XFILLER_18_39 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_12
XFILLER_11_239 vgnd vpwr scs8hd_decap_12
XANTENNA__64__A chanx_right_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_6_232 vgnd vpwr scs8hd_decap_12
X_24_ _24_/HI _24_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_158 vgnd vpwr scs8hd_fill_1
XFILLER_29_27 vgnd vpwr scs8hd_decap_4
XFILLER_10_62 vgnd vpwr scs8hd_decap_12
XFILLER_10_51 vgnd vpwr scs8hd_decap_8
XFILLER_3_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_125 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D mux_top_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__59__A chanx_right_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
XFILLER_19_93 vgnd vpwr scs8hd_decap_12
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_117 vpwr vgnd scs8hd_fill_2
XFILLER_33_183 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_14.mux_l2_in_0_/S mux_right_track_16.mux_l1_in_0_/S
+ mem_right_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_6
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_172 vgnd vpwr scs8hd_fill_1
XFILLER_24_150 vgnd vpwr scs8hd_decap_4
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[19] vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_175 vgnd vpwr scs8hd_decap_4
XFILLER_38_220 vgnd vpwr scs8hd_decap_6
XFILLER_38_264 vgnd vpwr scs8hd_decap_12
XFILLER_26_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_26.scs8hd_buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _42_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA__72__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_35_234 vgnd vpwr scs8hd_decap_6
XFILLER_35_245 vpwr vgnd scs8hd_fill_2
XFILLER_35_256 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_190 vgnd vpwr scs8hd_decap_8
XFILLER_37_27 vgnd vpwr scs8hd_decap_4
XFILLER_41_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_105 vgnd vpwr scs8hd_decap_12
XANTENNA__67__A chanx_right_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_32_204 vpwr vgnd scs8hd_fill_2
XFILLER_27_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D mux_top_track_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_171 vgnd vpwr scs8hd_decap_12
XFILLER_4_86 vgnd vpwr scs8hd_decap_12
XFILLER_23_259 vgnd vpwr scs8hd_decap_3
XFILLER_23_226 vgnd vpwr scs8hd_decap_8
XFILLER_23_215 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.scs8hd_buf_4_0_ mux_top_track_8.mux_l2_in_0_/X _71_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
X_40_ chany_top_in[14] chanx_right_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_1_141 vgnd vpwr scs8hd_decap_12
XFILLER_20_218 vgnd vpwr scs8hd_decap_8
XFILLER_13_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D mux_right_track_8.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
X_23_ _23_/HI _23_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_74 vgnd vpwr scs8hd_decap_12
XANTENNA__75__A _75_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_192 vgnd vpwr scs8hd_decap_3
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_184 vgnd vpwr scs8hd_decap_12
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_232 vgnd vpwr scs8hd_fill_1
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_276 vgnd vpwr scs8hd_fill_1
XFILLER_29_265 vpwr vgnd scs8hd_fill_2
XFILLER_16_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_110 vgnd vpwr scs8hd_decap_12
XFILLER_8_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.scs8hd_buf_4_0__A mux_top_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_224 vpwr vgnd scs8hd_fill_2
XFILLER_41_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_117 vgnd vpwr scs8hd_decap_12
XFILLER_17_235 vgnd vpwr scs8hd_decap_8
XFILLER_40_271 vgnd vpwr scs8hd_decap_6
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_98 vgnd vpwr scs8hd_decap_12
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
Xmem_right_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_10.scs8hd_buf_4_0__A mux_right_track_10.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_190 vgnd vpwr scs8hd_fill_1
XFILLER_24_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_1_ _34_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_62 vgnd vpwr scs8hd_decap_12
XFILLER_6_245 vgnd vpwr scs8hd_decap_12
X_22_ _22_/HI _22_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_149 vpwr vgnd scs8hd_fill_2
XFILLER_1_44 vgnd vpwr scs8hd_decap_12
XFILLER_28_138 vgnd vpwr scs8hd_decap_3
XFILLER_10_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_259 vpwr vgnd scs8hd_fill_2
XFILLER_3_215 vgnd vpwr scs8hd_decap_12
XFILLER_19_138 vgnd vpwr scs8hd_decap_12
XFILLER_19_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_1_ right_top_grid_pin_48_ mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_141 vgnd vpwr scs8hd_decap_12
XFILLER_30_111 vpwr vgnd scs8hd_fill_2
XFILLER_30_144 vgnd vpwr scs8hd_fill_1
XFILLER_30_199 vgnd vpwr scs8hd_decap_8
XFILLER_7_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_144 vpwr vgnd scs8hd_fill_2
XFILLER_21_177 vpwr vgnd scs8hd_fill_2
XFILLER_29_244 vpwr vgnd scs8hd_fill_2
XFILLER_32_51 vgnd vpwr scs8hd_decap_8
XFILLER_32_62 vgnd vpwr scs8hd_decap_12
XFILLER_16_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_159 vgnd vpwr scs8hd_decap_12
XFILLER_26_258 vpwr vgnd scs8hd_fill_2
XFILLER_26_236 vgnd vpwr scs8hd_decap_3
XFILLER_41_239 vgnd vpwr scs8hd_fill_1
XFILLER_5_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_247 vpwr vgnd scs8hd_fill_2
Xmem_right_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_24.mux_l1_in_0_/S mux_right_track_24.mux_l2_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_184 vgnd vpwr scs8hd_decap_12
Xmem_top_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_239 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l1_in_0__S mux_right_track_20.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_154 vgnd vpwr scs8hd_decap_8
XFILLER_13_250 vpwr vgnd scs8hd_fill_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
XFILLER_9_254 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_24.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_1_/S
+ mem_right_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_16.mux_l2_in_0_ _27_/HI mux_right_track_16.mux_l1_in_0_/X mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D mux_right_track_14.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_40_62 vgnd vpwr scs8hd_decap_12
XFILLER_40_51 vgnd vpwr scs8hd_decap_8
XFILLER_10_253 vpwr vgnd scs8hd_fill_2
XFILLER_10_220 vgnd vpwr scs8hd_decap_12
XFILLER_6_257 vgnd vpwr scs8hd_decap_12
X_21_ _21_/HI _21_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_128 vpwr vgnd scs8hd_fill_2
XFILLER_1_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_106 vpwr vgnd scs8hd_fill_2
XFILLER_3_227 vgnd vpwr scs8hd_decap_12
XFILLER_10_98 vgnd vpwr scs8hd_decap_12
XFILLER_19_117 vgnd vpwr scs8hd_decap_8
XFILLER_33_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_ right_top_grid_pin_46_ right_top_grid_pin_44_ mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_175 vgnd vpwr scs8hd_decap_8
XFILLER_24_142 vgnd vpwr scs8hd_decap_4
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_123 vgnd vpwr scs8hd_decap_3
XFILLER_7_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
XFILLER_29_223 vpwr vgnd scs8hd_fill_2
XFILLER_29_212 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vgnd vpwr scs8hd_decap_12
XFILLER_32_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__S mux_right_track_12.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D mux_right_track_14.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_240 vpwr vgnd scs8hd_fill_2
XFILLER_25_270 vgnd vpwr scs8hd_decap_4
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
Xmem_right_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_22.mux_l2_in_0_/S mux_right_track_24.mux_l1_in_0_/S
+ mem_right_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_4_196 vgnd vpwr scs8hd_decap_12
Xmem_top_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_0.mux_l2_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_31_240 vpwr vgnd scs8hd_fill_2
XFILLER_13_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_51 vgnd vpwr scs8hd_decap_8
XFILLER_38_62 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_8.mux_l1_in_1_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_18.scs8hd_buf_4_0__A mux_right_track_18.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_86 vgnd vpwr scs8hd_decap_12
XFILLER_10_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_74 vgnd vpwr scs8hd_decap_12
XFILLER_6_269 vgnd vpwr scs8hd_decap_8
X_20_ _20_/HI _20_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_1_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D mux_top_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_173 vpwr vgnd scs8hd_fill_2
XFILLER_3_239 vgnd vpwr scs8hd_decap_12
XFILLER_35_96 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_0_ right_top_grid_pin_46_ chany_top_in[7] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_154 vgnd vpwr scs8hd_decap_4
XFILLER_33_187 vpwr vgnd scs8hd_fill_2
XFILLER_18_195 vgnd vpwr scs8hd_decap_4
XFILLER_18_184 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[1] mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_110 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_32 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_154 vgnd vpwr scs8hd_decap_12
XFILLER_7_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_29_257 vpwr vgnd scs8hd_fill_2
XFILLER_16_98 vgnd vpwr scs8hd_decap_12
XFILLER_12_135 vgnd vpwr scs8hd_decap_12
XFILLER_32_86 vgnd vpwr scs8hd_decap_12
XFILLER_35_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_17_227 vgnd vpwr scs8hd_decap_6
XFILLER_32_208 vgnd vpwr scs8hd_decap_6
XFILLER_16_271 vgnd vpwr scs8hd_decap_6
XFILLER_14_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_44 vgnd vpwr scs8hd_decap_12
XFILLER_1_167 vpwr vgnd scs8hd_fill_2
XFILLER_38_74 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_1_/S
+ mem_right_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 _34_/HI vgnd vpwr scs8hd_diode_2
XFILLER_39_193 vpwr vgnd scs8hd_fill_2
XFILLER_24_98 vgnd vpwr scs8hd_decap_12
XFILLER_40_86 vgnd vpwr scs8hd_decap_12
XFILLER_36_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_32 vgnd vpwr scs8hd_decap_12
XFILLER_27_163 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_44 vgnd vpwr scs8hd_decap_12
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_30_147 vgnd vpwr scs8hd_decap_3
XFILLER_15_166 vgnd vpwr scs8hd_decap_12
XFILLER_7_68 vgnd vpwr scs8hd_decap_12
XFILLER_38_236 vgnd vpwr scs8hd_decap_6
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_6
XFILLER_12_147 vgnd vpwr scs8hd_decap_12
XFILLER_32_98 vgnd vpwr scs8hd_decap_6
XFILLER_20_191 vpwr vgnd scs8hd_fill_2
XFILLER_35_206 vpwr vgnd scs8hd_fill_2
XFILLER_26_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_261 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_27_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_110 vgnd vpwr scs8hd_decap_12
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D mux_top_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_264 vgnd vpwr scs8hd_decap_12
XFILLER_22_231 vpwr vgnd scs8hd_fill_2
XFILLER_13_56 vgnd vpwr scs8hd_decap_12
XFILLER_38_86 vgnd vpwr scs8hd_decap_12
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_224 vgnd vpwr scs8hd_decap_12
XFILLER_9_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_10_245 vgnd vpwr scs8hd_decap_8
XFILLER_40_98 vgnd vpwr scs8hd_decap_8
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_44 vgnd vpwr scs8hd_decap_12
XFILLER_19_11 vgnd vpwr scs8hd_decap_12
XFILLER_35_32 vgnd vpwr scs8hd_decap_12
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_145 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.scs8hd_buf_4_0__A mux_right_track_4.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 _25_/HI vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_30_104 vgnd vpwr scs8hd_fill_1
XFILLER_30_115 vgnd vpwr scs8hd_decap_6
XFILLER_30_159 vpwr vgnd scs8hd_fill_2
XFILLER_15_178 vgnd vpwr scs8hd_decap_12
XFILLER_21_148 vgnd vpwr scs8hd_decap_3
XFILLER_29_215 vpwr vgnd scs8hd_fill_2
XFILLER_12_159 vgnd vpwr scs8hd_decap_12
XFILLER_7_141 vgnd vpwr scs8hd_decap_12
XFILLER_34_251 vgnd vpwr scs8hd_fill_1
XFILLER_27_44 vgnd vpwr scs8hd_decap_12
XFILLER_25_262 vpwr vgnd scs8hd_fill_2
XFILLER_40_232 vgnd vpwr scs8hd_decap_8
XFILLER_4_59 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_210 vpwr vgnd scs8hd_fill_2
XFILLER_31_265 vpwr vgnd scs8hd_fill_2
XFILLER_31_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_68 vgnd vpwr scs8hd_decap_12
XFILLER_38_98 vgnd vpwr scs8hd_decap_6
XFILLER_13_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1__S mux_right_track_6.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_269 vgnd vpwr scs8hd_decap_6
XFILLER_9_236 vgnd vpwr scs8hd_decap_12
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_5_80 vgnd vpwr scs8hd_decap_12
XFILLER_39_162 vgnd vpwr scs8hd_decap_3
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 _18_/HI vgnd vpwr scs8hd_diode_2
XFILLER_36_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D mux_right_track_2.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_20.mux_l2_in_0__A0 _30_/HI vgnd vpwr scs8hd_diode_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vgnd vpwr scs8hd_decap_12
XFILLER_19_23 vgnd vpwr scs8hd_decap_8
XFILLER_35_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_2_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_4
XFILLER_18_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.scs8hd_buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _55_/A vgnd vpwr
+ scs8hd_buf_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_168 vgnd vpwr scs8hd_decap_4
XFILLER_24_146 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_26.scs8hd_buf_4_0__A mux_right_track_26.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__A1 mux_right_track_12.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_138 vgnd vpwr scs8hd_decap_6
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_105 vgnd vpwr scs8hd_decap_8
XFILLER_29_227 vpwr vgnd scs8hd_fill_2
XFILLER_29_205 vgnd vpwr scs8hd_fill_1
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_230 vgnd vpwr scs8hd_decap_12
XFILLER_17_208 vgnd vpwr scs8hd_decap_6
XFILLER_27_56 vgnd vpwr scs8hd_decap_12
XFILLER_25_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_123 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D mux_right_track_4.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_right_track_14.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_14.mux_l1_in_0_/S mux_right_track_14.mux_l2_in_0_/S
+ mem_right_track_14.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_9_248 vgnd vpwr scs8hd_decap_6
XFILLER_9_215 vgnd vpwr scs8hd_fill_1
XFILLER_5_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_36_155 vgnd vpwr scs8hd_decap_8
XFILLER_36_177 vgnd vpwr scs8hd_decap_6
XFILLER_36_199 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_20.mux_l2_in_0__A1 mux_right_track_20.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D mux_right_track_22.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_59 vpwr vgnd scs8hd_fill_2
XFILLER_35_56 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_19_68 vgnd vpwr scs8hd_decap_12
XFILLER_2_232 vgnd vpwr scs8hd_decap_12
XFILLER_33_103 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.scs8hd_buf_4_0_ mux_right_track_14.mux_l2_in_0_/X _48_/A vgnd
+ vpwr scs8hd_buf_1
X_59_ chanx_right_in[17] chany_top_out[16] vgnd vpwr scs8hd_buf_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_128 vgnd vpwr scs8hd_decap_8
XFILLER_23_191 vgnd vpwr scs8hd_decap_4
XFILLER_23_180 vgnd vpwr scs8hd_decap_4
XFILLER_7_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 _21_/HI vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_228 vgnd vpwr scs8hd_decap_4
XFILLER_21_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D mux_right_track_4.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_7_198 vgnd vpwr scs8hd_fill_1
XFILLER_7_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_242 vpwr vgnd scs8hd_fill_2
XFILLER_27_68 vgnd vpwr scs8hd_decap_12
XFILLER_40_245 vpwr vgnd scs8hd_fill_2
XFILLER_4_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_1_ _23_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_253 vpwr vgnd scs8hd_fill_2
XFILLER_16_220 vgnd vpwr scs8hd_decap_12
XFILLER_31_234 vgnd vpwr scs8hd_decap_4
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_190 vgnd vpwr scs8hd_decap_12
Xmem_right_track_14.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_12.mux_l2_in_0_/S mux_right_track_14.mux_l1_in_0_/S
+ mem_right_track_14.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D mux_right_track_22.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_105 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vgnd vpwr scs8hd_fill_1
XFILLER_5_93 vgnd vpwr scs8hd_decap_12
XFILLER_39_186 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_ right_bottom_grid_pin_1_ right_top_grid_pin_48_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XFILLER_6_208 vgnd vpwr scs8hd_decap_12
Xmux_right_track_22.scs8hd_buf_4_0_ mux_right_track_22.mux_l2_in_0_/X _44_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_5_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_75_ _75_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_36_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_167 vgnd vpwr scs8hd_decap_3
Xmux_top_track_24.mux_l2_in_0_ _20_/HI mux_top_track_24.mux_l1_in_0_/X mux_top_track_24.mux_l2_in_0_/S
+ mux_top_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_27 vgnd vpwr scs8hd_decap_12
XFILLER_35_68 vgnd vpwr scs8hd_decap_12
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_167 vgnd vpwr scs8hd_decap_4
XFILLER_27_145 vpwr vgnd scs8hd_fill_2
XANTENNA__40__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_18_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_58_ chanx_right_in[18] chany_top_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_24_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_21_15 vgnd vpwr scs8hd_decap_12
XFILLER_30_107 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.scs8hd_buf_4_0_ mux_top_track_4.mux_l2_in_0_/X _73_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_59 vpwr vgnd scs8hd_fill_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_20_195 vgnd vpwr scs8hd_decap_4
XFILLER_7_166 vgnd vpwr scs8hd_decap_12
XFILLER_34_210 vgnd vpwr scs8hd_decap_4
XFILLER_34_265 vgnd vpwr scs8hd_decap_12
XFILLER_19_251 vpwr vgnd scs8hd_fill_2
XFILLER_25_210 vpwr vgnd scs8hd_fill_2
Xmux_right_track_12.mux_l2_in_0_ _25_/HI mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_147 vgnd vpwr scs8hd_decap_12
XFILLER_17_80 vgnd vpwr scs8hd_decap_12
XFILLER_16_232 vgnd vpwr scs8hd_decap_12
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_213 vgnd vpwr scs8hd_decap_3
XFILLER_13_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_117 vgnd vpwr scs8hd_decap_12
XFILLER_13_202 vgnd vpwr scs8hd_decap_12
XANTENNA__43__A _43_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_121 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_ right_top_grid_pin_46_ right_top_grid_pin_44_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__38__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
X_74_ chanx_right_in[2] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_36_102 vgnd vpwr scs8hd_fill_1
XFILLER_36_135 vgnd vpwr scs8hd_fill_1
XFILLER_10_39 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_18_135 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_149 vpwr vgnd scs8hd_fill_2
XFILLER_25_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_62 vgnd vpwr scs8hd_decap_12
XFILLER_2_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[11] vgnd vpwr scs8hd_diode_2
X_57_ chanx_right_in[19] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_32_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_105 vgnd vpwr scs8hd_decap_12
XFILLER_23_171 vpwr vgnd scs8hd_fill_2
XFILLER_11_93 vgnd vpwr scs8hd_decap_12
XANTENNA__51__A _51_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_1_ mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_14_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_22.mux_l2_in_0__S mux_right_track_22.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_219 vpwr vgnd scs8hd_fill_2
XFILLER_29_208 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_12
XFILLER_32_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_241 vgnd vpwr scs8hd_decap_3
XANTENNA__46__A _46_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_141 vgnd vpwr scs8hd_decap_12
XFILLER_7_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_222 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_25_266 vpwr vgnd scs8hd_fill_2
XFILLER_25_200 vgnd vpwr scs8hd_fill_1
XFILLER_4_159 vgnd vpwr scs8hd_decap_12
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_6
XFILLER_33_80 vgnd vpwr scs8hd_decap_12
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_236 vgnd vpwr scs8hd_decap_8
XFILLER_22_225 vgnd vpwr scs8hd_decap_4
XFILLER_1_129 vgnd vpwr scs8hd_decap_12
XFILLER_13_258 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_ right_top_grid_pin_44_ chany_top_in[5] mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_133 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[19] mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_59 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__54__A _54_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_276 vgnd vpwr scs8hd_fill_1
X_73_ _73_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_36_114 vgnd vpwr scs8hd_decap_8
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_2_257 vgnd vpwr scs8hd_decap_12
XANTENNA__49__A _49_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
Xmem_right_track_22.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_22.mux_l1_in_0_/S mux_right_track_22.mux_l2_in_0_/S
+ mem_right_track_22.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_139 vgnd vpwr scs8hd_fill_1
XFILLER_18_147 vgnd vpwr scs8hd_decap_12
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_80 vgnd vpwr scs8hd_decap_12
X_56_ chanx_right_in[0] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_2_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_24.mux_l1_in_1_ _32_/HI right_bottom_grid_pin_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_172 vgnd vpwr scs8hd_decap_4
XFILLER_15_117 vgnd vpwr scs8hd_decap_12
Xmem_right_track_6.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l3_in_0_/S
+ mem_right_track_6.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A0 _28_/HI vgnd vpwr scs8hd_diode_2
X_39_ chany_top_in[15] chanx_right_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_16_39 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_12
XFILLER_20_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__62__A chanx_right_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_19_242 vgnd vpwr scs8hd_fill_1
XFILLER_34_245 vgnd vpwr scs8hd_decap_6
XFILLER_8_51 vgnd vpwr scs8hd_decap_8
XFILLER_8_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XANTENNA__57__A chanx_right_in[19] vgnd vpwr scs8hd_diode_2
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_93 vgnd vpwr scs8hd_decap_12
XFILLER_16_245 vgnd vpwr scs8hd_decap_8
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_59 vpwr vgnd scs8hd_fill_2
XFILLER_13_215 vgnd vpwr scs8hd_decap_12
XFILLER_39_101 vgnd vpwr scs8hd_decap_4
XFILLER_39_145 vpwr vgnd scs8hd_fill_2
XFILLER_24_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_12
XANTENNA__70__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
X_72_ chanx_right_in[4] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_39_80 vgnd vpwr scs8hd_decap_12
XFILLER_35_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
Xmem_right_track_22.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_20.mux_l2_in_0_/S mux_right_track_22.mux_l1_in_0_/S
+ mem_right_track_22.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_26.mux_l2_in_0__A0 _33_/HI vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_33_107 vgnd vpwr scs8hd_decap_3
XFILLER_18_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l3_in_0__S mux_right_track_6.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__65__A chanx_right_in[11] vgnd vpwr scs8hd_diode_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_93 vgnd vpwr scs8hd_decap_12
X_55_ _55_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_86 vgnd vpwr scs8hd_decap_12
Xmux_right_track_24.mux_l1_in_0_ right_top_grid_pin_42_ chany_top_in[11] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_129 vgnd vpwr scs8hd_decap_12
XFILLER_23_195 vgnd vpwr scs8hd_fill_1
Xmem_right_track_6.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l2_in_0_/S
+ mem_right_track_6.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_6.scs8hd_buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _52_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_14_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l2_in_0__A1 mux_right_track_18.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.scs8hd_buf_4_0__A mux_right_track_16.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
X_38_ chany_top_in[16] chanx_right_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_37_210 vgnd vpwr scs8hd_decap_4
XFILLER_37_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_39 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vpwr vgnd scs8hd_fill_2
XFILLER_20_165 vgnd vpwr scs8hd_decap_12
XFILLER_20_110 vgnd vpwr scs8hd_decap_12
XFILLER_11_154 vgnd vpwr scs8hd_decap_12
XFILLER_19_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_74 vgnd vpwr scs8hd_decap_12
XFILLER_40_249 vgnd vpwr scs8hd_fill_1
XFILLER_25_224 vpwr vgnd scs8hd_fill_2
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_93 vgnd vpwr scs8hd_decap_4
XANTENNA__73__A _73_/A vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_0__S mux_right_track_12.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_27 vgnd vpwr scs8hd_decap_12
XFILLER_21_260 vpwr vgnd scs8hd_fill_2
XFILLER_13_227 vgnd vpwr scs8hd_decap_12
XANTENNA__68__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_39_113 vpwr vgnd scs8hd_fill_2
XFILLER_10_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_14_62 vgnd vpwr scs8hd_decap_12
XFILLER_14_51 vgnd vpwr scs8hd_decap_8
X_71_ _71_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_27_149 vpwr vgnd scs8hd_fill_2
XFILLER_27_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D mux_right_track_10.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_26.mux_l2_in_0__A1 mux_right_track_26.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_141 vgnd vpwr scs8hd_decap_12
XFILLER_26_160 vpwr vgnd scs8hd_fill_2
XFILLER_41_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 right_bottom_grid_pin_1_ vgnd vpwr scs8hd_diode_2
X_54_ _54_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_98 vgnd vpwr scs8hd_decap_12
XFILLER_32_141 vgnd vpwr scs8hd_decap_4
XFILLER_23_163 vgnd vpwr scs8hd_decap_8
Xmem_right_track_6.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_1_/S
+ mem_right_track_6.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_200 vgnd vpwr scs8hd_fill_1
XFILLER_37_222 vpwr vgnd scs8hd_fill_2
X_37_ chany_top_in[17] chanx_right_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_20_177 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_233 vpwr vgnd scs8hd_fill_2
XFILLER_28_200 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _23_/HI vgnd vpwr scs8hd_diode_2
XFILLER_22_62 vgnd vpwr scs8hd_decap_12
XFILLER_22_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_211 vgnd vpwr scs8hd_fill_1
XFILLER_34_214 vgnd vpwr scs8hd_fill_1
XFILLER_8_86 vgnd vpwr scs8hd_decap_12
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XFILLER_25_236 vgnd vpwr scs8hd_fill_1
XFILLER_31_206 vpwr vgnd scs8hd_fill_2
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_286 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_39 vgnd vpwr scs8hd_decap_12
XFILLER_21_272 vgnd vpwr scs8hd_decap_3
XFILLER_13_239 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D mux_right_track_10.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_125 vpwr vgnd scs8hd_fill_2
XFILLER_5_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_74 vgnd vpwr scs8hd_decap_12
XFILLER_5_202 vgnd vpwr scs8hd_decap_12
XFILLER_30_62 vgnd vpwr scs8hd_decap_12
XFILLER_30_51 vgnd vpwr scs8hd_decap_8
X_70_ chanx_right_in[6] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_12
XFILLER_35_183 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_172 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
X_53_ _53_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D mux_top_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_164 vpwr vgnd scs8hd_fill_2
XFILLER_32_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_36_ chany_top_in[18] chanx_right_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_37_245 vpwr vgnd scs8hd_fill_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_123 vgnd vpwr scs8hd_decap_4
XFILLER_9_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_245 vgnd vpwr scs8hd_decap_3
XFILLER_28_212 vgnd vpwr scs8hd_decap_3
XFILLER_11_178 vgnd vpwr scs8hd_decap_12
XFILLER_7_105 vgnd vpwr scs8hd_decap_12
XFILLER_22_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_34_226 vpwr vgnd scs8hd_fill_2
XFILLER_8_98 vgnd vpwr scs8hd_decap_12
XFILLER_6_171 vgnd vpwr scs8hd_decap_12
X_19_ _19_/HI _19_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_270 vgnd vpwr scs8hd_decap_4
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_141 vgnd vpwr scs8hd_decap_12
XFILLER_30_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.scs8hd_buf_4_0__A mux_right_track_2.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_62 vgnd vpwr scs8hd_decap_12
XFILLER_28_51 vgnd vpwr scs8hd_decap_8
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_5_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_137 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_74 vgnd vpwr scs8hd_decap_12
XFILLER_14_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_129 vgnd vpwr scs8hd_fill_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_154 vgnd vpwr scs8hd_decap_12
XFILLER_26_184 vgnd vpwr scs8hd_decap_12
X_52_ _52_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_32_176 vgnd vpwr scs8hd_fill_1
XFILLER_23_198 vpwr vgnd scs8hd_fill_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_23_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.scs8hd_buf_4_0__A mux_top_track_24.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_32 vgnd vpwr scs8hd_decap_12
XFILLER_36_51 vgnd vpwr scs8hd_decap_8
XFILLER_36_62 vgnd vpwr scs8hd_decap_12
XFILLER_14_110 vgnd vpwr scs8hd_decap_12
X_35_ _35_/HI _35_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_117 vgnd vpwr scs8hd_decap_12
XFILLER_22_86 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
X_18_ _18_/HI _18_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_274 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.scs8hd_buf_4_0__A mux_right_track_24.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_252 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D mux_right_track_16.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_74 vgnd vpwr scs8hd_decap_12
XFILLER_8_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_193 vgnd vpwr scs8hd_decap_4
XFILLER_30_86 vgnd vpwr scs8hd_decap_12
XFILLER_14_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_259 vpwr vgnd scs8hd_fill_2
XFILLER_5_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_35_174 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
XFILLER_26_196 vgnd vpwr scs8hd_decap_4
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_166 vgnd vpwr scs8hd_decap_12
XFILLER_1_251 vgnd vpwr scs8hd_decap_4
X_51_ _51_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_17_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D mux_top_track_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_12.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_12.mux_l1_in_0_/S mux_right_track_12.mux_l2_in_0_/S
+ mem_right_track_12.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_24.scs8hd_buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _63_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_11_44 vgnd vpwr scs8hd_decap_12
XFILLER_36_74 vgnd vpwr scs8hd_decap_12
X_34_ _34_/HI _34_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_269 vgnd vpwr scs8hd_decap_8
XFILLER_22_98 vgnd vpwr scs8hd_decap_12
XFILLER_7_129 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D mux_right_track_16.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_217 vgnd vpwr scs8hd_decap_3
XFILLER_19_247 vpwr vgnd scs8hd_fill_2
XFILLER_19_203 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_6_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_1_ _35_/HI right_top_grid_pin_49_ mux_right_track_6.mux_l2_in_0_/S
+ mux_right_track_6.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_228 vgnd vpwr scs8hd_decap_8
XFILLER_25_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_17_32 vgnd vpwr scs8hd_decap_12
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_264 vgnd vpwr scs8hd_decap_8
Xmux_right_track_10.scs8hd_buf_4_0_ mux_right_track_10.mux_l2_in_0_/X _50_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_28_86 vgnd vpwr scs8hd_decap_12
XFILLER_12_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_257 vgnd vpwr scs8hd_decap_12
XFILLER_8_213 vgnd vpwr scs8hd_decap_12
XFILLER_5_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 _19_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_98 vgnd vpwr scs8hd_decap_6
XFILLER_5_227 vgnd vpwr scs8hd_decap_12
XFILLER_29_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_6
XFILLER_2_208 vgnd vpwr scs8hd_decap_12
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_26_175 vgnd vpwr scs8hd_decap_8
XFILLER_26_164 vgnd vpwr scs8hd_decap_8
XFILLER_25_32 vgnd vpwr scs8hd_decap_12
XFILLER_41_178 vgnd vpwr scs8hd_decap_12
XFILLER_1_263 vgnd vpwr scs8hd_decap_12
X_50_ _50_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
Xmem_right_track_12.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_10.mux_l2_in_0_/S mux_right_track_12.mux_l1_in_0_/S
+ mem_right_track_12.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_23_145 vpwr vgnd scs8hd_fill_2
XFILLER_11_56 vgnd vpwr scs8hd_decap_12
XFILLER_36_86 vgnd vpwr scs8hd_decap_12
XFILLER_14_123 vgnd vpwr scs8hd_decap_12
X_33_ _33_/HI _33_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_26.mux_l1_in_0__S mux_right_track_26.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_259 vpwr vgnd scs8hd_fill_2
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_237 vpwr vgnd scs8hd_fill_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
Xmux_right_track_18.mux_l2_in_0_ _28_/HI mux_right_track_18.mux_l1_in_0_/X mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_18.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_196 vgnd vpwr scs8hd_decap_12
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_20.mux_l2_in_0_ _30_/HI mux_right_track_20.mux_l1_in_0_/X mux_right_track_20.mux_l2_in_0_/S
+ mux_right_track_20.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_44 vgnd vpwr scs8hd_decap_12
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_32 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_251 vpwr vgnd scs8hd_fill_2
XFILLER_30_254 vpwr vgnd scs8hd_fill_2
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_221 vpwr vgnd scs8hd_fill_2
XFILLER_21_210 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_20.mux_l1_in_0__A0 right_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_28_98 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_269 vgnd vpwr scs8hd_decap_8
XFILLER_8_225 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_1_ right_top_grid_pin_47_ right_top_grid_pin_45_ mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_0.scs8hd_buf_4_0_ mux_top_track_0.mux_l2_in_0_/X _75_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D mux_right_track_0.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_239 vgnd vpwr scs8hd_decap_12
XFILLER_39_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_26_110 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_44 vgnd vpwr scs8hd_decap_12
XFILLER_41_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_2_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l2_in_0__S mux_right_track_18.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_168 vpwr vgnd scs8hd_fill_2
XFILLER_32_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_124 vpwr vgnd scs8hd_fill_2
XFILLER_11_68 vgnd vpwr scs8hd_decap_12
XFILLER_36_98 vgnd vpwr scs8hd_decap_4
XFILLER_14_135 vgnd vpwr scs8hd_decap_12
X_32_ _32_/HI _32_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_249 vpwr vgnd scs8hd_fill_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_4
XFILLER_20_127 vgnd vpwr scs8hd_fill_1
XFILLER_13_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_80 vgnd vpwr scs8hd_decap_12
XFILLER_11_105 vgnd vpwr scs8hd_decap_12
XFILLER_19_238 vgnd vpwr scs8hd_decap_4
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_27_260 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.scs8hd_buf_4_0__A mux_top_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A0 _35_/HI vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_241 vpwr vgnd scs8hd_fill_2
XFILLER_33_274 vgnd vpwr scs8hd_fill_1
XFILLER_18_271 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D mux_right_track_0.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_56 vgnd vpwr scs8hd_decap_12
XFILLER_16_208 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_44 vgnd vpwr scs8hd_decap_12
XFILLER_33_99 vpwr vgnd scs8hd_fill_2
XFILLER_24_274 vgnd vpwr scs8hd_decap_3
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_178 vgnd vpwr scs8hd_decap_12
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
XFILLER_30_266 vgnd vpwr scs8hd_decap_8
XFILLER_21_200 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
Xmux_right_track_18.mux_l1_in_0_ right_top_grid_pin_47_ chany_top_in[8] mux_right_track_18.mux_l1_in_0_/S
+ mux_right_track_18.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_6.mux_l3_in_0__A0 mux_right_track_6.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_237 vgnd vpwr scs8hd_decap_6
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_ right_top_grid_pin_43_ chany_top_in[2] mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_8.mux_l2_in_0_ _22_/HI mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_20.mux_l1_in_0_ right_top_grid_pin_48_ chany_top_in[9] mux_right_track_20.mux_l1_in_0_/S
+ mux_right_track_20.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D mux_right_track_18.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_163 vgnd vpwr scs8hd_fill_1
XFILLER_39_32 vgnd vpwr scs8hd_decap_12
XFILLER_29_152 vgnd vpwr scs8hd_fill_1
XFILLER_35_100 vpwr vgnd scs8hd_fill_2
XFILLER_35_166 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_25_56 vgnd vpwr scs8hd_decap_12
XFILLER_41_44 vgnd vpwr scs8hd_decap_12
XFILLER_2_27 vgnd vpwr scs8hd_decap_12
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_188 vpwr vgnd scs8hd_fill_2
XFILLER_17_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_147 vgnd vpwr scs8hd_decap_12
X_31_ _31_/HI _31_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_206 vpwr vgnd scs8hd_fill_2
XFILLER_28_217 vgnd vpwr scs8hd_decap_3
XFILLER_11_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_272 vgnd vpwr scs8hd_decap_3
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_59 vpwr vgnd scs8hd_fill_2
XFILLER_6_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 right_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_22.mux_l1_in_0__S mux_right_track_22.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_231 vgnd vpwr scs8hd_decap_8
XFILLER_17_68 vgnd vpwr scs8hd_decap_12
Xmem_right_track_20.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_20.mux_l1_in_0_/S mux_right_track_20.mux_l2_in_0_/S
+ mem_right_track_20.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_33_56 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_223 vpwr vgnd scs8hd_fill_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_80 vgnd vpwr scs8hd_decap_12
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_12_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_6.mux_l3_in_0__A1 mux_right_track_6.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_5_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_109 vpwr vgnd scs8hd_fill_2
XFILLER_38_175 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D mux_right_track_4.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 _26_/HI vgnd vpwr scs8hd_diode_2
XFILLER_39_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_197 vgnd vpwr scs8hd_decap_8
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_35_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_26_123 vgnd vpwr scs8hd_decap_12
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_41_56 vgnd vpwr scs8hd_decap_12
XFILLER_25_68 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[5] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_39 vgnd vpwr scs8hd_decap_12
XFILLER_32_104 vgnd vpwr scs8hd_fill_1
XFILLER_32_126 vgnd vpwr scs8hd_decap_8
XFILLER_32_137 vpwr vgnd scs8hd_fill_2
XFILLER_17_178 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_23_137 vgnd vpwr scs8hd_decap_6
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_159 vgnd vpwr scs8hd_decap_12
X_30_ _30_/HI _30_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_218 vpwr vgnd scs8hd_fill_2
XFILLER_9_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0__S mux_right_track_14.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_229 vpwr vgnd scs8hd_fill_2
XFILLER_3_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_129 vgnd vpwr scs8hd_decap_12
XFILLER_19_207 vgnd vpwr scs8hd_decap_4
XFILLER_8_27 vgnd vpwr scs8hd_decap_12
XFILLER_10_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_254 vpwr vgnd scs8hd_fill_2
XFILLER_33_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D mux_right_track_6.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_68 vgnd vpwr scs8hd_decap_12
XFILLER_24_254 vpwr vgnd scs8hd_fill_2
Xmem_right_track_20.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_18.mux_l2_in_0_/S mux_right_track_20.mux_l1_in_0_/S
+ mem_right_track_20.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_top_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_top_track_0.mux_l1_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_22.mux_l2_in_0__A0 _31_/HI vgnd vpwr scs8hd_diode_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l2_in_0_/S
+ mem_right_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.scs8hd_buf_4_0__A mux_right_track_14.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_2.scs8hd_buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _54_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_right_track_14.mux_l2_in_0__A1 mux_right_track_14.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_56 vgnd vpwr scs8hd_decap_12
XFILLER_29_165 vpwr vgnd scs8hd_fill_2
XFILLER_4_253 vpwr vgnd scs8hd_fill_2
XFILLER_4_220 vgnd vpwr scs8hd_decap_12
XFILLER_35_135 vgnd vpwr scs8hd_fill_1
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_41_105 vgnd vpwr scs8hd_decap_12
XFILLER_26_135 vgnd vpwr scs8hd_fill_1
XFILLER_41_68 vgnd vpwr scs8hd_decap_12
XFILLER_15_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_105 vgnd vpwr scs8hd_decap_12
XFILLER_31_171 vpwr vgnd scs8hd_fill_2
XFILLER_31_193 vpwr vgnd scs8hd_fill_2
XFILLER_23_149 vpwr vgnd scs8hd_fill_2
XFILLER_11_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D mux_right_track_6.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_193 vgnd vpwr scs8hd_decap_12
XANTENNA__41__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0__S mux_right_track_6.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_274 vgnd vpwr scs8hd_decap_3
XFILLER_22_59 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA__36__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_42_244 vgnd vpwr scs8hd_decap_4
XFILLER_8_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_196 vgnd vpwr scs8hd_decap_12
XFILLER_6_123 vgnd vpwr scs8hd_decap_12
XFILLER_33_200 vpwr vgnd scs8hd_fill_2
XFILLER_33_222 vgnd vpwr scs8hd_decap_12
XFILLER_33_266 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D mux_right_track_24.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_236 vpwr vgnd scs8hd_fill_2
XFILLER_30_258 vgnd vpwr scs8hd_decap_4
XFILLER_23_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_22.mux_l2_in_0__A1 mux_right_track_22.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_225 vpwr vgnd scs8hd_fill_2
XFILLER_9_93 vgnd vpwr scs8hd_decap_12
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
Xmem_top_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_right_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_1_/S
+ mem_right_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_269 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.scs8hd_buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _47_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_7_251 vgnd vpwr scs8hd_decap_12
XFILLER_38_199 vpwr vgnd scs8hd_fill_2
XFILLER_14_27 vgnd vpwr scs8hd_decap_12
XFILLER_30_59 vpwr vgnd scs8hd_fill_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_68 vgnd vpwr scs8hd_decap_12
XFILLER_29_133 vgnd vpwr scs8hd_fill_1
XANTENNA__44__A _44_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 right_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_41_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_213 vgnd vpwr scs8hd_fill_1
XANTENNA__39__A chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_31_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_117 vgnd vpwr scs8hd_fill_1
XFILLER_9_154 vgnd vpwr scs8hd_decap_12
XFILLER_22_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_264 vgnd vpwr scs8hd_decap_8
XFILLER_6_135 vgnd vpwr scs8hd_decap_12
XANTENNA__52__A _52_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_212 vpwr vgnd scs8hd_fill_2
XFILLER_18_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_190 vgnd vpwr scs8hd_decap_12
Xmem_top_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_4.mux_l2_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.mux_l2_in_0__S mux_right_track_10.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_24.scs8hd_buf_4_0_ mux_right_track_24.mux_l2_in_0_/X _43_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA__47__A _47_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XFILLER_21_248 vpwr vgnd scs8hd_fill_2
XFILLER_21_215 vgnd vpwr scs8hd_decap_3
Xmem_top_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_8.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_208 vgnd vpwr scs8hd_fill_1
XFILLER_7_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 right_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_38_123 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_12
XFILLER_14_39 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_145 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__60__A chanx_right_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_29_80 vgnd vpwr scs8hd_decap_12
XFILLER_6_62 vgnd vpwr scs8hd_decap_12
XFILLER_6_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_27 vgnd vpwr scs8hd_decap_4
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_32_118 vgnd vpwr scs8hd_decap_4
XANTENNA__55__A _55_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_184 vgnd vpwr scs8hd_decap_12
XFILLER_40_173 vpwr vgnd scs8hd_fill_2
XFILLER_25_192 vgnd vpwr scs8hd_decap_8
XFILLER_15_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.scs8hd_buf_4_0__A mux_right_track_0.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l2_in_1_ _29_/HI right_top_grid_pin_49_ mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_59 vpwr vgnd scs8hd_fill_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_9_166 vgnd vpwr scs8hd_decap_12
XFILLER_36_243 vgnd vpwr scs8hd_fill_1
XFILLER_36_254 vgnd vpwr scs8hd_decap_8
XFILLER_22_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_210 vpwr vgnd scs8hd_fill_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
XFILLER_27_243 vpwr vgnd scs8hd_fill_2
XFILLER_10_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_147 vgnd vpwr scs8hd_decap_12
XFILLER_37_80 vgnd vpwr scs8hd_decap_12
XFILLER_18_232 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__63__A _63_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_28_27 vgnd vpwr scs8hd_decap_12
XFILLER_20_271 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D mux_top_track_8.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA__58__A chanx_right_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_38_135 vgnd vpwr scs8hd_fill_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_30_39 vgnd vpwr scs8hd_decap_12
XFILLER_39_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XFILLER_4_245 vgnd vpwr scs8hd_decap_8
XFILLER_35_138 vpwr vgnd scs8hd_fill_2
XFILLER_6_74 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_138 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_34_193 vpwr vgnd scs8hd_fill_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_17_105 vgnd vpwr scs8hd_decap_12
XFILLER_40_196 vgnd vpwr scs8hd_fill_1
XANTENNA__71__A _71_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XFILLER_31_93 vgnd vpwr scs8hd_decap_8
Xmux_right_track_14.mux_l2_in_0_ _26_/HI mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_14.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_163 vpwr vgnd scs8hd_fill_2
XFILLER_16_171 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_right_track_22.scs8hd_buf_4_0__A mux_right_track_22.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_12
XANTENNA__66__A chanx_right_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_13_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XFILLER_9_178 vgnd vpwr scs8hd_decap_12
XFILLER_36_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_62 vgnd vpwr scs8hd_decap_12
XFILLER_12_51 vgnd vpwr scs8hd_decap_8
XFILLER_6_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_ right_top_grid_pin_47_ right_top_grid_pin_45_ mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_258 vpwr vgnd scs8hd_fill_2
X_69_ chanx_right_in[7] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_258 vgnd vpwr scs8hd_decap_4
XFILLER_3_129 vgnd vpwr scs8hd_decap_12
XFILLER_2_184 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_10.mux_l1_in_0_/S mux_right_track_10.mux_l2_in_0_/S
+ mem_right_track_10.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_39 vgnd vpwr scs8hd_decap_12
XANTENNA__74__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_39_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_169 vgnd vpwr scs8hd_decap_3
XFILLER_20_62 vgnd vpwr scs8hd_decap_12
XANTENNA__69__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_93 vgnd vpwr scs8hd_decap_12
XFILLER_6_86 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_19_180 vpwr vgnd scs8hd_fill_2
XFILLER_1_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.scs8hd_buf_4_0__A mux_right_track_8.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_164 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_242 vpwr vgnd scs8hd_fill_2
XFILLER_36_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_3_32 vgnd vpwr scs8hd_decap_12
XFILLER_36_212 vgnd vpwr scs8hd_decap_8
XFILLER_27_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_123 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_ right_top_grid_pin_45_ chany_top_in[6] mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_12_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_201 vgnd vpwr scs8hd_decap_12
Xmux_right_track_2.mux_l1_in_0_ right_top_grid_pin_43_ chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_204 vpwr vgnd scs8hd_fill_2
XFILLER_33_237 vpwr vgnd scs8hd_fill_2
XFILLER_37_93 vgnd vpwr scs8hd_decap_8
XFILLER_18_245 vgnd vpwr scs8hd_decap_8
Xmux_top_track_4.mux_l2_in_0_ _21_/HI mux_top_track_4.mux_l1_in_0_/X mux_top_track_4.mux_l2_in_0_/S
+ mux_top_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_right_track_26.mux_l2_in_0_ _33_/HI mux_right_track_26.mux_l1_in_0_/X ccff_tail
+ mux_right_track_26.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
X_68_ chanx_right_in[8] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_24_215 vpwr vgnd scs8hd_fill_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XFILLER_15_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_207 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_2_196 vgnd vpwr scs8hd_decap_12
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.scs8hd_dfxbp_1_0_ prog_clk mux_right_track_8.mux_l2_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ mem_right_track_10.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_51 vgnd vpwr scs8hd_decap_8
XFILLER_11_251 vpwr vgnd scs8hd_fill_2
XFILLER_7_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_104 vgnd vpwr scs8hd_fill_1
XFILLER_38_159 vgnd vpwr scs8hd_decap_4
XFILLER_37_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D mux_right_track_12.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.scs8hd_buf_4_0_ mux_right_track_8.mux_l2_in_0_/X _51_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_20_74 vgnd vpwr scs8hd_decap_12
XFILLER_28_192 vgnd vpwr scs8hd_decap_8
XFILLER_6_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_34_151 vgnd vpwr scs8hd_decap_12
XFILLER_1_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_184 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_265 vpwr vgnd scs8hd_fill_2
XFILLER_39_210 vgnd vpwr scs8hd_decap_4
XFILLER_22_110 vgnd vpwr scs8hd_decap_12
XFILLER_26_62 vgnd vpwr scs8hd_decap_12
XFILLER_26_51 vgnd vpwr scs8hd_decap_8
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D mux_top_track_4.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_235 vgnd vpwr scs8hd_decap_8
XFILLER_3_44 vgnd vpwr scs8hd_decap_12
XFILLER_27_224 vpwr vgnd scs8hd_fill_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_12_86 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_213 vpwr vgnd scs8hd_fill_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
X_67_ chanx_right_in[9] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 right_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_30_219 vpwr vgnd scs8hd_fill_2
XFILLER_15_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D mux_right_track_12.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_18.scs8hd_dfxbp_1_1_ prog_clk mux_right_track_18.mux_l1_in_0_/S mux_right_track_18.mux_l2_in_0_/S
+ mem_right_track_18.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_14_271 vgnd vpwr scs8hd_decap_6
XFILLER_9_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_208 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_26.mux_l1_in_0_ right_top_grid_pin_43_ chany_top_in[12] mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_51 vgnd vpwr scs8hd_decap_8
XFILLER_34_62 vgnd vpwr scs8hd_decap_12
XFILLER_29_149 vgnd vpwr scs8hd_fill_1
XFILLER_29_127 vgnd vpwr scs8hd_decap_6
XFILLER_29_105 vgnd vpwr scs8hd_fill_1
XFILLER_20_86 vgnd vpwr scs8hd_decap_12
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_182 vgnd vpwr scs8hd_fill_1
XFILLER_34_163 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 _29_/HI vgnd vpwr scs8hd_diode_2
XFILLER_1_207 vgnd vpwr scs8hd_decap_6
XFILLER_40_199 vpwr vgnd scs8hd_fill_2
XFILLER_40_177 vgnd vpwr scs8hd_decap_6
XFILLER_40_111 vgnd vpwr scs8hd_decap_8
XFILLER_31_122 vpwr vgnd scs8hd_fill_2
XFILLER_16_196 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_188 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
.ends

