* NGSPICE file created from cbx_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt cbx_1__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_grid_pin_0_ bottom_grid_pin_4_ bottom_grid_pin_8_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] data_in
+ enable top_grid_pin_14_ top_grid_pin_2_ top_grid_pin_6_ vpwr vgnd
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_56 vpwr vgnd scs8hd_fill_2
XFILLER_5_354 vgnd vpwr scs8hd_decap_12
XFILLER_3_67 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _062_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_129 vgnd vpwr scs8hd_fill_1
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_2_346 vpwr vgnd scs8hd_fill_2
XFILLER_5_140 vpwr vgnd scs8hd_fill_2
XFILLER_5_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _087_/Y vgnd vpwr
+ scs8hd_diode_2
X_062_ _074_/A _074_/B _040_/X _058_/D _062_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_11 vgnd vpwr scs8hd_decap_4
XFILLER_9_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_242 vgnd vpwr scs8hd_decap_6
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
X_045_ address[0] _059_/C vgnd vpwr scs8hd_buf_1
X_114_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_19_342 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XFILLER_16_312 vgnd vpwr scs8hd_decap_12
XFILLER_16_389 vgnd vpwr scs8hd_decap_8
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XFILLER_3_260 vpwr vgnd scs8hd_fill_2
XFILLER_3_271 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _092_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XANTENNA__042__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_43 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_0_274 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__037__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_35 vpwr vgnd scs8hd_fill_2
XFILLER_5_377 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_193 vpwr vgnd scs8hd_fill_2
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_163 vpwr vgnd scs8hd_fill_2
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
XFILLER_17_281 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA__050__A _071_/A vgnd vpwr scs8hd_diode_2
X_061_ address[2] _074_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_122 vgnd vpwr scs8hd_fill_1
XFILLER_2_100 vgnd vpwr scs8hd_decap_6
XFILLER_2_199 vpwr vgnd scs8hd_fill_2
XFILLER_2_133 vgnd vpwr scs8hd_decap_3
XFILLER_0_47 vgnd vpwr scs8hd_decap_12
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XANTENNA__045__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_225 vpwr vgnd scs8hd_fill_2
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
X_113_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_044_ _046_/A _046_/B _040_/X _046_/D _044_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_269 vgnd vpwr scs8hd_decap_12
XFILLER_19_354 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_324 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_1_209 vpwr vgnd scs8hd_fill_2
XANTENNA__042__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_55 vgnd vpwr scs8hd_decap_6
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__053__A address[4] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _070_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_106 vgnd vpwr scs8hd_decap_12
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_5_367 vgnd vpwr scs8hd_decap_6
XFILLER_12_190 vgnd vpwr scs8hd_decap_12
XANTENNA__048__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_304 vpwr vgnd scs8hd_fill_2
XFILLER_10_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_315 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _088_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_293 vgnd vpwr scs8hd_decap_12
XANTENNA__050__B _058_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_decap_4
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
X_060_ address[1] _074_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_167 vpwr vgnd scs8hd_fill_2
XFILLER_0_59 vgnd vpwr scs8hd_decap_3
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_20_211 vgnd vpwr scs8hd_decap_6
XANTENNA__061__A address[2] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _046_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
X_043_ _043_/A _046_/D vgnd vpwr scs8hd_buf_1
X_112_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__056__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_218 vpwr vgnd scs8hd_fill_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
XFILLER_3_295 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_1.LATCH_0_.latch data_in _089_/A _083_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XANTENNA__042__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_306 vgnd vpwr scs8hd_decap_12
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_12_361 vgnd vpwr scs8hd_decap_12
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XFILLER_9_118 vgnd vpwr scs8hd_decap_4
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_3_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _040_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_0_.latch data_in _087_/A _079_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
XANTENNA__050__C _059_/C vgnd vpwr scs8hd_diode_2
XANTENNA__059__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_16 vgnd vpwr scs8hd_fill_1
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_47 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _090_/A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
X_042_ address[4] address[5] address[3] _081_/B _043_/A vgnd vpwr scs8hd_or4_4
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
X_111_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_12
XFILLER_6_293 vgnd vpwr scs8hd_decap_12
XFILLER_1_92 vpwr vgnd scs8hd_fill_2
XANTENNA__056__B _046_/B vgnd vpwr scs8hd_diode_2
XANTENNA__072__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_337 vgnd vpwr scs8hd_decap_12
XANTENNA__042__D _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_318 vgnd vpwr scs8hd_decap_12
XFILLER_0_266 vpwr vgnd scs8hd_fill_2
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XFILLER_8_300 vgnd vpwr scs8hd_decap_12
XFILLER_8_377 vgnd vpwr scs8hd_decap_12
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _086_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_303 vpwr vgnd scs8hd_fill_2
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XFILLER_8_163 vgnd vpwr scs8hd_decap_8
XFILLER_8_174 vgnd vpwr scs8hd_decap_12
XFILLER_2_328 vgnd vpwr scs8hd_decap_8
XANTENNA__080__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _057_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_144 vpwr vgnd scs8hd_fill_2
XFILLER_5_199 vpwr vgnd scs8hd_fill_2
XANTENNA__050__D _046_/D vgnd vpwr scs8hd_diode_2
XANTENNA__059__B _058_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_405 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
X_110_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_041_ enable _081_/B vgnd vpwr scs8hd_inv_8
XFILLER_19_379 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _092_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA__056__C _040_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_16_349 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_220 vpwr vgnd scs8hd_fill_2
XFILLER_3_231 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _044_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_278 vgnd vpwr scs8hd_fill_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_312 vgnd vpwr scs8hd_decap_12
XFILLER_8_389 vgnd vpwr scs8hd_decap_8
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _075_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _088_/A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_178 vgnd vpwr scs8hd_decap_3
XANTENNA__059__C _059_/C vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_288 vgnd vpwr scs8hd_decap_12
XFILLER_1_170 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_281 vgnd vpwr scs8hd_decap_12
XFILLER_7_229 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_12
XFILLER_1_3 vgnd vpwr scs8hd_decap_3
X_040_ _040_/A _040_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__056__D _058_/D vgnd vpwr scs8hd_diode_2
XANTENNA__072__C _074_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_287 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__083__B _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_0_202 vpwr vgnd scs8hd_fill_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_324 vgnd vpwr scs8hd_decap_12
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_71 vgnd vpwr scs8hd_decap_12
XANTENNA__078__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_132 vpwr vgnd scs8hd_fill_2
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_2_308 vgnd vpwr scs8hd_decap_4
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_61 vgnd vpwr scs8hd_decap_8
XANTENNA__059__D _058_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_7 vgnd vpwr scs8hd_fill_1
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XFILLER_0_19 vpwr vgnd scs8hd_fill_2
XFILLER_9_17 vpwr vgnd scs8hd_fill_2
XFILLER_9_293 vgnd vpwr scs8hd_decap_12
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _059_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_208 vpwr vgnd scs8hd_fill_2
XFILLER_3_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_230 vpwr vgnd scs8hd_fill_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_6_285 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_099_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__072__D _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C _081_/X vgnd vpwr scs8hd_diode_2
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_94 vgnd vpwr scs8hd_decap_4
XANTENNA__078__C _078_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_306 vgnd vpwr scs8hd_decap_12
XFILLER_4_361 vgnd vpwr scs8hd_decap_12
XFILLER_5_103 vpwr vgnd scs8hd_fill_2
XFILLER_1_353 vgnd vpwr scs8hd_decap_12
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_106 vgnd vpwr scs8hd_fill_1
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
X_098_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_96 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_3_201 vpwr vgnd scs8hd_fill_2
XFILLER_3_256 vpwr vgnd scs8hd_fill_2
XFILLER_3_267 vpwr vgnd scs8hd_fill_2
XFILLER_15_330 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XANTENNA__083__D _074_/C vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_300 vgnd vpwr scs8hd_decap_12
XFILLER_12_377 vgnd vpwr scs8hd_decap_12
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XANTENNA__078__D _078_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_318 vgnd vpwr scs8hd_decap_12
XFILLER_17_403 vgnd vpwr scs8hd_decap_4
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_112 vgnd vpwr scs8hd_decap_12
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_141 vgnd vpwr scs8hd_decap_12
XFILLER_4_373 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _091_/A mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _062_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_18 vgnd vpwr scs8hd_decap_12
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_365 vgnd vpwr scs8hd_fill_1
XFILLER_1_332 vgnd vpwr scs8hd_decap_4
XFILLER_1_321 vpwr vgnd scs8hd_fill_2
XFILLER_5_159 vpwr vgnd scs8hd_fill_2
XFILLER_4_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_129 vpwr vgnd scs8hd_fill_2
XFILLER_2_118 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _068_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_306 vgnd vpwr scs8hd_decap_12
X_097_ _097_/HI _097_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_243 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vgnd vpwr scs8hd_decap_6
XFILLER_18_361 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _094_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _050_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XFILLER_3_235 vpwr vgnd scs8hd_fill_2
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_342 vgnd vpwr scs8hd_decap_12
XFILLER_15_375 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_312 vgnd vpwr scs8hd_decap_12
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _044_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XFILLER_12_389 vgnd vpwr scs8hd_decap_8
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_124 vgnd vpwr scs8hd_fill_1
XFILLER_4_385 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_1_.latch data_in _088_/A _082_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_300 vgnd vpwr scs8hd_decap_3
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_160 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_281 vgnd vpwr scs8hd_decap_12
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_19_318 vgnd vpwr scs8hd_decap_12
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_096_ _096_/HI _096_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_266 vgnd vpwr scs8hd_decap_8
XFILLER_18_373 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_1_.latch data_in _086_/A _078_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_10_52 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _089_/A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_354 vgnd vpwr scs8hd_decap_12
XFILLER_15_387 vgnd vpwr scs8hd_decap_12
X_079_ _075_/X address[5] _078_/C _074_/C _079_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_15_19 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_324 vgnd vpwr scs8hd_decap_12
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_191 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _097_/HI _090_/Y mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_231 vgnd vpwr scs8hd_decap_12
XFILLER_13_293 vgnd vpwr scs8hd_decap_12
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XFILLER_1_8 vgnd vpwr scs8hd_decap_3
X_095_ _095_/HI _095_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
XFILLER_6_289 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_385 vgnd vpwr scs8hd_decap_12
XFILLER_10_64 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_399 vgnd vpwr scs8hd_decap_8
X_078_ _075_/X address[5] _078_/C _078_/D _078_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__106__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_218 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_43 vpwr vgnd scs8hd_fill_2
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_166 vgnd vpwr scs8hd_decap_12
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XFILLER_4_140 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_31 vgnd vpwr scs8hd_decap_12
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_176 vpwr vgnd scs8hd_fill_2
XFILLER_1_132 vgnd vpwr scs8hd_decap_4
XANTENNA__109__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
X_094_ _094_/HI _094_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vpwr vgnd scs8hd_fill_2
XFILLER_1_45 vpwr vgnd scs8hd_fill_2
XFILLER_1_67 vpwr vgnd scs8hd_fill_2
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_10_76 vgnd vpwr scs8hd_decap_12
XFILLER_10_98 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_15_367 vgnd vpwr scs8hd_decap_6
X_077_ _076_/X _078_/C vgnd vpwr scs8hd_buf_1
XFILLER_2_271 vpwr vgnd scs8hd_fill_2
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_337 vgnd vpwr scs8hd_decap_12
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _096_/HI _088_/Y mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_11 vpwr vgnd scs8hd_fill_2
XFILLER_7_55 vgnd vpwr scs8hd_decap_4
XFILLER_7_330 vgnd vpwr scs8hd_decap_12
XFILLER_11_381 vgnd vpwr scs8hd_decap_12
XFILLER_8_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_178 vgnd vpwr scs8hd_decap_12
XFILLER_1_336 vgnd vpwr scs8hd_fill_1
XFILLER_4_23 vpwr vgnd scs8hd_fill_2
XFILLER_4_185 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _074_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__040__A _040_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_43 vgnd vpwr scs8hd_decap_12
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XFILLER_6_247 vgnd vpwr scs8hd_decap_6
X_093_ _093_/HI _093_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_276 vgnd vpwr scs8hd_decap_12
XFILLER_1_13 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_239 vgnd vpwr scs8hd_decap_3
XFILLER_10_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
X_076_ _066_/C _081_/B _076_/X vgnd vpwr scs8hd_or2_4
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _052_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_349 vgnd vpwr scs8hd_decap_12
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _058_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_342 vgnd vpwr scs8hd_decap_12
XFILLER_7_375 vgnd vpwr scs8hd_decap_12
XFILLER_11_393 vgnd vpwr scs8hd_decap_12
X_059_ _071_/A _058_/B _059_/C _058_/D _059_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__043__A _043_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_8_128 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__038__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_315 vgnd vpwr scs8hd_decap_4
XFILLER_0_370 vpwr vgnd scs8hd_fill_2
XFILLER_4_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__051__A _046_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_6_226 vpwr vgnd scs8hd_fill_2
XFILLER_10_211 vgnd vpwr scs8hd_decap_3
X_092_ _092_/HI _092_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_288 vgnd vpwr scs8hd_decap_12
XFILLER_18_300 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _091_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__046__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vgnd vpwr scs8hd_decap_8
XFILLER_10_45 vgnd vpwr scs8hd_decap_4
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
X_075_ address[4] _075_/X vgnd vpwr scs8hd_buf_1
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_8 vgnd vpwr scs8hd_decap_3
X_058_ _071_/A _058_/B _040_/X _058_/D _058_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_387 vgnd vpwr scs8hd_decap_12
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_313 vgnd vpwr scs8hd_decap_8
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vpwr vgnd scs8hd_fill_2
XFILLER_7_195 vpwr vgnd scs8hd_fill_2
XANTENNA__054__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_349 vpwr vgnd scs8hd_fill_2
XFILLER_9_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_110 vgnd vpwr scs8hd_decap_3
XFILLER_4_154 vgnd vpwr scs8hd_decap_4
XFILLER_4_69 vpwr vgnd scs8hd_fill_2
XANTENNA__049__A _071_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_202 vpwr vgnd scs8hd_fill_2
XFILLER_9_213 vpwr vgnd scs8hd_fill_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__051__B _058_/B vgnd vpwr scs8hd_diode_2
X_091_ _091_/A _091_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_312 vgnd vpwr scs8hd_decap_12
XFILLER_5_282 vpwr vgnd scs8hd_fill_2
XANTENNA__046__B _046_/B vgnd vpwr scs8hd_diode_2
XANTENNA__062__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ _074_/A _074_/B _074_/C _067_/X _074_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__057__A _046_/A vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
X_057_ _046_/A _046_/B _059_/C _058_/D _057_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_47 vpwr vgnd scs8hd_fill_2
XFILLER_7_399 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _091_/Y mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_108 vpwr vgnd scs8hd_fill_2
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_130 vgnd vpwr scs8hd_decap_4
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_109_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_19_281 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__054__B _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_339 vgnd vpwr scs8hd_fill_1
XFILLER_4_144 vgnd vpwr scs8hd_decap_3
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA__049__B _058_/B vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_12
XANTENNA__051__C _040_/X vgnd vpwr scs8hd_diode_2
X_090_ _090_/A _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_206 vgnd vpwr scs8hd_decap_3
XFILLER_6_3 vgnd vpwr scs8hd_decap_3
XFILLER_1_38 vpwr vgnd scs8hd_fill_2
XFILLER_1_49 vpwr vgnd scs8hd_fill_2
XFILLER_18_324 vgnd vpwr scs8hd_decap_12
XANTENNA__046__C _059_/C vgnd vpwr scs8hd_diode_2
XANTENNA__062__B _074_/B vgnd vpwr scs8hd_diode_2
X_073_ _074_/A _074_/B _078_/D _067_/X _073_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_253 vpwr vgnd scs8hd_fill_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_70 vgnd vpwr scs8hd_decap_3
XANTENNA__057__B _046_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A _074_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XFILLER_7_26 vpwr vgnd scs8hd_fill_2
XFILLER_11_330 vgnd vpwr scs8hd_decap_12
X_056_ _046_/A _046_/B _040_/X _058_/D _056_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_367 vgnd vpwr scs8hd_decap_6
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XANTENNA__068__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
XFILLER_7_164 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
X_108_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_11_171 vgnd vpwr scs8hd_decap_12
X_039_ address[0] _040_/A vgnd vpwr scs8hd_inv_8
XFILLER_19_293 vgnd vpwr scs8hd_decap_12
XANTENNA__070__B _046_/B vgnd vpwr scs8hd_diode_2
XANTENNA__054__C _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_0_362 vgnd vpwr scs8hd_decap_8
XFILLER_0_351 vgnd vpwr scs8hd_decap_8
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__049__C _040_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_104 vgnd vpwr scs8hd_fill_1
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_3
XANTENNA__051__D _046_/D vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _066_/C vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _089_/Y mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_295 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_391 vgnd vpwr scs8hd_decap_12
XANTENNA__046__D _046_/D vgnd vpwr scs8hd_diode_2
XANTENNA__062__C _040_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_306 vgnd vpwr scs8hd_decap_12
XFILLER_2_210 vpwr vgnd scs8hd_fill_2
X_072_ _071_/A _074_/B _074_/C _067_/X _072_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_287 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _096_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_361 vgnd vpwr scs8hd_decap_12
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XANTENNA__057__C _059_/C vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XANTENNA__073__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
X_055_ _054_/X _058_/D vgnd vpwr scs8hd_buf_1
XFILLER_11_342 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B _046_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
X_038_ address[2] _046_/B vgnd vpwr scs8hd_inv_8
X_107_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__054__D address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__070__C _074_/C vgnd vpwr scs8hd_diode_2
XANTENNA__079__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_4_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _090_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__049__D _046_/D vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vgnd vpwr scs8hd_decap_4
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _058_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__076__B _081_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_5_252 vpwr vgnd scs8hd_fill_2
XANTENNA__062__D _058_/D vgnd vpwr scs8hd_diode_2
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_318 vgnd vpwr scs8hd_decap_12
X_071_ _071_/A _074_/B _078_/D _067_/X _071_/Y vgnd vpwr scs8hd_nor4_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XANTENNA__057__D _058_/D vgnd vpwr scs8hd_diode_2
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
XANTENNA__073__C _078_/D vgnd vpwr scs8hd_diode_2
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
X_054_ address[3] _081_/B _066_/A address[5] _054_/X vgnd vpwr scs8hd_or4_4
XFILLER_11_354 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _083_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_12
XANTENNA__068__C _078_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XANTENNA__084__B _080_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _046_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vpwr vgnd scs8hd_fill_2
X_037_ address[1] _046_/A vgnd vpwr scs8hd_buf_1
X_106_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_8_93 vgnd vpwr scs8hd_decap_6
XANTENNA__070__D _067_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__079__B address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_0_320 vgnd vpwr scs8hd_decap_3
XFILLER_16_276 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_217 vgnd vpwr scs8hd_decap_3
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_8_261 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
XFILLER_5_231 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _073_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _074_/A _046_/B _074_/C _067_/X _070_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_267 vpwr vgnd scs8hd_fill_2
XFILLER_4_3 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _097_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_2_62 vgnd vpwr scs8hd_decap_8
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XANTENNA__073__D _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
XANTENNA__098__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
X_053_ address[4] _066_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_60 vgnd vpwr scs8hd_fill_1
XFILLER_11_377 vpwr vgnd scs8hd_fill_2
XANTENNA__068__D _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA__084__C _078_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_101 vgnd vpwr scs8hd_fill_1
X_105_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _051_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__079__C _078_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_115 vpwr vgnd scs8hd_fill_2
XFILLER_16_288 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _057_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_12
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_240 vgnd vpwr scs8hd_fill_1
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_84 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_265 vpwr vgnd scs8hd_fill_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_2_257 vgnd vpwr scs8hd_fill_1
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_96 vpwr vgnd scs8hd_fill_2
XFILLER_2_41 vpwr vgnd scs8hd_fill_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
XFILLER_11_367 vgnd vpwr scs8hd_decap_4
X_052_ _046_/A _058_/B _059_/C _046_/D _052_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__084__D _078_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _091_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_168 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
X_104_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_3_330 vgnd vpwr scs8hd_decap_12
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_84 vgnd vpwr scs8hd_decap_8
XANTENNA__079__D _074_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_333 vpwr vgnd scs8hd_fill_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _095_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_163 vpwr vgnd scs8hd_fill_2
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XFILLER_6_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_19 vpwr vgnd scs8hd_fill_2
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_051_ _046_/A _058_/B _040_/X _046_/D _051_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_306 vgnd vpwr scs8hd_decap_12
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_361 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
XFILLER_11_110 vgnd vpwr scs8hd_decap_12
XFILLER_7_147 vpwr vgnd scs8hd_fill_2
X_103_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_3_342 vgnd vpwr scs8hd_decap_12
XFILLER_14_7 vgnd vpwr scs8hd_decap_12
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _063_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_209 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _086_/A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_278 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_330 vgnd vpwr scs8hd_decap_12
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_300 vgnd vpwr scs8hd_decap_12
XFILLER_14_377 vgnd vpwr scs8hd_decap_12
XFILLER_2_32 vgnd vpwr scs8hd_decap_6
XFILLER_1_292 vgnd vpwr scs8hd_fill_1
XFILLER_1_270 vgnd vpwr scs8hd_fill_1
XFILLER_17_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_381 vgnd vpwr scs8hd_decap_4
X_050_ _071_/A _058_/B _059_/C _046_/D _050_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_318 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_3
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_19_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _051_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_19 vgnd vpwr scs8hd_decap_12
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_354 vgnd vpwr scs8hd_decap_12
XFILLER_7_115 vgnd vpwr scs8hd_decap_4
XFILLER_7_126 vpwr vgnd scs8hd_fill_2
X_102_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_64 vgnd vpwr scs8hd_decap_12
XFILLER_0_302 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__104__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_405 vpwr vgnd scs8hd_fill_2
XFILLER_0_198 vpwr vgnd scs8hd_fill_2
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_265 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XFILLER_5_32 vpwr vgnd scs8hd_fill_2
XFILLER_5_65 vpwr vgnd scs8hd_fill_2
XFILLER_5_235 vpwr vgnd scs8hd_fill_2
XFILLER_17_342 vgnd vpwr scs8hd_decap_12
XFILLER_2_249 vpwr vgnd scs8hd_fill_2
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_312 vgnd vpwr scs8hd_decap_12
XFILLER_14_389 vgnd vpwr scs8hd_decap_8
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_2_22 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_decap_4
XFILLER_9_393 vgnd vpwr scs8hd_decap_12
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
XFILLER_11_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_6_385 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
X_101_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_6_171 vgnd vpwr scs8hd_decap_4
XFILLER_8_76 vgnd vpwr scs8hd_decap_4
XFILLER_6_193 vpwr vgnd scs8hd_fill_2
XFILLER_4_119 vpwr vgnd scs8hd_fill_2
XFILLER_0_325 vpwr vgnd scs8hd_fill_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_281 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_11 vpwr vgnd scs8hd_fill_2
XFILLER_8_244 vgnd vpwr scs8hd_decap_8
XFILLER_8_288 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_88 vpwr vgnd scs8hd_fill_2
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_6
XFILLER_17_354 vgnd vpwr scs8hd_decap_12
XFILLER_2_228 vpwr vgnd scs8hd_fill_2
XFILLER_2_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _090_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_324 vgnd vpwr scs8hd_decap_12
XFILLER_2_12 vgnd vpwr scs8hd_decap_3
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_98 vgnd vpwr scs8hd_decap_12
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
X_100_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_6
XFILLER_0_337 vpwr vgnd scs8hd_fill_2
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_12_7 vgnd vpwr scs8hd_decap_8
XFILLER_15_293 vgnd vpwr scs8hd_decap_12
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_167 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XANTENNA__041__A enable vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_248 vpwr vgnd scs8hd_fill_2
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_1_284 vpwr vgnd scs8hd_fill_2
XFILLER_1_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_12
XFILLER_11_11 vpwr vgnd scs8hd_fill_2
XFILLER_11_22 vpwr vgnd scs8hd_fill_2
XFILLER_11_33 vgnd vpwr scs8hd_decap_4
XFILLER_11_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_361 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_9_170 vpwr vgnd scs8hd_fill_2
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_192 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_0_3 vgnd vpwr scs8hd_decap_3
XFILLER_3_313 vpwr vgnd scs8hd_fill_2
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _072_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_269 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_45 vgnd vpwr scs8hd_decap_4
XANTENNA__044__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XFILLER_3_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__039__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_113 vgnd vpwr scs8hd_decap_4
XFILLER_8_224 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _050_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_367 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A _046_/A vgnd vpwr scs8hd_diode_2
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _056_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_12
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_1_296 vpwr vgnd scs8hd_fill_2
XFILLER_9_330 vgnd vpwr scs8hd_decap_12
XANTENNA__047__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_318 vgnd vpwr scs8hd_decap_12
XFILLER_11_56 vgnd vpwr scs8hd_decap_4
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
XFILLER_9_182 vgnd vpwr scs8hd_fill_1
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _087_/A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_7_119 vgnd vpwr scs8hd_fill_1
XFILLER_11_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_089_ _089_/A _089_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_141 vpwr vgnd scs8hd_fill_2
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__044__B _046_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
XANTENNA__060__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_100 vpwr vgnd scs8hd_fill_2
XANTENNA__055__A _054_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_decap_12
XFILLER_5_36 vgnd vpwr scs8hd_decap_4
XFILLER_5_69 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_239 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_379 vgnd vpwr scs8hd_decap_12
XFILLER_4_283 vpwr vgnd scs8hd_fill_2
XANTENNA__052__B _058_/B vgnd vpwr scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XFILLER_14_349 vgnd vpwr scs8hd_decap_12
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_2_26 vgnd vpwr scs8hd_decap_4
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_342 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _056_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__063__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
XANTENNA__058__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_326 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_120 vgnd vpwr scs8hd_decap_3
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
X_088_ _088_/A _088_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA__044__C _040_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_329 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_159 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_288 vgnd vpwr scs8hd_decap_12
XFILLER_10_7 vgnd vpwr scs8hd_decap_8
XFILLER_7_281 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_218 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_251 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__052__C _059_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_decap_4
XFILLER_6_91 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_38 vgnd vpwr scs8hd_fill_1
XFILLER_9_354 vgnd vpwr scs8hd_decap_12
XANTENNA__063__B _074_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_335 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_8
XANTENNA__058__B _058_/B vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _089_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_087_ _087_/A _087_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__044__D _046_/D vgnd vpwr scs8hd_diode_2
XANTENNA__069__A address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _093_/HI _086_/Y mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_146 vpwr vgnd scs8hd_fill_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__071__B _074_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _095_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_293 vgnd vpwr scs8hd_decap_12
XANTENNA__066__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_403 vgnd vpwr scs8hd_decap_4
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_4_296 vgnd vpwr scs8hd_decap_8
XANTENNA__052__D _046_/D vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__077__A _076_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_288 vpwr vgnd scs8hd_fill_2
XFILLER_1_266 vgnd vpwr scs8hd_decap_4
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_9_377 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _093_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__063__C _059_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_174 vgnd vpwr scs8hd_decap_8
XFILLER_3_71 vpwr vgnd scs8hd_fill_2
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
XANTENNA__058__C _040_/X vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _074_/B vgnd vpwr scs8hd_diode_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_086_ _086_/A _086_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_2_394 vgnd vpwr scs8hd_decap_3
XFILLER_2_350 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_0_.latch data_in _091_/A _085_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__085__A _075_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
X_069_ address[0] _074_/C vgnd vpwr scs8hd_buf_1
XFILLER_0_94 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_117 vgnd vpwr scs8hd_fill_1
XFILLER_0_128 vgnd vpwr scs8hd_decap_4
XANTENNA__071__C _078_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_206 vpwr vgnd scs8hd_fill_2
XFILLER_8_228 vgnd vpwr scs8hd_decap_12
XFILLER_12_202 vgnd vpwr scs8hd_decap_12
XANTENNA__066__C _066_/C vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _080_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _063_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_93 vgnd vpwr scs8hd_decap_6
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_201 vpwr vgnd scs8hd_fill_2
XFILLER_2_18 vpwr vgnd scs8hd_fill_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _087_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_330 vgnd vpwr scs8hd_decap_12
XFILLER_9_367 vgnd vpwr scs8hd_decap_4
XFILLER_9_389 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XANTENNA__063__D _058_/D vgnd vpwr scs8hd_diode_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_300 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_6_337 vgnd vpwr scs8hd_decap_12
XFILLER_10_377 vgnd vpwr scs8hd_decap_12
XFILLER_9_131 vpwr vgnd scs8hd_fill_2
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XFILLER_5_381 vgnd vpwr scs8hd_decap_12
XANTENNA__058__D _058_/D vgnd vpwr scs8hd_diode_2
XANTENNA__074__C _074_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_8 vgnd vpwr scs8hd_decap_8
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_6_101 vpwr vgnd scs8hd_fill_2
X_085_ _075_/X _080_/Y _078_/C _074_/C _085_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_112 vgnd vpwr scs8hd_decap_8
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_167 vpwr vgnd scs8hd_fill_2
XFILLER_6_189 vpwr vgnd scs8hd_fill_2
XFILLER_2_362 vgnd vpwr scs8hd_decap_12
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XANTENNA__085__B _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_104 vpwr vgnd scs8hd_fill_2
X_068_ _074_/A _046_/B _078_/D _067_/X _068_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _068_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XANTENNA__071__D _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_19_391 vgnd vpwr scs8hd_decap_12
XANTENNA__066__D _081_/B vgnd vpwr scs8hd_diode_2
XANTENNA__082__C _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_306 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_361 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_1_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _059_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_342 vgnd vpwr scs8hd_decap_12
XFILLER_13_375 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_312 vgnd vpwr scs8hd_decap_12
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_6_305 vgnd vpwr scs8hd_decap_12
XFILLER_6_349 vgnd vpwr scs8hd_decap_12
XFILLER_10_389 vgnd vpwr scs8hd_decap_8
XFILLER_9_165 vpwr vgnd scs8hd_fill_2
XFILLER_9_198 vpwr vgnd scs8hd_fill_2
XFILLER_5_393 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
XANTENNA__074__D _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA__099__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_374 vgnd vpwr scs8hd_decap_12
X_084_ _075_/X _080_/Y _078_/C _078_/D _084_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XANTENNA__085__C _078_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_171 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _049_/Y vgnd vpwr scs8hd_diode_2
X_067_ _067_/A _067_/X vgnd vpwr scs8hd_buf_1
XFILLER_0_63 vgnd vpwr scs8hd_decap_6
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_9_94 vgnd vpwr scs8hd_fill_1
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_252 vpwr vgnd scs8hd_fill_2
XFILLER_11_281 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _071_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__082__D _078_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_318 vgnd vpwr scs8hd_decap_12
XFILLER_4_222 vpwr vgnd scs8hd_fill_2
XFILLER_4_266 vgnd vpwr scs8hd_decap_8
XFILLER_6_51 vgnd vpwr scs8hd_fill_1
XFILLER_6_84 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _088_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_159 vgnd vpwr scs8hd_decap_12
XFILLER_13_354 vgnd vpwr scs8hd_decap_12
XFILLER_13_387 vgnd vpwr scs8hd_decap_12
XFILLER_0_291 vpwr vgnd scs8hd_fill_2
XFILLER_11_18 vpwr vgnd scs8hd_fill_2
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_317 vgnd vpwr scs8hd_decap_12
XFILLER_10_324 vgnd vpwr scs8hd_decap_12
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_52 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _049_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_96 vpwr vgnd scs8hd_fill_2
XFILLER_3_309 vpwr vgnd scs8hd_fill_2
X_083_ _075_/X _080_/Y _081_/X _074_/C _083_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_110 vgnd vpwr scs8hd_decap_12
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_386 vgnd vpwr scs8hd_decap_8
XFILLER_18_276 vgnd vpwr scs8hd_decap_12
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XANTENNA__085__D _074_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_066_ _066_/A address[5] _066_/C _081_/B _067_/A vgnd vpwr scs8hd_or4_4
XFILLER_9_51 vpwr vgnd scs8hd_fill_2
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_293 vgnd vpwr scs8hd_decap_12
X_049_ _071_/A _058_/B _040_/X _046_/D _049_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_63 vgnd vpwr scs8hd_decap_6
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_13_399 vgnd vpwr scs8hd_decap_8
XFILLER_0_270 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _087_/Y mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_6_329 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_9_123 vgnd vpwr scs8hd_decap_8
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_75 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vpwr vgnd scs8hd_fill_2
X_082_ _075_/X _080_/Y _081_/X _078_/D _082_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_10_122 vgnd vpwr scs8hd_decap_12
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_199 vgnd vpwr scs8hd_decap_12
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_288 vgnd vpwr scs8hd_decap_12
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_269 vgnd vpwr scs8hd_decap_12
X_065_ address[3] _066_/C vgnd vpwr scs8hd_inv_8
XFILLER_2_195 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_30 vpwr vgnd scs8hd_fill_2
XFILLER_9_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _086_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _094_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_048_ address[2] _058_/B vgnd vpwr scs8hd_buf_1
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
XFILLER_14_19 vgnd vpwr scs8hd_decap_12
XFILLER_4_279 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_1_205 vpwr vgnd scs8hd_fill_2
XFILLER_13_367 vgnd vpwr scs8hd_decap_6
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_337 vgnd vpwr scs8hd_decap_12
XFILLER_9_102 vpwr vgnd scs8hd_fill_2
XFILLER_9_157 vgnd vpwr scs8hd_decap_8
XFILLER_5_330 vgnd vpwr scs8hd_decap_12
XFILLER_3_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_134 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_081_ address[3] _081_/B _081_/X vgnd vpwr scs8hd_or2_4
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_108 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
X_064_ _040_/A _078_/D vgnd vpwr scs8hd_buf_1
XFILLER_0_44 vgnd vpwr scs8hd_fill_1
XANTENNA__110__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_9_86 vgnd vpwr scs8hd_decap_8
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XANTENNA__105__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
X_047_ address[1] _071_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _089_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_247 vpwr vgnd scs8hd_fill_2
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_6_43 vgnd vpwr scs8hd_decap_8
XFILLER_6_87 vgnd vpwr scs8hd_decap_4
XFILLER_3_291 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_9_306 vgnd vpwr scs8hd_decap_12
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_10_349 vgnd vpwr scs8hd_decap_12
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XFILLER_5_342 vgnd vpwr scs8hd_decap_12
XANTENNA__113__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_080_ address[5] _080_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_312 vgnd vpwr scs8hd_fill_1
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _052_/Y vgnd vpwr scs8hd_diode_2
X_063_ _074_/A _074_/B _059_/C _058_/D _063_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_175 vgnd vpwr scs8hd_fill_1
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_78 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vgnd vpwr scs8hd_decap_4
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
X_046_ _046_/A _046_/B _059_/C _046_/D _046_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_212 vpwr vgnd scs8hd_fill_2
XFILLER_7_245 vgnd vpwr scs8hd_decap_4
XFILLER_7_256 vpwr vgnd scs8hd_fill_2
X_115_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_330 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_1_.latch data_in _090_/A _084_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_226 vpwr vgnd scs8hd_fill_2
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XFILLER_16_300 vgnd vpwr scs8hd_decap_12
XFILLER_16_377 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_318 vgnd vpwr scs8hd_decap_12
XFILLER_15_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_0_295 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

