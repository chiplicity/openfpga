* NGSPICE file created from sb_3__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt sb_3__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_
+ bottom_right_grid_pin_15_ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_
+ bottom_right_grid_pin_7_ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_12_ left_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ top_right_grid_pin_13_ top_right_grid_pin_15_ top_right_grid_pin_1_ top_right_grid_pin_3_
+ top_right_grid_pin_5_ top_right_grid_pin_7_ top_right_grid_pin_9_ vpwr vgnd
XFILLER_22_122 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_85 vgnd vpwr scs8hd_decap_6
XFILLER_13_133 vpwr vgnd scs8hd_fill_2
XFILLER_9_137 vpwr vgnd scs8hd_fill_2
XFILLER_9_159 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _110_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_1_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _166_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_107 vpwr vgnd scs8hd_fill_2
XFILLER_10_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_206 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _156_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _066_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_131_ _101_/A _135_/B _131_/Y vgnd vpwr scs8hd_nor2_4
X_062_ address[5] _152_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_165 vgnd vpwr scs8hd_fill_1
XFILLER_2_132 vgnd vpwr scs8hd_fill_1
XANTENNA__119__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
XFILLER_14_272 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _183_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_213 vpwr vgnd scs8hd_fill_2
XFILLER_11_231 vpwr vgnd scs8hd_fill_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
X_114_ _106_/A _110_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _080_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _116_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_4_205 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _164_/HI _070_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__116__B _148_/C vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_25_142 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_98 vpwr vgnd scs8hd_fill_2
XFILLER_0_252 vpwr vgnd scs8hd_fill_2
XFILLER_0_241 vgnd vpwr scs8hd_decap_6
XFILLER_31_156 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_186 vgnd vpwr scs8hd_decap_8
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_234 vgnd vpwr scs8hd_decap_8
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _156_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_145 vpwr vgnd scs8hd_fill_2
XFILLER_22_101 vpwr vgnd scs8hd_fill_2
XFILLER_26_64 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_3
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_13_178 vgnd vpwr scs8hd_decap_3
XFILLER_3_68 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_160 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _158_/HI _067_/Y mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _172_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_215 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _082_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
X_130_ address[6] _152_/B _100_/B _135_/B vgnd vpwr scs8hd_or3_4
XFILLER_15_229 vpwr vgnd scs8hd_fill_2
X_061_ address[6] _145_/A vgnd vpwr scs8hd_inv_8
XFILLER_2_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XFILLER_9_34 vgnd vpwr scs8hd_decap_4
XANTENNA__135__A _105_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _176_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _073_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_210 vpwr vgnd scs8hd_fill_2
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
X_113_ _105_/A _110_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_66 vpwr vgnd scs8hd_fill_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_42 vpwr vgnd scs8hd_fill_2
XFILLER_28_184 vpwr vgnd scs8hd_fill_2
XANTENNA__132__B _135_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _069_/A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_140 vpwr vgnd scs8hd_fill_2
XFILLER_19_173 vgnd vpwr scs8hd_decap_4
XFILLER_19_195 vgnd vpwr scs8hd_decap_4
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.LATCH_1_.latch data_in _070_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_154 vpwr vgnd scs8hd_fill_2
XFILLER_31_32 vgnd vpwr scs8hd_decap_12
XFILLER_16_121 vpwr vgnd scs8hd_fill_2
XFILLER_31_168 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _128_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XFILLER_16_165 vgnd vpwr scs8hd_decap_6
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_39_224 vgnd vpwr scs8hd_decap_3
XFILLER_22_168 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_146 vgnd vpwr scs8hd_decap_4
XFILLER_13_157 vgnd vpwr scs8hd_decap_4
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_21_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _179_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _073_/Y mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_8_183 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_138 vgnd vpwr scs8hd_decap_6
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _075_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_271 vgnd vpwr scs8hd_decap_4
XFILLER_18_205 vgnd vpwr scs8hd_fill_1
XFILLER_18_227 vpwr vgnd scs8hd_fill_2
XFILLER_5_197 vgnd vpwr scs8hd_decap_3
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vpwr vgnd scs8hd_fill_2
XFILLER_23_263 vgnd vpwr scs8hd_decap_12
XFILLER_23_241 vgnd vpwr scs8hd_decap_3
XFILLER_23_44 vpwr vgnd scs8hd_fill_2
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
X_060_ address[0] _145_/D vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
X_189_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_244 vgnd vpwr scs8hd_decap_8
XANTENNA__061__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vpwr vgnd scs8hd_fill_2
XFILLER_18_22 vgnd vpwr scs8hd_decap_4
XFILLER_18_44 vgnd vpwr scs8hd_fill_1
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_112_ _104_/A _110_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_108 vgnd vpwr scs8hd_decap_8
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_163 vgnd vpwr scs8hd_decap_8
XFILLER_6_36 vgnd vpwr scs8hd_decap_4
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
XFILLER_25_188 vpwr vgnd scs8hd_fill_2
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XFILLER_31_66 vgnd vpwr scs8hd_decap_6
XFILLER_31_44 vgnd vpwr scs8hd_decap_6
XFILLER_31_11 vgnd vpwr scs8hd_decap_12
XFILLER_0_276 vgnd vpwr scs8hd_fill_1
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_158 vgnd vpwr scs8hd_fill_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_107 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_103 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__138__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__064__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_12_35 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _098_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _148_/C vgnd vpwr scs8hd_diode_2
Xmem_left_track_15.LATCH_0_.latch data_in _081_/A _152_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_250 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_80 vgnd vpwr scs8hd_decap_12
XFILLER_23_220 vpwr vgnd scs8hd_fill_2
XANTENNA__059__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_168 vgnd vpwr scs8hd_decap_6
XFILLER_2_157 vpwr vgnd scs8hd_fill_2
XFILLER_2_135 vgnd vpwr scs8hd_fill_1
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_188_ _188_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__151__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_212 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
X_111_ _103_/A _110_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_6_260 vgnd vpwr scs8hd_decap_12
XFILLER_4_219 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_12
XFILLER_29_77 vgnd vpwr scs8hd_decap_4
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_89 vpwr vgnd scs8hd_fill_2
XFILLER_31_78 vgnd vpwr scs8hd_decap_3
XFILLER_31_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_233 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_204 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _068_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_80 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _083_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in _066_/A _137_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__C _145_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__154__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _170_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XANTENNA__140__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_14_232 vpwr vgnd scs8hd_fill_2
XFILLER_14_243 vgnd vpwr scs8hd_decap_8
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__151__C _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_180 vgnd vpwr scs8hd_decap_3
XFILLER_1_191 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _102_/A _110_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_235 vpwr vgnd scs8hd_fill_2
XFILLER_11_257 vgnd vpwr scs8hd_decap_3
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA__146__C _145_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_209 vgnd vpwr scs8hd_decap_4
XFILLER_29_23 vgnd vpwr scs8hd_decap_12
XFILLER_3_242 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vpwr vgnd scs8hd_fill_2
XFILLER_19_165 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _159_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_146 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vgnd vpwr scs8hd_decap_4
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_69 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_256 vgnd vpwr scs8hd_decap_12
XFILLER_0_223 vpwr vgnd scs8hd_fill_2
XFILLER_31_105 vgnd vpwr scs8hd_decap_6
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__D _145_/D vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_216 vpwr vgnd scs8hd_fill_2
XFILLER_22_149 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _067_/A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_26_68 vpwr vgnd scs8hd_fill_2
XFILLER_26_13 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_182 vgnd vpwr scs8hd_fill_1
XFILLER_21_171 vgnd vpwr scs8hd_decap_4
XANTENNA__138__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_131 vpwr vgnd scs8hd_fill_2
XFILLER_8_164 vpwr vgnd scs8hd_fill_2
XFILLER_8_186 vpwr vgnd scs8hd_fill_2
XFILLER_12_193 vpwr vgnd scs8hd_fill_2
XANTENNA__154__C _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_119 vgnd vpwr scs8hd_decap_8
XFILLER_12_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _072_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_208 vgnd vpwr scs8hd_decap_6
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__149__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_263 vgnd vpwr scs8hd_decap_12
XANTENNA__181__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_233 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _071_/Y mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_16 vgnd vpwr scs8hd_decap_4
X_186_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_13_91 vgnd vpwr scs8hd_fill_1
XANTENNA__151__D _145_/D vgnd vpwr scs8hd_diode_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _077_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_11_214 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _169_/HI _169_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XFILLER_1_72 vpwr vgnd scs8hd_fill_2
XFILLER_20_15 vpwr vgnd scs8hd_fill_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_46 vgnd vpwr scs8hd_decap_4
XFILLER_29_35 vgnd vpwr scs8hd_decap_4
XFILLER_28_122 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_188 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_17 vgnd vpwr scs8hd_decap_12
XFILLER_10_70 vpwr vgnd scs8hd_fill_2
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XFILLER_19_199 vgnd vpwr scs8hd_fill_1
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_158 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _074_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_268 vgnd vpwr scs8hd_decap_8
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_30_194 vgnd vpwr scs8hd_decap_12
XFILLER_30_183 vgnd vpwr scs8hd_decap_8
XFILLER_15_191 vpwr vgnd scs8hd_fill_2
XANTENNA__184__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_47 vgnd vpwr scs8hd_decap_6
XFILLER_26_25 vgnd vpwr scs8hd_fill_1
XANTENNA__094__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XANTENNA__154__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _111_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XFILLER_5_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__D _145_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_4
XFILLER_17_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_8
XFILLER_23_26 vgnd vpwr scs8hd_decap_3
XANTENNA__091__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
X_185_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_29_6 vgnd vpwr scs8hd_decap_3
XFILLER_20_215 vgnd vpwr scs8hd_decap_4
XFILLER_20_204 vgnd vpwr scs8hd_decap_8
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_26 vgnd vpwr scs8hd_fill_1
XANTENNA__086__B address[4] vgnd vpwr scs8hd_diode_2
X_168_ _168_/HI _168_/LO vgnd vpwr scs8hd_conb_1
X_099_ _115_/A address[4] _115_/C _100_/B vgnd vpwr scs8hd_or3_4
XFILLER_37_134 vgnd vpwr scs8hd_decap_12
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
XFILLER_1_62 vgnd vpwr scs8hd_decap_4
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XFILLER_28_134 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
XFILLER_3_222 vgnd vpwr scs8hd_decap_12
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_115 vpwr vgnd scs8hd_fill_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_15_38 vgnd vpwr scs8hd_decap_4
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_104 vpwr vgnd scs8hd_fill_2
XFILLER_16_148 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XFILLER_24_192 vgnd vpwr scs8hd_fill_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_30_140 vgnd vpwr scs8hd_decap_12
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_140 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_129 vpwr vgnd scs8hd_fill_2
XFILLER_21_184 vgnd vpwr scs8hd_decap_4
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_fill_1
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XFILLER_12_162 vgnd vpwr scs8hd_fill_1
XANTENNA__195__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__089__B _059_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _066_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_254 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__091__C _145_/D vgnd vpwr scs8hd_diode_2
XFILLER_2_139 vgnd vpwr scs8hd_decap_12
XFILLER_2_128 vgnd vpwr scs8hd_decap_4
XFILLER_14_202 vpwr vgnd scs8hd_fill_2
X_184_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_1_194 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__C _115_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_167_ _167_/HI _167_/LO vgnd vpwr scs8hd_conb_1
X_098_ _090_/A _106_/A _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_146 vgnd vpwr scs8hd_decap_12
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
XFILLER_1_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _082_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__097__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_234 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_92 vgnd vpwr scs8hd_decap_3
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_237 vpwr vgnd scs8hd_fill_2
XFILLER_0_204 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vgnd vpwr scs8hd_decap_8
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _168_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XFILLER_21_71 vgnd vpwr scs8hd_decap_4
XFILLER_21_60 vgnd vpwr scs8hd_fill_1
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__089__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_148 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _178_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_107 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_1_151 vgnd vpwr scs8hd_decap_3
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_228 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_239 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_9_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_71 vpwr vgnd scs8hd_fill_2
X_166_ _166_/HI _166_/LO vgnd vpwr scs8hd_conb_1
X_097_ address[1] address[2] address[0] _106_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _069_/Y mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_158 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _075_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__097__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vgnd vpwr scs8hd_decap_6
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_19_169 vpwr vgnd scs8hd_fill_2
X_149_ _145_/A _152_/B _142_/C _145_/D _149_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _160_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_29 vgnd vpwr scs8hd_decap_3
XFILLER_31_28 vpwr vgnd scs8hd_fill_2
XFILLER_0_227 vgnd vpwr scs8hd_decap_6
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XFILLER_24_161 vgnd vpwr scs8hd_fill_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_183 vgnd vpwr scs8hd_fill_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _157_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_17 vgnd vpwr scs8hd_decap_8
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_6
XFILLER_16_83 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_135 vgnd vpwr scs8hd_fill_1
XFILLER_8_179 vgnd vpwr scs8hd_decap_4
XFILLER_12_197 vgnd vpwr scs8hd_decap_4
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_3
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_259 vpwr vgnd scs8hd_fill_2
XFILLER_23_237 vpwr vgnd scs8hd_fill_2
XFILLER_23_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_119 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_182_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_226 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_252 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_13_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
XFILLER_24_50 vgnd vpwr scs8hd_decap_4
X_165_ _165_/HI _165_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_211 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _090_/A _105_/A _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_27_6 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _096_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_19 vpwr vgnd scs8hd_fill_2
Xmem_left_track_15.LATCH_1_.latch data_in _080_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_10_74 vgnd vpwr scs8hd_fill_1
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XFILLER_27_170 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _067_/A vgnd vpwr
+ scs8hd_diode_2
X_148_ _145_/A address[5] _148_/C address[0] _148_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_25_3 vgnd vpwr scs8hd_fill_1
X_079_ _079_/A _079_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_129 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_51 vpwr vgnd scs8hd_fill_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _090_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_110 vpwr vgnd scs8hd_fill_2
XFILLER_12_121 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_180 vgnd vpwr scs8hd_fill_1
XFILLER_26_235 vgnd vpwr scs8hd_decap_12
XFILLER_26_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_224 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_194 vpwr vgnd scs8hd_fill_2
XFILLER_4_161 vgnd vpwr scs8hd_decap_3
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
X_181_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_22_260 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_131 vgnd vpwr scs8hd_decap_4
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA__100__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_264 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_164_ _164_/HI _164_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
X_095_ address[1] address[2] _145_/D _105_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_201 vpwr vgnd scs8hd_fill_2
XFILLER_1_22 vgnd vpwr scs8hd_decap_12
XANTENNA__111__A _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ _145_/A address[5] _148_/C _145_/D _147_/Y vgnd vpwr scs8hd_nor4_4
X_078_ _078_/A _078_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_119 vgnd vpwr scs8hd_decap_3
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
XFILLER_16_108 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_10 vpwr vgnd scs8hd_fill_2
XFILLER_7_21 vgnd vpwr scs8hd_decap_4
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
XFILLER_7_76 vpwr vgnd scs8hd_fill_2
XFILLER_21_144 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_62 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _082_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XANTENNA__103__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_26_247 vgnd vpwr scs8hd_decap_12
XFILLER_5_118 vgnd vpwr scs8hd_decap_4
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_84 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_151 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_206 vpwr vgnd scs8hd_fill_2
XFILLER_22_272 vgnd vpwr scs8hd_decap_3
X_180_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_143 vgnd vpwr scs8hd_decap_8
XFILLER_1_176 vpwr vgnd scs8hd_fill_2
XFILLER_1_187 vgnd vpwr scs8hd_decap_4
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XANTENNA__109__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_276 vgnd vpwr scs8hd_fill_1
XFILLER_6_224 vgnd vpwr scs8hd_decap_12
X_094_ _090_/A _104_/A _094_/Y vgnd vpwr scs8hd_nor2_4
X_163_ _163_/HI _163_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__111__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _169_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_34 vgnd vpwr scs8hd_decap_12
XFILLER_1_89 vgnd vpwr scs8hd_decap_4
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _104_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_3
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_27_194 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_52 vgnd vpwr scs8hd_decap_4
XFILLER_19_106 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
X_077_ _077_/A _077_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__106__B _100_/X vgnd vpwr scs8hd_diode_2
X_146_ _145_/A address[5] _145_/C address[0] _146_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__122__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_109 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _067_/Y mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_8
XFILLER_24_186 vgnd vpwr scs8hd_decap_6
XFILLER_24_164 vpwr vgnd scs8hd_fill_2
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
Xmem_left_track_11.LATCH_1_.latch data_in _076_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
XFILLER_30_178 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vpwr vgnd scs8hd_fill_2
X_129_ _106_/A _128_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_178 vpwr vgnd scs8hd_fill_2
XFILLER_21_167 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
XFILLER_29_212 vgnd vpwr scs8hd_decap_12
XFILLER_16_53 vpwr vgnd scs8hd_fill_2
XFILLER_32_74 vgnd vpwr scs8hd_decap_6
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
XFILLER_12_178 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_26_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _077_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_52 vpwr vgnd scs8hd_fill_2
XFILLER_27_74 vpwr vgnd scs8hd_fill_2
Xmem_left_track_7.LATCH_0_.latch data_in _073_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_259 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _074_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_87 vgnd vpwr scs8hd_decap_4
XFILLER_1_100 vgnd vpwr scs8hd_decap_12
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
X_162_ _162_/HI _162_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_75 vgnd vpwr scs8hd_decap_6
X_093_ _091_/A address[2] address[0] _104_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_236 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_46 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_68 vpwr vgnd scs8hd_fill_2
XFILLER_10_55 vpwr vgnd scs8hd_fill_2
XFILLER_10_66 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_fill_1
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A address[5] _145_/C _145_/D _145_/Y vgnd vpwr scs8hd_nor4_4
X_076_ _076_/A _076_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
XFILLER_18_184 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _161_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_102 vgnd vpwr scs8hd_decap_12
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
X_128_ _105_/A _128_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__A _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
X_059_ address[2] _059_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_224 vgnd vpwr scs8hd_decap_12
XFILLER_12_102 vgnd vpwr scs8hd_decap_8
XFILLER_16_87 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_172 vpwr vgnd scs8hd_fill_2
XFILLER_7_194 vpwr vgnd scs8hd_fill_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_216 vpwr vgnd scs8hd_fill_2
XFILLER_4_175 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_68 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_274 vgnd vpwr scs8hd_decap_3
XFILLER_13_22 vgnd vpwr scs8hd_decap_3
XFILLER_1_112 vgnd vpwr scs8hd_decap_8
XFILLER_1_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _066_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__125__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_201 vgnd vpwr scs8hd_fill_1
XANTENNA__141__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_43 vgnd vpwr scs8hd_decap_4
XFILLER_10_200 vgnd vpwr scs8hd_decap_4
X_161_ _161_/HI _161_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_248 vgnd vpwr scs8hd_decap_12
X_092_ _090_/A _103_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_174 vgnd vpwr scs8hd_fill_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _169_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_144_ _145_/A address[5] _100_/B address[0] _144_/Y vgnd vpwr scs8hd_nor4_4
X_075_ _075_/A _075_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_177 vgnd vpwr scs8hd_decap_6
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_55 vgnd vpwr scs8hd_decap_3
XFILLER_21_88 vgnd vpwr scs8hd_decap_3
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_114 vgnd vpwr scs8hd_decap_6
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
X_127_ _104_/A _128_/B _127_/Y vgnd vpwr scs8hd_nor2_4
X_058_ address[1] _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _187_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[4] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_236 vgnd vpwr scs8hd_decap_8
XFILLER_16_11 vgnd vpwr scs8hd_fill_1
XFILLER_12_125 vgnd vpwr scs8hd_decap_4
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_fill_1
XANTENNA__128__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_184 vgnd vpwr scs8hd_fill_1
XFILLER_26_206 vgnd vpwr scs8hd_decap_8
XFILLER_27_21 vpwr vgnd scs8hd_fill_2
XFILLER_27_10 vgnd vpwr scs8hd_decap_4
XFILLER_4_198 vgnd vpwr scs8hd_decap_4
XFILLER_4_143 vgnd vpwr scs8hd_decap_8
XANTENNA__130__C _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_16_250 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _080_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_fill_1
XFILLER_1_168 vgnd vpwr scs8hd_decap_6
XFILLER_13_231 vgnd vpwr scs8hd_decap_3
XFILLER_9_213 vpwr vgnd scs8hd_fill_2
XFILLER_9_224 vpwr vgnd scs8hd_fill_2
XFILLER_9_235 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B address[5] vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.LATCH_0_.latch data_in _069_/A _140_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
X_091_ _091_/A address[2] _145_/D _103_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_205 vgnd vpwr scs8hd_decap_6
X_160_ _160_/HI _160_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_15 vgnd vpwr scs8hd_decap_4
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA__062__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_153 vgnd vpwr scs8hd_fill_1
XFILLER_19_44 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
X_074_ _074_/A _074_/Y vgnd vpwr scs8hd_inv_8
X_143_ _145_/A address[5] _100_/B _145_/D _143_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_2_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XFILLER_24_123 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_12 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_126_ _103_/A _128_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vgnd vpwr scs8hd_decap_8
XFILLER_12_148 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__144__B address[5] vgnd vpwr scs8hd_diode_2
X_109_ _101_/A _110_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_88 vpwr vgnd scs8hd_fill_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_221 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_122 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_262 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XANTENNA__065__A enable vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XANTENNA__141__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_56 vpwr vgnd scs8hd_fill_2
XFILLER_24_23 vgnd vpwr scs8hd_decap_6
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_235 vgnd vpwr scs8hd_decap_12
X_090_ _090_/A _102_/A _090_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_209 vpwr vgnd scs8hd_fill_2
XFILLER_10_36 vpwr vgnd scs8hd_fill_2
XFILLER_19_12 vgnd vpwr scs8hd_decap_4
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _083_/A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_23 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vgnd vpwr scs8hd_fill_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_198 vgnd vpwr scs8hd_decap_4
X_142_ _145_/A address[5] _142_/C address[0] _142_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
X_073_ _073_/A _073_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_242 vgnd vpwr scs8hd_decap_12
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _171_/A vgnd vpwr scs8hd_inv_1
XANTENNA__147__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_165 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XFILLER_24_157 vgnd vpwr scs8hd_decap_4
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _076_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_24 vgnd vpwr scs8hd_decap_4
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_168 vpwr vgnd scs8hd_fill_2
X_125_ _102_/A _128_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_14_190 vgnd vpwr scs8hd_fill_1
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _175_/A vgnd vpwr scs8hd_inv_1
XANTENNA__144__C _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_160 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
X_108_ _100_/A _145_/C _110_/B vgnd vpwr scs8hd_or2_4
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _192_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _067_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_233 vgnd vpwr scs8hd_decap_12
XFILLER_27_78 vgnd vpwr scs8hd_decap_4
XFILLER_27_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__139__C _148_/C vgnd vpwr scs8hd_diode_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_248 vpwr vgnd scs8hd_fill_2
XANTENNA__141__D _145_/D vgnd vpwr scs8hd_diode_2
XANTENNA__076__A _076_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _100_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_59 vgnd vpwr scs8hd_decap_4
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_177 vgnd vpwr scs8hd_decap_4
XFILLER_27_166 vpwr vgnd scs8hd_fill_2
X_141_ _145_/A address[5] _142_/C _145_/D _141_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_254 vgnd vpwr scs8hd_decap_12
X_072_ _072_/A _072_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_188 vpwr vgnd scs8hd_fill_2
XANTENNA__147__C _148_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _162_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _069_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_124_ _101_/A _128_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__084__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_176 vgnd vpwr scs8hd_decap_4
XFILLER_7_198 vpwr vgnd scs8hd_fill_2
XANTENNA__144__D address[0] vgnd vpwr scs8hd_diode_2
X_107_ address[3] _115_/B _115_/C _145_/C vgnd vpwr scs8hd_or3_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_35 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_242 vpwr vgnd scs8hd_fill_2
XFILLER_4_157 vpwr vgnd scs8hd_fill_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_3
XFILLER_4_179 vpwr vgnd scs8hd_fill_2
XANTENNA__139__D _145_/D vgnd vpwr scs8hd_diode_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _067_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_127 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XFILLER_13_212 vgnd vpwr scs8hd_decap_3
XANTENNA__182__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_260 vgnd vpwr scs8hd_decap_12
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_39_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.INVTX1_2_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_47 vgnd vpwr scs8hd_fill_1
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _078_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _090_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_230 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_156 vgnd vpwr scs8hd_fill_1
XANTENNA__087__A _100_/A vgnd vpwr scs8hd_diode_2
X_071_ _071_/A _071_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_140_ address[6] _152_/B _148_/C address[0] _140_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_266 vgnd vpwr scs8hd_decap_8
XFILLER_2_211 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XANTENNA__147__D _145_/D vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_104 vpwr vgnd scs8hd_fill_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _162_/HI _082_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_17 vpwr vgnd scs8hd_fill_2
XFILLER_7_28 vpwr vgnd scs8hd_fill_2
X_123_ address[6] _152_/B _142_/C _128_/B vgnd vpwr scs8hd_or3_4
XFILLER_16_7 vpwr vgnd scs8hd_fill_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__084__B _059_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_173 vgnd vpwr scs8hd_decap_4
X_106_ _106_/A _100_/X _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_155 vpwr vgnd scs8hd_fill_2
XFILLER_19_240 vgnd vpwr scs8hd_decap_4
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_60 vpwr vgnd scs8hd_fill_2
XFILLER_27_25 vgnd vpwr scs8hd_fill_1
XFILLER_40_257 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vgnd vpwr scs8hd_decap_12
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_191 vgnd vpwr scs8hd_decap_3
XFILLER_22_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_139 vpwr vgnd scs8hd_fill_2
XFILLER_9_217 vpwr vgnd scs8hd_fill_2
XFILLER_9_228 vgnd vpwr scs8hd_decap_4
XFILLER_9_239 vpwr vgnd scs8hd_fill_2
XFILLER_8_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_143 vgnd vpwr scs8hd_decap_12
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_24_15 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_6 vgnd vpwr scs8hd_decap_8
XFILLER_1_19 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
XFILLER_14_70 vpwr vgnd scs8hd_fill_2
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.LATCH_1_.latch data_in _072_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _077_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__193__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_19_48 vpwr vgnd scs8hd_fill_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA__087__B _142_/C vgnd vpwr scs8hd_diode_2
X_070_ _070_/A _070_/Y vgnd vpwr scs8hd_inv_8
XFILLER_33_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_102 vgnd vpwr scs8hd_decap_4
XFILLER_18_135 vgnd vpwr scs8hd_fill_1
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_16 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _090_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_122_ _106_/A _116_/X _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _081_/A mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_14_182 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XANTENNA__084__C _145_/D vgnd vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_49 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
XFILLER_20_174 vgnd vpwr scs8hd_decap_6
XFILLER_20_196 vpwr vgnd scs8hd_fill_2
XFILLER_28_274 vgnd vpwr scs8hd_fill_1
X_105_ _105_/A _100_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XFILLER_25_222 vpwr vgnd scs8hd_fill_2
XFILLER_40_269 vgnd vpwr scs8hd_decap_6
XANTENNA__095__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_258 vpwr vgnd scs8hd_fill_2
XFILLER_16_222 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _079_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_236 vgnd vpwr scs8hd_decap_8
XFILLER_22_203 vpwr vgnd scs8hd_fill_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_39_155 vgnd vpwr scs8hd_decap_12
XFILLER_5_84 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_6
XFILLER_10_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_81 vgnd vpwr scs8hd_decap_8
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_19_16 vgnd vpwr scs8hd_fill_1
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_117 vgnd vpwr scs8hd_decap_4
XFILLER_26_191 vgnd vpwr scs8hd_fill_1
XFILLER_26_180 vgnd vpwr scs8hd_decap_4
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_92 vpwr vgnd scs8hd_fill_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _155_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_74 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _066_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__B _106_/A vgnd vpwr scs8hd_diode_2
X_121_ _105_/A _116_/X _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_104_ _104_/A _100_/X _104_/Y vgnd vpwr scs8hd_nor2_4
Xmem_left_track_17.LATCH_0_.latch data_in _083_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vgnd vpwr scs8hd_fill_1
XFILLER_22_71 vpwr vgnd scs8hd_fill_2
XFILLER_7_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_8_73 vpwr vgnd scs8hd_fill_2
XFILLER_8_84 vgnd vpwr scs8hd_decap_6
XFILLER_40_215 vgnd vpwr scs8hd_decap_3
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_25_234 vgnd vpwr scs8hd_decap_8
XANTENNA__095__C _145_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XFILLER_33_81 vgnd vpwr scs8hd_decap_12
XFILLER_22_248 vgnd vpwr scs8hd_decap_12
XFILLER_5_30 vgnd vpwr scs8hd_decap_8
XFILLER_39_167 vgnd vpwr scs8hd_decap_12
XFILLER_39_101 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _068_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_80 vgnd vpwr scs8hd_fill_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _076_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _188_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_140 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_1_.latch data_in _068_/A _139_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_195 vpwr vgnd scs8hd_fill_2
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
XFILLER_23_151 vgnd vpwr scs8hd_decap_3
X_120_ _104_/A _116_/X _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_62 vgnd vpwr scs8hd_decap_4
XFILLER_11_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _103_/A _100_/X _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_143 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _161_/HI _080_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_221 vgnd vpwr scs8hd_decap_4
XFILLER_8_41 vpwr vgnd scs8hd_fill_2
XFILLER_6_191 vgnd vpwr scs8hd_fill_1
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XFILLER_27_17 vpwr vgnd scs8hd_fill_2
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_93 vgnd vpwr scs8hd_decap_12
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _158_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_179 vgnd vpwr scs8hd_decap_4
XFILLER_39_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_5_234 vgnd vpwr scs8hd_decap_8
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_149 vgnd vpwr scs8hd_decap_4
XFILLER_27_105 vgnd vpwr scs8hd_decap_4
XFILLER_4_6 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
X_196_ _196_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_3_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_108 vpwr vgnd scs8hd_fill_2
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _155_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _179_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
X_102_ _102_/A _100_/X _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_203 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _079_/A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_107 vpwr vgnd scs8hd_fill_2
XFILLER_17_62 vgnd vpwr scs8hd_decap_4
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _076_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_228 vgnd vpwr scs8hd_decap_4
Xmem_left_track_13.LATCH_0_.latch data_in _079_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_83 vgnd vpwr scs8hd_fill_1
XFILLER_0_143 vgnd vpwr scs8hd_decap_12
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_98 vgnd vpwr scs8hd_decap_4
XFILLER_5_43 vgnd vpwr scs8hd_decap_12
XFILLER_24_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _173_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _083_/Y mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_40 vpwr vgnd scs8hd_fill_2
XFILLER_5_213 vpwr vgnd scs8hd_fill_2
XFILLER_14_74 vgnd vpwr scs8hd_fill_1
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B _100_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_7_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_194 vgnd vpwr scs8hd_decap_3
XFILLER_26_161 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_161 vpwr vgnd scs8hd_fill_2
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _177_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_53 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _078_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_164 vpwr vgnd scs8hd_fill_2
XFILLER_14_186 vgnd vpwr scs8hd_decap_4
X_178_ _178_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_20_123 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_256 vgnd vpwr scs8hd_decap_12
XFILLER_28_223 vgnd vpwr scs8hd_decap_8
XFILLER_28_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_101_ _101_/A _100_/X _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_3
XFILLER_11_156 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_8
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_204 vpwr vgnd scs8hd_fill_2
XFILLER_16_215 vpwr vgnd scs8hd_fill_2
XFILLER_16_226 vgnd vpwr scs8hd_fill_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XANTENNA__104__B _100_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _069_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__120__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _074_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_207 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_122 vpwr vgnd scs8hd_fill_2
XFILLER_0_133 vpwr vgnd scs8hd_fill_2
XFILLER_0_199 vpwr vgnd scs8hd_fill_2
XFILLER_5_55 vgnd vpwr scs8hd_decap_6
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_88 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _136_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_53 vpwr vgnd scs8hd_fill_2
XFILLER_30_30 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_97 vpwr vgnd scs8hd_fill_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _067_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_184 vgnd vpwr scs8hd_fill_1
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_96 vpwr vgnd scs8hd_fill_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _071_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_154 vgnd vpwr scs8hd_fill_1
X_177_ _177_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA__107__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__123__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_28_213 vgnd vpwr scs8hd_fill_1
XFILLER_28_268 vgnd vpwr scs8hd_decap_6
X_100_ _100_/A _100_/B _100_/X vgnd vpwr scs8hd_or2_4
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_22_97 vpwr vgnd scs8hd_fill_2
XFILLER_19_202 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_183 vpwr vgnd scs8hd_fill_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_42 vgnd vpwr scs8hd_decap_3
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_142 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _160_/HI _078_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _069_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_63 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _102_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_241 vgnd vpwr scs8hd_decap_4
XFILLER_12_252 vgnd vpwr scs8hd_decap_8
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_67 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_127 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
XFILLER_30_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_108 vpwr vgnd scs8hd_fill_2
XFILLER_18_119 vgnd vpwr scs8hd_decap_4
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vgnd vpwr scs8hd_decap_4
X_193_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_68 vgnd vpwr scs8hd_decap_4
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_199 vgnd vpwr scs8hd_decap_4
XFILLER_11_66 vgnd vpwr scs8hd_fill_1
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
X_176_ _176_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__107__C _115_/C vgnd vpwr scs8hd_diode_2
XANTENNA__123__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_236 vgnd vpwr scs8hd_decap_12
XFILLER_11_103 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_45 vpwr vgnd scs8hd_fill_2
X_159_ _159_/HI _159_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__134__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_173 vgnd vpwr scs8hd_fill_1
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_8
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vgnd vpwr scs8hd_fill_1
XFILLER_3_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vpwr scs8hd_fill_1
XANTENNA__129__A _106_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _077_/A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_102 vgnd vpwr scs8hd_decap_12
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XFILLER_28_75 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_8_224 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _163_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _115_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_139 vpwr vgnd scs8hd_fill_2
XFILLER_14_22 vpwr vgnd scs8hd_fill_2
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_8
XFILLER_39_85 vpwr vgnd scs8hd_fill_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _128_/B vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_32 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _079_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _081_/Y mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_1_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_17_142 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_156 vgnd vpwr scs8hd_decap_4
XFILLER_23_134 vpwr vgnd scs8hd_fill_2
XFILLER_23_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_101 vpwr vgnd scs8hd_fill_2
XFILLER_14_112 vpwr vgnd scs8hd_fill_2
X_175_ _175_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__123__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_37_215 vgnd vpwr scs8hd_decap_12
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_248 vgnd vpwr scs8hd_decap_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_6
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_22_55 vgnd vpwr scs8hd_fill_1
XFILLER_22_22 vgnd vpwr scs8hd_decap_3
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_10_170 vpwr vgnd scs8hd_fill_2
XANTENNA__134__B _135_/B vgnd vpwr scs8hd_diode_2
X_089_ address[1] _059_/Y address[0] _102_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
X_158_ _158_/HI _158_/LO vgnd vpwr scs8hd_conb_1
XFILLER_26_3 vgnd vpwr scs8hd_fill_1
XANTENNA__150__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_207 vgnd vpwr scs8hd_decap_4
XANTENNA__060__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_229 vgnd vpwr scs8hd_fill_1
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_65 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__129__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_240 vgnd vpwr scs8hd_decap_4
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_232 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _081_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_114 vgnd vpwr scs8hd_decap_8
XFILLER_0_125 vgnd vpwr scs8hd_decap_8
XFILLER_8_236 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in _082_/A _153_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _072_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_29_195 vpwr vgnd scs8hd_fill_2
XFILLER_29_184 vpwr vgnd scs8hd_fill_2
XFILLER_29_140 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _167_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_6_90 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_187 vgnd vpwr scs8hd_decap_4
XFILLER_26_165 vgnd vpwr scs8hd_decap_4
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_4
XFILLER_1_253 vgnd vpwr scs8hd_decap_12
XFILLER_17_165 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_124 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_24 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_168 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _068_/Y vgnd vpwr
+ scs8hd_diode_2
X_174_ _174_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_37_227 vgnd vpwr scs8hd_decap_12
XFILLER_28_7 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _069_/A mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_127 vgnd vpwr scs8hd_decap_3
XFILLER_28_205 vpwr vgnd scs8hd_fill_2
XFILLER_3_91 vpwr vgnd scs8hd_fill_2
XANTENNA__058__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_22_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _157_/HI _157_/LO vgnd vpwr scs8hd_conb_1
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_120 vgnd vpwr scs8hd_decap_3
XFILLER_8_69 vpwr vgnd scs8hd_fill_2
XANTENNA__150__B _152_/B vgnd vpwr scs8hd_diode_2
X_088_ _101_/A _090_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_208 vpwr vgnd scs8hd_fill_2
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_89 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_156 vgnd vpwr scs8hd_decap_3
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_252 vpwr vgnd scs8hd_fill_2
XFILLER_15_263 vgnd vpwr scs8hd_decap_12
XANTENNA__145__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_222 vgnd vpwr scs8hd_fill_1
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_248 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_45 vgnd vpwr scs8hd_decap_8
XFILLER_30_12 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_30_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _070_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_152 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _159_/HI _076_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__C _142_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_right_grid_pin_5_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_80 vgnd vpwr scs8hd_decap_8
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
X_190_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_265 vgnd vpwr scs8hd_decap_12
XANTENNA__137__C _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_180 vgnd vpwr scs8hd_decap_3
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_173_ _173_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_37_239 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _075_/A mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _164_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A _074_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_139 vpwr vgnd scs8hd_fill_2
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_156_ _156_/HI _156_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_143 vpwr vgnd scs8hd_fill_2
XFILLER_10_183 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_087_ _100_/A _142_/C _090_/A vgnd vpwr scs8hd_or2_4
XFILLER_6_187 vgnd vpwr scs8hd_decap_4
XANTENNA__150__C _142_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XFILLER_18_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_242 vgnd vpwr scs8hd_decap_12
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_17_68 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_168 vpwr vgnd scs8hd_fill_2
XFILLER_3_146 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__C _145_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
X_139_ address[6] _152_/B _148_/C _145_/D _139_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_0_71 vgnd vpwr scs8hd_fill_1
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_256 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_205 vgnd vpwr scs8hd_decap_8
XFILLER_5_38 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_4
XFILLER_30_24 vgnd vpwr scs8hd_decap_6
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XFILLER_29_175 vpwr vgnd scs8hd_fill_2
XFILLER_29_164 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__142__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_112 vgnd vpwr scs8hd_fill_1
XFILLER_25_24 vpwr vgnd scs8hd_fill_2
XFILLER_25_13 vpwr vgnd scs8hd_fill_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
Xmem_left_track_13.LATCH_1_.latch data_in _078_/A _149_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_211 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_112 vpwr vgnd scs8hd_fill_2
XANTENNA__137__D _145_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _090_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_148 vgnd vpwr scs8hd_decap_3
X_172_ _172_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_141 vpwr vgnd scs8hd_fill_2
XANTENNA__148__C _148_/C vgnd vpwr scs8hd_diode_2
XANTENNA__180__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_163 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _079_/Y mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_14 vpwr vgnd scs8hd_fill_2
XFILLER_11_107 vpwr vgnd scs8hd_fill_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in _075_/A _146_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_251 vgnd vpwr scs8hd_fill_1
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XFILLER_8_49 vpwr vgnd scs8hd_fill_2
X_155_ _155_/HI _155_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_151 vpwr vgnd scs8hd_fill_2
X_086_ address[3] address[4] _115_/C _142_/C vgnd vpwr scs8hd_or3_4
XANTENNA__150__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XFILLER_18_273 vpwr vgnd scs8hd_fill_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_25 vpwr vgnd scs8hd_fill_2
XFILLER_17_47 vgnd vpwr scs8hd_decap_3
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_24_254 vgnd vpwr scs8hd_fill_1
XFILLER_24_210 vpwr vgnd scs8hd_fill_2
XANTENNA__085__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__145__D _145_/D vgnd vpwr scs8hd_diode_2
X_138_ address[6] _152_/B _145_/C address[0] _138_/Y vgnd vpwr scs8hd_nor4_4
X_069_ _069_/A _069_/Y vgnd vpwr scs8hd_inv_8
XFILLER_24_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_191 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_83 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_268 vgnd vpwr scs8hd_decap_8
XFILLER_9_81 vgnd vpwr scs8hd_decap_3
XFILLER_0_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _078_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_79 vgnd vpwr scs8hd_decap_4
XFILLER_28_57 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_26 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_89 vgnd vpwr scs8hd_decap_12
XFILLER_39_34 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _196_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_124 vpwr vgnd scs8hd_fill_2
XFILLER_25_47 vgnd vpwr scs8hd_decap_4
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_fill_1
XFILLER_17_146 vpwr vgnd scs8hd_fill_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _070_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__D _145_/D vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vpwr vgnd scs8hd_fill_2
XFILLER_23_116 vgnd vpwr scs8hd_decap_4
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XFILLER_11_49 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_116 vpwr vgnd scs8hd_fill_2
XFILLER_22_193 vgnd vpwr scs8hd_fill_1
X_171_ _171_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _135_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__148__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vgnd vpwr scs8hd_decap_4
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _080_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__090__B _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_274 vgnd vpwr scs8hd_decap_3
XFILLER_27_230 vgnd vpwr scs8hd_decap_3
XFILLER_6_167 vgnd vpwr scs8hd_decap_6
X_085_ address[6] address[5] _100_/A vgnd vpwr scs8hd_or2_4
X_154_ _145_/A _152_/B _145_/C address[0] _154_/Y vgnd vpwr scs8hd_nor4_4
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _166_/HI _074_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_69 vgnd vpwr scs8hd_decap_12
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _067_/A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__B address[5] vgnd vpwr scs8hd_diode_2
X_137_ address[6] _152_/B _145_/C _145_/D _137_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_068_ _068_/A _068_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_236 vgnd vpwr scs8hd_decap_8
XFILLER_21_214 vpwr vgnd scs8hd_fill_2
XFILLER_21_203 vgnd vpwr scs8hd_decap_8
XANTENNA__186__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _071_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _170_/A vgnd vpwr scs8hd_inv_1
XANTENNA__096__A _090_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_247 vpwr vgnd scs8hd_fill_2
XFILLER_5_18 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_49 vpwr vgnd scs8hd_fill_2
XFILLER_39_46 vgnd vpwr scs8hd_decap_12
XFILLER_29_144 vgnd vpwr scs8hd_fill_1
XFILLER_29_199 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_70 vgnd vpwr scs8hd_decap_3
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _174_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_50 vgnd vpwr scs8hd_decap_12
XPHY_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_19 vgnd vpwr scs8hd_fill_1
XFILLER_32_128 vgnd vpwr scs8hd_decap_12
XFILLER_32_117 vgnd vpwr scs8hd_decap_4
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _069_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__194__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_28 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_172 vgnd vpwr scs8hd_decap_4
X_170_ _170_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XFILLER_9_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_150 vgnd vpwr scs8hd_fill_1
XFILLER_28_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_95 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _073_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_49 vgnd vpwr scs8hd_decap_6
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _115_/A vgnd vpwr scs8hd_diode_2
X_153_ _145_/A _152_/B _145_/C _145_/D _153_/Y vgnd vpwr scs8hd_nor4_4
X_084_ address[1] _059_/Y _145_/D _101_/A vgnd vpwr scs8hd_or3_4
XFILLER_18_231 vgnd vpwr scs8hd_decap_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_15_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _073_/A mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_212 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.LATCH_0_.latch data_in _071_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ _106_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_067_ _067_/A _067_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_63 vgnd vpwr scs8hd_decap_8
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_21_248 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _167_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _103_/A _116_/X _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_230 vpwr vgnd scs8hd_fill_2
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_17 vgnd vpwr scs8hd_decap_3
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_40 vgnd vpwr scs8hd_fill_1
XFILLER_6_62 vgnd vpwr scs8hd_decap_4
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_8
XFILLER_26_81 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_85 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _165_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_254 vgnd vpwr scs8hd_decap_12
XFILLER_27_243 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_083_ _083_/A _083_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_125 vgnd vpwr scs8hd_decap_3
XFILLER_6_147 vgnd vpwr scs8hd_decap_6
XFILLER_10_154 vgnd vpwr scs8hd_decap_3
XFILLER_10_187 vpwr vgnd scs8hd_fill_2
X_152_ _145_/A _152_/B _100_/B address[0] _152_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _077_/Y mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_128 vpwr vgnd scs8hd_fill_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_066_ _066_/A _066_/Y vgnd vpwr scs8hd_inv_8
X_135_ _105_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_183 vgnd vpwr scs8hd_decap_8
XFILLER_2_161 vgnd vpwr scs8hd_decap_4
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_28_49 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
X_118_ _102_/A _116_/X _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_242 vpwr vgnd scs8hd_fill_2
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_4_223 vgnd vpwr scs8hd_decap_12
XFILLER_29_81 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_17 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_28 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_7 vgnd vpwr scs8hd_decap_3
XFILLER_25_171 vpwr vgnd scs8hd_fill_2
XFILLER_17_116 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XFILLER_31_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _081_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_182 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_230 vpwr vgnd scs8hd_fill_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_185 vgnd vpwr scs8hd_decap_8
XFILLER_22_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_3
XFILLER_13_174 vpwr vgnd scs8hd_fill_2
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _068_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_18 vpwr vgnd scs8hd_fill_2
XANTENNA__099__C _115_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_266 vgnd vpwr scs8hd_decap_8
XFILLER_10_144 vgnd vpwr scs8hd_fill_1
XFILLER_10_166 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vgnd vpwr scs8hd_decap_8
X_151_ _145_/A _152_/B _100_/B _145_/D _151_/Y vgnd vpwr scs8hd_nor4_4
X_082_ _082_/A _082_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _168_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_244 vgnd vpwr scs8hd_decap_8
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_29 vpwr vgnd scs8hd_fill_2
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_225 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_225 vpwr vgnd scs8hd_fill_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
XFILLER_23_83 vgnd vpwr scs8hd_fill_1
X_134_ _104_/A _135_/B _134_/Y vgnd vpwr scs8hd_nor2_4
X_065_ enable _115_/C vgnd vpwr scs8hd_inv_8
XFILLER_2_195 vpwr vgnd scs8hd_fill_2
XFILLER_2_151 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
XFILLER_28_28 vgnd vpwr scs8hd_decap_3
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _165_/HI _072_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_6
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _083_/A vgnd vpwr
+ scs8hd_diode_2
X_117_ _101_/A _116_/X _117_/Y vgnd vpwr scs8hd_nor2_4
Xmem_left_track_1.LATCH_0_.latch data_in _067_/A _138_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_37_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_235 vgnd vpwr scs8hd_decap_12
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_29_93 vpwr vgnd scs8hd_fill_2
XFILLER_26_128 vgnd vpwr scs8hd_decap_4
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XFILLER_31_83 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _163_/HI _069_/Y mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_194 vgnd vpwr scs8hd_fill_1
XFILLER_39_242 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vpwr vgnd scs8hd_fill_2
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _070_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_190 vpwr vgnd scs8hd_fill_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_6
X_150_ _145_/A _152_/B _142_/C address[0] _150_/Y vgnd vpwr scs8hd_nor4_4
X_081_ _081_/A _081_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_52 vgnd vpwr scs8hd_decap_4
XFILLER_12_63 vpwr vgnd scs8hd_fill_2
XFILLER_18_201 vgnd vpwr scs8hd_decap_4
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_5_160 vpwr vgnd scs8hd_fill_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_right_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_248 vpwr vgnd scs8hd_fill_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_95 vpwr vgnd scs8hd_fill_2
XFILLER_23_73 vgnd vpwr scs8hd_decap_4
XFILLER_23_51 vgnd vpwr scs8hd_decap_4
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
X_133_ _103_/A _135_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_064_ address[4] _115_/B vgnd vpwr scs8hd_inv_8
XANTENNA__110__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_7 vgnd vpwr scs8hd_decap_3
XFILLER_21_218 vpwr vgnd scs8hd_fill_2
XFILLER_9_20 vgnd vpwr scs8hd_fill_1
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_86 vpwr vgnd scs8hd_fill_2
XFILLER_28_18 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _071_/A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_40 vpwr vgnd scs8hd_fill_2
XFILLER_18_62 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_262 vgnd vpwr scs8hd_decap_12
X_116_ _100_/A _148_/C _116_/X vgnd vpwr scs8hd_or2_4
XFILLER_29_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_104 vpwr vgnd scs8hd_fill_2
XFILLER_37_170 vgnd vpwr scs8hd_decap_12
XFILLER_4_247 vgnd vpwr scs8hd_decap_12
XFILLER_6_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _072_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _106_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_217 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_129 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _075_/Y mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_132 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_154 vgnd vpwr scs8hd_decap_4
XFILLER_7_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_103 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_99 vgnd vpwr scs8hd_decap_4
XFILLER_3_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_235 vgnd vpwr scs8hd_decap_8
XFILLER_27_213 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_10_102 vgnd vpwr scs8hd_decap_8
X_080_ _080_/A _080_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _100_/A vgnd vpwr scs8hd_diode_2
X_132_ _102_/A _135_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_063_ address[3] _115_/A vgnd vpwr scs8hd_inv_8
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_0_78 vgnd vpwr scs8hd_fill_1
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_260 vgnd vpwr scs8hd_decap_12
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_20_252 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__105__B _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_234 vgnd vpwr scs8hd_decap_8
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_11_274 vgnd vpwr scs8hd_decap_3
X_115_ _115_/A _115_/B _115_/C _148_/C vgnd vpwr scs8hd_or3_4
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_1_.latch data_in _074_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__121__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_182 vgnd vpwr scs8hd_fill_1
XFILLER_4_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XFILLER_29_73 vpwr vgnd scs8hd_fill_2
XFILLER_28_171 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _100_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_66 vgnd vpwr scs8hd_fill_1
XFILLER_6_99 vgnd vpwr scs8hd_decap_6
XFILLER_26_108 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_fill_1
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_1_229 vgnd vpwr scs8hd_decap_12
XFILLER_17_108 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XFILLER_31_144 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _157_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

