magic
tech EFS8A
magscale 1 2
timestamp 1604337784
<< viali >>
rect 2329 12393 2363 12427
rect 17233 12325 17267 12359
rect 2145 12257 2179 12291
rect 16957 12257 16991 12291
rect 1593 11849 1627 11883
rect 2697 11849 2731 11883
rect 14105 11849 14139 11883
rect 20453 11849 20487 11883
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 2513 11645 2547 11679
rect 13921 11645 13955 11679
rect 20269 11645 20303 11679
rect 3157 11577 3191 11611
rect 2421 11509 2455 11543
rect 14565 11509 14599 11543
rect 17049 11509 17083 11543
rect 20913 11509 20947 11543
rect 2329 11305 2363 11339
rect 17491 11305 17525 11339
rect 17969 11237 18003 11271
rect 26792 11237 26826 11271
rect 2145 11169 2179 11203
rect 18061 11169 18095 11203
rect 26525 11169 26559 11203
rect 17877 11101 17911 11135
rect 27905 11033 27939 11067
rect 3341 10761 3375 10795
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 3157 10557 3191 10591
rect 3709 10557 3743 10591
rect 2145 10421 2179 10455
rect 17785 10421 17819 10455
rect 26617 10421 26651 10455
rect 26985 10421 27019 10455
rect 1593 10217 1627 10251
rect 8309 10217 8343 10251
rect 32321 10217 32355 10251
rect 1409 10081 1443 10115
rect 8125 10081 8159 10115
rect 32137 10081 32171 10115
rect 18153 9877 18187 9911
rect 18153 9673 18187 9707
rect 5733 9605 5767 9639
rect 7481 9605 7515 9639
rect 7941 9537 7975 9571
rect 17509 9537 17543 9571
rect 18613 9537 18647 9571
rect 5549 9469 5583 9503
rect 7297 9469 7331 9503
rect 18613 9401 18647 9435
rect 18705 9401 18739 9435
rect 1685 9333 1719 9367
rect 6193 9333 6227 9367
rect 8309 9333 8343 9367
rect 17877 9333 17911 9367
rect 32137 9333 32171 9367
rect 1685 9129 1719 9163
rect 21465 9061 21499 9095
rect 1501 8993 1535 9027
rect 21557 8993 21591 9027
rect 21373 8925 21407 8959
rect 21005 8857 21039 8891
rect 18153 8789 18187 8823
rect 1593 8585 1627 8619
rect 18153 8585 18187 8619
rect 21373 8585 21407 8619
rect 30665 8585 30699 8619
rect 32321 8585 32355 8619
rect 2329 8517 2363 8551
rect 21465 8449 21499 8483
rect 1409 8381 1443 8415
rect 1961 8381 1995 8415
rect 17785 8381 17819 8415
rect 18429 8381 18463 8415
rect 18705 8381 18739 8415
rect 20637 8381 20671 8415
rect 29009 8381 29043 8415
rect 29285 8381 29319 8415
rect 29541 8381 29575 8415
rect 32137 8381 32171 8415
rect 32689 8381 32723 8415
rect 17509 8313 17543 8347
rect 21005 8313 21039 8347
rect 18613 8245 18647 8279
rect 8677 8041 8711 8075
rect 9873 8041 9907 8075
rect 17785 8041 17819 8075
rect 29377 8041 29411 8075
rect 17877 7973 17911 8007
rect 1409 7905 1443 7939
rect 8493 7905 8527 7939
rect 9689 7905 9723 7939
rect 17785 7837 17819 7871
rect 1593 7769 1627 7803
rect 17325 7769 17359 7803
rect 1961 7497 1995 7531
rect 9137 7497 9171 7531
rect 17325 7497 17359 7531
rect 32321 7497 32355 7531
rect 1593 7429 1627 7463
rect 1409 7293 1443 7327
rect 2329 7293 2363 7327
rect 8953 7293 8987 7327
rect 16957 7293 16991 7327
rect 32137 7293 32171 7327
rect 32689 7293 32723 7327
rect 8493 7157 8527 7191
rect 9689 7157 9723 7191
rect 17601 7157 17635 7191
rect 19441 6885 19475 6919
rect 1501 6817 1535 6851
rect 19257 6817 19291 6851
rect 8953 6749 8987 6783
rect 19533 6749 19567 6783
rect 1685 6681 1719 6715
rect 18981 6681 19015 6715
rect 15945 6613 15979 6647
rect 1593 6409 1627 6443
rect 16037 6409 16071 6443
rect 18889 6409 18923 6443
rect 19349 6409 19383 6443
rect 32321 6409 32355 6443
rect 15853 6273 15887 6307
rect 16589 6273 16623 6307
rect 1409 6205 1443 6239
rect 32137 6205 32171 6239
rect 32689 6205 32723 6239
rect 16313 6137 16347 6171
rect 2053 6069 2087 6103
rect 16497 6069 16531 6103
rect 19717 6069 19751 6103
rect 1685 5865 1719 5899
rect 4261 5865 4295 5899
rect 5365 5865 5399 5899
rect 6469 5865 6503 5899
rect 7573 5865 7607 5899
rect 16037 5865 16071 5899
rect 21465 5865 21499 5899
rect 29653 5865 29687 5899
rect 32321 5865 32355 5899
rect 21281 5797 21315 5831
rect 4077 5729 4111 5763
rect 5181 5729 5215 5763
rect 6285 5729 6319 5763
rect 7389 5729 7423 5763
rect 28540 5729 28574 5763
rect 32137 5729 32171 5763
rect 21557 5661 21591 5695
rect 28273 5661 28307 5695
rect 21005 5593 21039 5627
rect 15577 5525 15611 5559
rect 1593 5321 1627 5355
rect 15577 5321 15611 5355
rect 21005 5321 21039 5355
rect 21741 5321 21775 5355
rect 28641 5321 28675 5355
rect 32137 5321 32171 5355
rect 21281 5253 21315 5287
rect 1409 5117 1443 5151
rect 4169 5117 4203 5151
rect 2053 5049 2087 5083
rect 15853 5049 15887 5083
rect 16129 5049 16163 5083
rect 5181 4981 5215 5015
rect 6285 4981 6319 5015
rect 7389 4981 7423 5015
rect 15393 4981 15427 5015
rect 16037 4981 16071 5015
rect 28273 4981 28307 5015
rect 1593 4777 1627 4811
rect 15485 4777 15519 4811
rect 16681 4777 16715 4811
rect 16773 4709 16807 4743
rect 1409 4641 1443 4675
rect 16589 4573 16623 4607
rect 16221 4505 16255 4539
rect 16589 4233 16623 4267
rect 16957 4165 16991 4199
rect 16221 4097 16255 4131
rect 1409 4029 1443 4063
rect 2053 3961 2087 3995
rect 1593 3893 1627 3927
rect 9873 3689 9907 3723
rect 8401 3553 8435 3587
rect 9689 3553 9723 3587
rect 1685 3485 1719 3519
rect 8585 3349 8619 3383
rect 1593 3145 1627 3179
rect 8401 3145 8435 3179
rect 9689 3145 9723 3179
rect 27445 3145 27479 3179
rect 2697 3077 2731 3111
rect 1409 2941 1443 2975
rect 2513 2941 2547 2975
rect 3065 2941 3099 2975
rect 26065 2941 26099 2975
rect 26310 2873 26344 2907
rect 2053 2805 2087 2839
rect 25881 2805 25915 2839
rect 2881 2601 2915 2635
rect 4261 2601 4295 2635
rect 26065 2601 26099 2635
rect 1409 2465 1443 2499
rect 1961 2465 1995 2499
rect 2697 2465 2731 2499
rect 4077 2465 4111 2499
rect 18337 2465 18371 2499
rect 18981 2465 19015 2499
rect 1593 2329 1627 2363
rect 3341 2261 3375 2295
rect 4721 2261 4755 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 1762 14152 1768 14204
rect 1820 14192 1826 14204
rect 34514 14192 34520 14204
rect 1820 14164 34520 14192
rect 1820 14152 1826 14164
rect 34514 14152 34520 14164
rect 34572 14152 34578 14204
rect 3326 14084 3332 14136
rect 3384 14124 3390 14136
rect 14090 14124 14096 14136
rect 3384 14096 14096 14124
rect 3384 14084 3390 14096
rect 14090 14084 14096 14096
rect 14148 14084 14154 14136
rect 28902 14084 28908 14136
rect 28960 14124 28966 14136
rect 34882 14124 34888 14136
rect 28960 14096 34888 14124
rect 28960 14084 28966 14096
rect 34882 14084 34888 14096
rect 34940 14084 34946 14136
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 20438 14056 20444 14068
rect 3476 14028 20444 14056
rect 3476 14016 3482 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 27982 14016 27988 14068
rect 28040 14056 28046 14068
rect 34790 14056 34796 14068
rect 28040 14028 34796 14056
rect 28040 14016 28046 14028
rect 34790 14016 34796 14028
rect 34848 14016 34854 14068
rect 3326 13948 3332 14000
rect 3384 13988 3390 14000
rect 34606 13988 34612 14000
rect 3384 13960 34612 13988
rect 3384 13948 3390 13960
rect 34606 13948 34612 13960
rect 34664 13948 34670 14000
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 34698 13920 34704 13932
rect 1636 13892 34704 13920
rect 1636 13880 1642 13892
rect 34698 13880 34704 13892
rect 34756 13880 34762 13932
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5718 13852 5724 13864
rect 4120 13824 5724 13852
rect 4120 13812 4126 13824
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 32306 13812 32312 13864
rect 32364 13852 32370 13864
rect 34514 13852 34520 13864
rect 32364 13824 34520 13852
rect 32364 13812 32370 13824
rect 34514 13812 34520 13824
rect 34572 13812 34578 13864
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9180 12804 12480 12832
rect 9180 12792 9186 12804
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 12452 12764 12480 12804
rect 34698 12764 34704 12776
rect 8720 12736 11836 12764
rect 12452 12736 34704 12764
rect 8720 12724 8726 12736
rect 1946 12656 1952 12708
rect 2004 12696 2010 12708
rect 11808 12696 11836 12736
rect 34698 12724 34704 12736
rect 34756 12724 34762 12776
rect 34514 12696 34520 12708
rect 2004 12668 11744 12696
rect 11808 12668 34520 12696
rect 2004 12656 2010 12668
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 8294 12628 8300 12640
rect 3108 12600 8300 12628
rect 3108 12588 3114 12600
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 11716 12628 11744 12668
rect 34514 12656 34520 12668
rect 34572 12656 34578 12708
rect 34606 12628 34612 12640
rect 11716 12600 34612 12628
rect 34606 12588 34612 12600
rect 34664 12588 34670 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 2314 12424 2320 12436
rect 2275 12396 2320 12424
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 17218 12356 17224 12368
rect 17179 12328 17224 12356
rect 17218 12316 17224 12328
rect 17276 12316 17282 12368
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2498 12288 2504 12300
rect 2179 12260 2504 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12288 17003 12291
rect 17034 12288 17040 12300
rect 16991 12260 17040 12288
rect 16991 12257 17003 12260
rect 16945 12251 17003 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2682 11880 2688 11892
rect 2643 11852 2688 11880
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 14090 11880 14096 11892
rect 14051 11852 14096 11880
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 20438 11880 20444 11892
rect 20399 11852 20444 11880
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1854 11676 1860 11688
rect 1443 11648 1860 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1854 11636 1860 11648
rect 1912 11676 1918 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1912 11648 1961 11676
rect 1912 11636 1918 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 13909 11679 13967 11685
rect 2547 11648 3188 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 3160 11617 3188 11648
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 20257 11679 20315 11685
rect 13955 11648 14596 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 3145 11611 3203 11617
rect 3145 11577 3157 11611
rect 3191 11608 3203 11611
rect 3418 11608 3424 11620
rect 3191 11580 3424 11608
rect 3191 11577 3203 11580
rect 3145 11571 3203 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11540 2467 11543
rect 2498 11540 2504 11552
rect 2455 11512 2504 11540
rect 2455 11509 2467 11512
rect 2409 11503 2467 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 14568 11549 14596 11648
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 20303 11648 20944 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 14553 11543 14611 11549
rect 14553 11509 14565 11543
rect 14599 11540 14611 11543
rect 14642 11540 14648 11552
rect 14599 11512 14648 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 17034 11540 17040 11552
rect 16995 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 20916 11549 20944 11648
rect 20901 11543 20959 11549
rect 20901 11509 20913 11543
rect 20947 11540 20959 11543
rect 21266 11540 21272 11552
rect 20947 11512 21272 11540
rect 20947 11509 20959 11512
rect 20901 11503 20959 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2317 11339 2375 11345
rect 2317 11336 2329 11339
rect 2280 11308 2329 11336
rect 2280 11296 2286 11308
rect 2317 11305 2329 11308
rect 2363 11305 2375 11339
rect 2317 11299 2375 11305
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17479 11339 17537 11345
rect 17479 11336 17491 11339
rect 17092 11308 17491 11336
rect 17092 11296 17098 11308
rect 17479 11305 17491 11308
rect 17525 11305 17537 11339
rect 17479 11299 17537 11305
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 17957 11271 18015 11277
rect 17957 11268 17969 11271
rect 17736 11240 17969 11268
rect 17736 11228 17742 11240
rect 17957 11237 17969 11240
rect 18003 11237 18015 11271
rect 17957 11231 18015 11237
rect 26780 11271 26838 11277
rect 26780 11237 26792 11271
rect 26826 11268 26838 11271
rect 26970 11268 26976 11280
rect 26826 11240 26976 11268
rect 26826 11237 26838 11240
rect 26780 11231 26838 11237
rect 26970 11228 26976 11240
rect 27028 11228 27034 11280
rect 2130 11200 2136 11212
rect 2091 11172 2136 11200
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 18046 11200 18052 11212
rect 17828 11172 18052 11200
rect 17828 11160 17834 11172
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 26513 11203 26571 11209
rect 26513 11169 26525 11203
rect 26559 11200 26571 11203
rect 26602 11200 26608 11212
rect 26559 11172 26608 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 27890 11064 27896 11076
rect 27851 11036 27896 11064
rect 27890 11024 27896 11036
rect 27948 11024 27954 11076
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 3326 10792 3332 10804
rect 3287 10764 3332 10792
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17770 10792 17776 10804
rect 17543 10764 17776 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18012 10764 18245 10792
rect 18012 10752 18018 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 3142 10588 3148 10600
rect 3103 10560 3148 10588
rect 3142 10548 3148 10560
rect 3200 10588 3206 10600
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3200 10560 3709 10588
rect 3200 10548 3206 10560
rect 3697 10557 3709 10560
rect 3743 10557 3755 10591
rect 3697 10551 3755 10557
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17678 10452 17684 10464
rect 17368 10424 17684 10452
rect 17368 10412 17374 10424
rect 17678 10412 17684 10424
rect 17736 10452 17742 10464
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17736 10424 17785 10452
rect 17736 10412 17742 10424
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 17773 10415 17831 10421
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 26970 10452 26976 10464
rect 26931 10424 26976 10452
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1581 10251 1639 10257
rect 1581 10248 1593 10251
rect 1544 10220 1593 10248
rect 1544 10208 1550 10220
rect 1581 10217 1593 10220
rect 1627 10217 1639 10251
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 1581 10211 1639 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 32306 10248 32312 10260
rect 32267 10220 32312 10248
rect 32306 10208 32312 10220
rect 32364 10208 32370 10260
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8202 10112 8208 10124
rect 8159 10084 8208 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 32122 10112 32128 10124
rect 32083 10084 32128 10112
rect 32122 10072 32128 10084
rect 32180 10072 32186 10124
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 18598 9908 18604 9920
rect 18187 9880 18604 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18141 9707 18199 9713
rect 18141 9704 18153 9707
rect 18012 9676 18153 9704
rect 18012 9664 18018 9676
rect 18141 9673 18153 9676
rect 18187 9673 18199 9707
rect 18141 9667 18199 9673
rect 5718 9636 5724 9648
rect 5679 9608 5724 9636
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 7466 9636 7472 9648
rect 7427 9608 7472 9636
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 7926 9568 7932 9580
rect 7300 9540 7932 9568
rect 7300 9509 7328 9540
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 17543 9540 18613 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 18601 9537 18613 9540
rect 18647 9568 18659 9571
rect 18690 9568 18696 9580
rect 18647 9540 18696 9568
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 7285 9503 7343 9509
rect 5583 9472 6224 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 1452 9336 1685 9364
rect 1452 9324 1458 9336
rect 1673 9333 1685 9336
rect 1719 9364 1731 9367
rect 2682 9364 2688 9376
rect 1719 9336 2688 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 6196 9373 6224 9472
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 18598 9432 18604 9444
rect 18559 9404 18604 9432
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 18782 9432 18788 9444
rect 18739 9404 18788 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6822 9364 6828 9376
rect 6227 9336 6828 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 8294 9364 8300 9376
rect 8255 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 17862 9364 17868 9376
rect 17775 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9364 17926 9376
rect 18708 9364 18736 9395
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 32122 9364 32128 9376
rect 17920 9336 18736 9364
rect 32083 9336 32128 9364
rect 17920 9324 17926 9336
rect 32122 9324 32128 9336
rect 32180 9324 32186 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1762 9160 1768 9172
rect 1719 9132 1768 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 21266 9052 21272 9104
rect 21324 9092 21330 9104
rect 21453 9095 21511 9101
rect 21453 9092 21465 9095
rect 21324 9064 21465 9092
rect 21324 9052 21330 9064
rect 21453 9061 21465 9064
rect 21499 9061 21511 9095
rect 21453 9055 21511 9061
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 1489 9027 1547 9033
rect 1489 9024 1501 9027
rect 1452 8996 1501 9024
rect 1452 8984 1458 8996
rect 1489 8993 1501 8996
rect 1535 8993 1547 9027
rect 21542 9024 21548 9036
rect 21503 8996 21548 9024
rect 1489 8987 1547 8993
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 20990 8888 20996 8900
rect 20951 8860 20996 8888
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18506 8820 18512 8832
rect 18187 8792 18512 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1946 8616 1952 8628
rect 1627 8588 1952 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18598 8616 18604 8628
rect 18187 8588 18604 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 21358 8616 21364 8628
rect 21319 8588 21364 8616
rect 21358 8576 21364 8588
rect 21416 8616 21422 8628
rect 30650 8616 30656 8628
rect 21416 8588 21496 8616
rect 30611 8588 30656 8616
rect 21416 8576 21422 8588
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 2317 8551 2375 8557
rect 2317 8548 2329 8551
rect 1452 8520 2329 8548
rect 1452 8508 1458 8520
rect 2317 8517 2329 8520
rect 2363 8517 2375 8551
rect 2317 8511 2375 8517
rect 21468 8489 21496 8588
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 32309 8619 32367 8625
rect 32309 8585 32321 8619
rect 32355 8616 32367 8619
rect 32398 8616 32404 8628
rect 32355 8588 32404 8616
rect 32355 8585 32367 8588
rect 32309 8579 32367 8585
rect 32398 8576 32404 8588
rect 32456 8576 32462 8628
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8449 21511 8483
rect 21453 8443 21511 8449
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1486 8412 1492 8424
rect 1443 8384 1492 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1486 8372 1492 8384
rect 1544 8412 1550 8424
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1544 8384 1961 8412
rect 1544 8372 1550 8384
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 17770 8412 17776 8424
rect 17731 8384 17776 8412
rect 1949 8375 2007 8381
rect 17770 8372 17776 8384
rect 17828 8412 17834 8424
rect 18414 8412 18420 8424
rect 17828 8384 18420 8412
rect 17828 8372 17834 8384
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 19518 8412 19524 8424
rect 18739 8384 19524 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 17494 8344 17500 8356
rect 17407 8316 17500 8344
rect 17494 8304 17500 8316
rect 17552 8344 17558 8356
rect 18708 8344 18736 8375
rect 19518 8372 19524 8384
rect 19576 8412 19582 8424
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 19576 8384 20637 8412
rect 19576 8372 19582 8384
rect 20625 8381 20637 8384
rect 20671 8412 20683 8415
rect 21542 8412 21548 8424
rect 20671 8384 21548 8412
rect 20671 8381 20683 8384
rect 20625 8375 20683 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 28994 8412 29000 8424
rect 28955 8384 29000 8412
rect 28994 8372 29000 8384
rect 29052 8412 29058 8424
rect 29273 8415 29331 8421
rect 29273 8412 29285 8415
rect 29052 8384 29285 8412
rect 29052 8372 29058 8384
rect 29273 8381 29285 8384
rect 29319 8381 29331 8415
rect 29273 8375 29331 8381
rect 29362 8372 29368 8424
rect 29420 8412 29426 8424
rect 29529 8415 29587 8421
rect 29529 8412 29541 8415
rect 29420 8384 29541 8412
rect 29420 8372 29426 8384
rect 29529 8381 29541 8384
rect 29575 8381 29587 8415
rect 29529 8375 29587 8381
rect 32030 8372 32036 8424
rect 32088 8412 32094 8424
rect 32125 8415 32183 8421
rect 32125 8412 32137 8415
rect 32088 8384 32137 8412
rect 32088 8372 32094 8384
rect 32125 8381 32137 8384
rect 32171 8412 32183 8415
rect 32677 8415 32735 8421
rect 32677 8412 32689 8415
rect 32171 8384 32689 8412
rect 32171 8381 32183 8384
rect 32125 8375 32183 8381
rect 32677 8381 32689 8384
rect 32723 8381 32735 8415
rect 32677 8375 32735 8381
rect 17552 8316 18736 8344
rect 20993 8347 21051 8353
rect 17552 8304 17558 8316
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21266 8344 21272 8356
rect 21039 8316 21272 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 18598 8276 18604 8288
rect 18559 8248 18604 8276
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 8662 8072 8668 8084
rect 8623 8044 8668 8072
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9858 8072 9864 8084
rect 9819 8044 9864 8072
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17644 8044 17785 8072
rect 17644 8032 17650 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 29362 8072 29368 8084
rect 29323 8044 29368 8072
rect 17773 8035 17831 8041
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 17862 8004 17868 8016
rect 17823 7976 17868 8004
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 17770 7868 17776 7880
rect 17731 7840 17776 7868
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 1578 7800 1584 7812
rect 1539 7772 1584 7800
rect 1578 7760 1584 7772
rect 1636 7760 1642 7812
rect 17310 7800 17316 7812
rect 17271 7772 17316 7800
rect 17310 7760 17316 7772
rect 17368 7760 17374 7812
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 1854 7528 1860 7540
rect 1452 7500 1860 7528
rect 1452 7488 1458 7500
rect 1854 7488 1860 7500
rect 1912 7528 1918 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1912 7500 1961 7528
rect 1912 7488 1918 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 9122 7528 9128 7540
rect 9083 7500 9128 7528
rect 1949 7491 2007 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17862 7528 17868 7540
rect 17359 7500 17868 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 32306 7528 32312 7540
rect 32267 7500 32312 7528
rect 32306 7488 32312 7500
rect 32364 7488 32370 7540
rect 1581 7463 1639 7469
rect 1581 7429 1593 7463
rect 1627 7460 1639 7463
rect 1670 7460 1676 7472
rect 1627 7432 1676 7460
rect 1627 7429 1639 7432
rect 1581 7423 1639 7429
rect 1670 7420 1676 7432
rect 1728 7420 1734 7472
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1443 7296 2329 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 2317 7293 2329 7296
rect 2363 7324 2375 7327
rect 2406 7324 2412 7336
rect 2363 7296 2412 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 8938 7324 8944 7336
rect 8899 7296 8944 7324
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 17770 7324 17776 7336
rect 16991 7296 17776 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 32122 7324 32128 7336
rect 32083 7296 32128 7324
rect 32122 7284 32128 7296
rect 32180 7324 32186 7336
rect 32677 7327 32735 7333
rect 32677 7324 32689 7327
rect 32180 7296 32689 7324
rect 32180 7284 32186 7296
rect 32677 7293 32689 7296
rect 32723 7293 32735 7327
rect 32677 7287 32735 7293
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 2222 7256 2228 7268
rect 1544 7228 2228 7256
rect 1544 7216 1550 7228
rect 2222 7216 2228 7228
rect 2280 7216 2286 7268
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 2038 7188 2044 7200
rect 1820 7160 2044 7188
rect 1820 7148 1826 7160
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14734 7188 14740 7200
rect 14148 7160 14740 7188
rect 14148 7148 14154 7160
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 17586 7188 17592 7200
rect 16632 7160 17592 7188
rect 16632 7148 16638 7160
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 27430 7148 27436 7200
rect 27488 7188 27494 7200
rect 28074 7188 28080 7200
rect 27488 7160 28080 7188
rect 27488 7148 27494 7160
rect 28074 7148 28080 7160
rect 28132 7148 28138 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2314 6984 2320 6996
rect 2004 6956 2320 6984
rect 2004 6944 2010 6956
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 19429 6919 19487 6925
rect 19429 6885 19441 6919
rect 19475 6885 19487 6919
rect 19429 6879 19487 6885
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6848 1547 6851
rect 2038 6848 2044 6860
rect 1535 6820 2044 6848
rect 1535 6817 1547 6820
rect 1489 6811 1547 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2314 6808 2320 6860
rect 2372 6848 2378 6860
rect 2498 6848 2504 6860
rect 2372 6820 2504 6848
rect 2372 6808 2378 6820
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18932 6820 19257 6848
rect 18932 6808 18938 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19444 6848 19472 6879
rect 19702 6848 19708 6860
rect 19444 6820 19708 6848
rect 19245 6811 19303 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 566 6740 572 6792
rect 624 6780 630 6792
rect 8938 6780 8944 6792
rect 624 6752 8944 6780
rect 624 6740 630 6752
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1946 6712 1952 6724
rect 1719 6684 1952 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18969 6715 19027 6721
rect 18969 6712 18981 6715
rect 18012 6684 18981 6712
rect 18012 6672 18018 6684
rect 18969 6681 18981 6684
rect 19015 6681 19027 6715
rect 18969 6675 19027 6681
rect 20530 6672 20536 6724
rect 20588 6712 20594 6724
rect 21542 6712 21548 6724
rect 20588 6684 21548 6712
rect 20588 6672 20594 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 8386 6644 8392 6656
rect 7524 6616 8392 6644
rect 7524 6604 7530 6616
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 15930 6644 15936 6656
rect 15891 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 16482 6440 16488 6452
rect 16071 6412 16488 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 18874 6440 18880 6452
rect 18835 6412 18880 6440
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 19518 6440 19524 6452
rect 19383 6412 19524 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 32309 6443 32367 6449
rect 32309 6409 32321 6443
rect 32355 6440 32367 6443
rect 32490 6440 32496 6452
rect 32355 6412 32496 6440
rect 32355 6409 32367 6412
rect 32309 6403 32367 6409
rect 32490 6400 32496 6412
rect 32548 6400 32554 6452
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6304 15899 6307
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 15887 6276 16589 6304
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 16577 6273 16589 6276
rect 16623 6304 16635 6307
rect 17494 6304 17500 6316
rect 16623 6276 17500 6304
rect 16623 6273 16635 6276
rect 16577 6267 16635 6273
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1670 6236 1676 6248
rect 1443 6208 1676 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1670 6196 1676 6208
rect 1728 6236 1734 6248
rect 2498 6236 2504 6248
rect 1728 6208 2504 6236
rect 1728 6196 1734 6208
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 32122 6236 32128 6248
rect 32083 6208 32128 6236
rect 32122 6196 32128 6208
rect 32180 6236 32186 6248
rect 32677 6239 32735 6245
rect 32677 6236 32689 6239
rect 32180 6208 32689 6236
rect 32180 6196 32186 6208
rect 32677 6205 32689 6208
rect 32723 6205 32735 6239
rect 32677 6199 32735 6205
rect 15562 6128 15568 6180
rect 15620 6168 15626 6180
rect 15930 6168 15936 6180
rect 15620 6140 15936 6168
rect 15620 6128 15626 6140
rect 15930 6128 15936 6140
rect 15988 6168 15994 6180
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 15988 6140 16313 6168
rect 15988 6128 15994 6140
rect 16301 6137 16313 6140
rect 16347 6137 16359 6171
rect 16301 6131 16359 6137
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 16482 6100 16488 6112
rect 16443 6072 16488 6100
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 19702 6100 19708 6112
rect 19663 6072 19708 6100
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 1670 5896 1676 5908
rect 1631 5868 1676 5896
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 6454 5896 6460 5908
rect 6415 5868 6460 5896
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 7558 5896 7564 5908
rect 7519 5868 7564 5896
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 16482 5896 16488 5908
rect 16071 5868 16488 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 21450 5896 21456 5908
rect 21411 5868 21456 5896
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 29362 5856 29368 5908
rect 29420 5896 29426 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 29420 5868 29653 5896
rect 29420 5856 29426 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 29641 5859 29699 5865
rect 32309 5899 32367 5905
rect 32309 5865 32321 5899
rect 32355 5896 32367 5899
rect 32398 5896 32404 5908
rect 32355 5868 32404 5896
rect 32355 5865 32367 5868
rect 32309 5859 32367 5865
rect 32398 5856 32404 5868
rect 32456 5856 32462 5908
rect 20806 5788 20812 5840
rect 20864 5828 20870 5840
rect 21266 5828 21272 5840
rect 20864 5800 21272 5828
rect 20864 5788 20870 5800
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 28902 5828 28908 5840
rect 28276 5800 28908 5828
rect 4062 5760 4068 5772
rect 4023 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 5166 5760 5172 5772
rect 5127 5732 5172 5760
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 6270 5760 6276 5772
rect 6231 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7340 5732 7389 5760
rect 7340 5720 7346 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 28276 5704 28304 5800
rect 28902 5788 28908 5800
rect 28960 5788 28966 5840
rect 28534 5769 28540 5772
rect 28528 5760 28540 5769
rect 28495 5732 28540 5760
rect 28528 5723 28540 5732
rect 28534 5720 28540 5723
rect 28592 5720 28598 5772
rect 32122 5760 32128 5772
rect 32083 5732 32128 5760
rect 32122 5720 32128 5732
rect 32180 5720 32186 5772
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21726 5692 21732 5704
rect 21591 5664 21732 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 28258 5692 28264 5704
rect 28219 5664 28264 5692
rect 28258 5652 28264 5664
rect 28316 5652 28322 5704
rect 19702 5584 19708 5636
rect 19760 5624 19766 5636
rect 20993 5627 21051 5633
rect 20993 5624 21005 5627
rect 19760 5596 21005 5624
rect 19760 5584 19766 5596
rect 20993 5593 21005 5596
rect 21039 5593 21051 5627
rect 20993 5587 21051 5593
rect 15565 5559 15623 5565
rect 15565 5525 15577 5559
rect 15611 5556 15623 5559
rect 16114 5556 16120 5568
rect 15611 5528 16120 5556
rect 15611 5525 15623 5528
rect 15565 5519 15623 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1762 5352 1768 5364
rect 1627 5324 1768 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 15562 5352 15568 5364
rect 15523 5324 15568 5352
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20864 5324 21005 5352
rect 20864 5312 20870 5324
rect 20993 5321 21005 5324
rect 21039 5352 21051 5355
rect 21450 5352 21456 5364
rect 21039 5324 21456 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 21726 5352 21732 5364
rect 21687 5324 21732 5352
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 28626 5352 28632 5364
rect 28587 5324 28632 5352
rect 28626 5312 28632 5324
rect 28684 5312 28690 5364
rect 32122 5352 32128 5364
rect 32083 5324 32128 5352
rect 32122 5312 32128 5324
rect 32180 5312 32186 5364
rect 21266 5284 21272 5296
rect 21227 5256 21272 5284
rect 21266 5244 21272 5256
rect 21324 5284 21330 5296
rect 21818 5284 21824 5296
rect 21324 5256 21824 5284
rect 21324 5244 21330 5256
rect 21818 5244 21824 5256
rect 21876 5244 21882 5296
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 1412 5080 1440 5111
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4157 5151 4215 5157
rect 4157 5148 4169 5151
rect 4120 5120 4169 5148
rect 4120 5108 4126 5120
rect 4157 5117 4169 5120
rect 4203 5148 4215 5151
rect 4246 5148 4252 5160
rect 4203 5120 4252 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 2041 5083 2099 5089
rect 2041 5080 2053 5083
rect 1412 5052 2053 5080
rect 2041 5049 2053 5052
rect 2087 5080 2099 5083
rect 4338 5080 4344 5092
rect 2087 5052 4344 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 15470 5040 15476 5092
rect 15528 5080 15534 5092
rect 15841 5083 15899 5089
rect 15841 5080 15853 5083
rect 15528 5052 15853 5080
rect 15528 5040 15534 5052
rect 15841 5049 15853 5052
rect 15887 5049 15899 5083
rect 16114 5080 16120 5092
rect 16027 5052 16120 5080
rect 15841 5043 15899 5049
rect 16114 5040 16120 5052
rect 16172 5080 16178 5092
rect 16942 5080 16948 5092
rect 16172 5052 16948 5080
rect 16172 5040 16178 5052
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 5166 5012 5172 5024
rect 4212 4984 5172 5012
rect 4212 4972 4218 4984
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 6270 5012 6276 5024
rect 6231 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 7374 5012 7380 5024
rect 7335 4984 7380 5012
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 15378 5012 15384 5024
rect 15291 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 5012 15442 5024
rect 16022 5012 16028 5024
rect 15436 4984 16028 5012
rect 15436 4972 15442 4984
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 28258 5012 28264 5024
rect 28219 4984 28264 5012
rect 28258 4972 28264 4984
rect 28316 4972 28322 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1544 4780 1593 4808
rect 1544 4768 1550 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 8202 4808 8208 4820
rect 6880 4780 8208 4808
rect 6880 4768 6886 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 16666 4808 16672 4820
rect 16627 4780 16672 4808
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 16942 4740 16948 4752
rect 16807 4712 16948 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 16942 4700 16948 4712
rect 17000 4740 17006 4752
rect 17310 4740 17316 4752
rect 17000 4712 17316 4740
rect 17000 4700 17006 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1670 4672 1676 4684
rect 1443 4644 1676 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 16574 4604 16580 4616
rect 16535 4576 16580 4604
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 16209 4539 16267 4545
rect 16209 4505 16221 4539
rect 16255 4536 16267 4539
rect 16482 4536 16488 4548
rect 16255 4508 16488 4536
rect 16255 4505 16267 4508
rect 16209 4499 16267 4505
rect 16482 4496 16488 4508
rect 16540 4496 16546 4548
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 21358 4468 21364 4480
rect 20772 4440 21364 4468
rect 20772 4428 20778 4440
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 16574 4264 16580 4276
rect 16535 4236 16580 4264
rect 16574 4224 16580 4236
rect 16632 4264 16638 4276
rect 17862 4264 17868 4276
rect 16632 4236 17868 4264
rect 16632 4224 16638 4236
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 16666 4196 16672 4208
rect 16592 4168 16672 4196
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 16209 4131 16267 4137
rect 16209 4128 16221 4131
rect 14148 4100 16221 4128
rect 14148 4088 14154 4100
rect 16209 4097 16221 4100
rect 16255 4128 16267 4131
rect 16592 4128 16620 4168
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 16942 4196 16948 4208
rect 16903 4168 16948 4196
rect 16942 4156 16948 4168
rect 17000 4156 17006 4208
rect 16255 4100 16620 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 1412 3992 1440 4023
rect 2038 3992 2044 4004
rect 1412 3964 2044 3992
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2682 3924 2688 3936
rect 1627 3896 2688 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 27430 3680 27436 3732
rect 27488 3720 27494 3732
rect 28350 3720 28356 3732
rect 27488 3692 28356 3720
rect 27488 3680 27494 3692
rect 28350 3680 28356 3692
rect 28408 3680 28414 3732
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 8570 3380 8576 3392
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 2590 3176 2596 3188
rect 1627 3148 2596 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 8386 3176 8392 3188
rect 8347 3148 8392 3176
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 27433 3179 27491 3185
rect 27433 3145 27445 3179
rect 27479 3176 27491 3179
rect 27522 3176 27528 3188
rect 27479 3148 27528 3176
rect 27479 3145 27491 3148
rect 27433 3139 27491 3145
rect 27522 3136 27528 3148
rect 27580 3136 27586 3188
rect 2682 3108 2688 3120
rect 2643 3080 2688 3108
rect 2682 3068 2688 3080
rect 2740 3068 2746 3120
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2501 2975 2559 2981
rect 1443 2944 2084 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2056 2848 2084 2944
rect 2501 2941 2513 2975
rect 2547 2972 2559 2975
rect 2774 2972 2780 2984
rect 2547 2944 2780 2972
rect 2547 2941 2559 2944
rect 2501 2935 2559 2941
rect 2774 2932 2780 2944
rect 2832 2972 2838 2984
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2832 2944 3065 2972
rect 2832 2932 2838 2944
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 26050 2972 26056 2984
rect 26011 2944 26056 2972
rect 3053 2935 3111 2941
rect 26050 2932 26056 2944
rect 26108 2932 26114 2984
rect 26298 2907 26356 2913
rect 26298 2904 26310 2907
rect 25884 2876 26310 2904
rect 25884 2848 25912 2876
rect 26298 2873 26310 2876
rect 26344 2873 26356 2907
rect 26298 2867 26356 2873
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 25866 2836 25872 2848
rect 25827 2808 25872 2836
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3142 2632 3148 2644
rect 2915 2604 3148 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 4249 2635 4307 2641
rect 4249 2632 4261 2635
rect 3660 2604 4261 2632
rect 3660 2592 3666 2604
rect 4249 2601 4261 2604
rect 4295 2601 4307 2635
rect 26050 2632 26056 2644
rect 26011 2604 26056 2632
rect 4249 2595 4307 2601
rect 26050 2592 26056 2604
rect 26108 2592 26114 2644
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2496 1458 2508
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1452 2468 1961 2496
rect 1452 2456 1458 2468
rect 1949 2465 1961 2468
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 3326 2496 3332 2508
rect 2731 2468 3332 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4706 2496 4712 2508
rect 4111 2468 4712 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18966 2496 18972 2508
rect 18371 2468 18972 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 1578 2360 1584 2372
rect 1539 2332 1584 2360
rect 1578 2320 1584 2332
rect 1636 2320 1642 2372
rect 3326 2292 3332 2304
rect 3287 2264 3332 2292
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 4706 2292 4712 2304
rect 4667 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 18506 2292 18512 2304
rect 18467 2264 18512 2292
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 1768 14152 1820 14204
rect 34520 14152 34572 14204
rect 3332 14084 3384 14136
rect 14096 14084 14148 14136
rect 28908 14084 28960 14136
rect 34888 14084 34940 14136
rect 3424 14016 3476 14068
rect 20444 14016 20496 14068
rect 27988 14016 28040 14068
rect 34796 14016 34848 14068
rect 3332 13948 3384 14000
rect 34612 13948 34664 14000
rect 1584 13880 1636 13932
rect 34704 13880 34756 13932
rect 4068 13812 4120 13864
rect 5724 13812 5776 13864
rect 32312 13812 32364 13864
rect 34520 13812 34572 13864
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 9128 12792 9180 12844
rect 8668 12724 8720 12776
rect 1952 12656 2004 12708
rect 34704 12724 34756 12776
rect 3056 12588 3108 12640
rect 8300 12588 8352 12640
rect 34520 12656 34572 12708
rect 34612 12588 34664 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 2320 12427 2372 12436
rect 2320 12393 2329 12427
rect 2329 12393 2363 12427
rect 2363 12393 2372 12427
rect 2320 12384 2372 12393
rect 17224 12359 17276 12368
rect 17224 12325 17233 12359
rect 17233 12325 17267 12359
rect 17267 12325 17276 12359
rect 17224 12316 17276 12325
rect 2504 12248 2556 12300
rect 17040 12248 17092 12300
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 1860 11636 1912 11688
rect 3424 11568 3476 11620
rect 2504 11500 2556 11552
rect 14648 11500 14700 11552
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 21272 11500 21324 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 2228 11296 2280 11348
rect 17040 11296 17092 11348
rect 17684 11228 17736 11280
rect 26976 11228 27028 11280
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 17776 11160 17828 11212
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 26608 11160 26660 11212
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 27896 11067 27948 11076
rect 27896 11033 27905 11067
rect 27905 11033 27939 11067
rect 27939 11033 27948 11067
rect 27896 11024 27948 11033
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 17776 10752 17828 10804
rect 17960 10752 18012 10804
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 17316 10412 17368 10464
rect 17684 10412 17736 10464
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 26976 10455 27028 10464
rect 26976 10421 26985 10455
rect 26985 10421 27019 10455
rect 27019 10421 27028 10455
rect 26976 10412 27028 10421
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1492 10208 1544 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 32312 10251 32364 10260
rect 32312 10217 32321 10251
rect 32321 10217 32355 10251
rect 32355 10217 32364 10251
rect 32312 10208 32364 10217
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 8208 10072 8260 10124
rect 32128 10115 32180 10124
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 18604 9868 18656 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 17960 9664 18012 9716
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 18696 9528 18748 9580
rect 1400 9324 1452 9376
rect 2688 9324 2740 9376
rect 18604 9435 18656 9444
rect 18604 9401 18613 9435
rect 18613 9401 18647 9435
rect 18647 9401 18656 9435
rect 18604 9392 18656 9401
rect 6828 9324 6880 9376
rect 8300 9367 8352 9376
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 18788 9392 18840 9444
rect 32128 9367 32180 9376
rect 17868 9324 17920 9333
rect 32128 9333 32137 9367
rect 32137 9333 32171 9367
rect 32171 9333 32180 9367
rect 32128 9324 32180 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1768 9120 1820 9172
rect 21272 9052 21324 9104
rect 1400 8984 1452 9036
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 20996 8891 21048 8900
rect 20996 8857 21005 8891
rect 21005 8857 21039 8891
rect 21039 8857 21048 8891
rect 20996 8848 21048 8857
rect 18512 8780 18564 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1952 8576 2004 8628
rect 18604 8576 18656 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 30656 8619 30708 8628
rect 21364 8576 21416 8585
rect 1400 8508 1452 8560
rect 30656 8585 30665 8619
rect 30665 8585 30699 8619
rect 30699 8585 30708 8619
rect 30656 8576 30708 8585
rect 32404 8576 32456 8628
rect 1492 8372 1544 8424
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 18420 8415 18472 8424
rect 17776 8372 17828 8381
rect 18420 8381 18429 8415
rect 18429 8381 18463 8415
rect 18463 8381 18472 8415
rect 18420 8372 18472 8381
rect 17500 8347 17552 8356
rect 17500 8313 17509 8347
rect 17509 8313 17543 8347
rect 17543 8313 17552 8347
rect 19524 8372 19576 8424
rect 21548 8372 21600 8424
rect 29000 8415 29052 8424
rect 29000 8381 29009 8415
rect 29009 8381 29043 8415
rect 29043 8381 29052 8415
rect 29000 8372 29052 8381
rect 29368 8372 29420 8424
rect 32036 8372 32088 8424
rect 17500 8304 17552 8313
rect 21272 8304 21324 8356
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 17592 8032 17644 8084
rect 29368 8075 29420 8084
rect 29368 8041 29377 8075
rect 29377 8041 29411 8075
rect 29411 8041 29420 8075
rect 29368 8032 29420 8041
rect 17868 8007 17920 8016
rect 17868 7973 17877 8007
rect 17877 7973 17911 8007
rect 17911 7973 17920 8007
rect 17868 7964 17920 7973
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 1584 7803 1636 7812
rect 1584 7769 1593 7803
rect 1593 7769 1627 7803
rect 1627 7769 1636 7803
rect 1584 7760 1636 7769
rect 17316 7803 17368 7812
rect 17316 7769 17325 7803
rect 17325 7769 17359 7803
rect 17359 7769 17368 7803
rect 17316 7760 17368 7769
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 1400 7488 1452 7540
rect 1860 7488 1912 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 17868 7488 17920 7540
rect 32312 7531 32364 7540
rect 32312 7497 32321 7531
rect 32321 7497 32355 7531
rect 32355 7497 32364 7531
rect 32312 7488 32364 7497
rect 1676 7420 1728 7472
rect 2412 7284 2464 7336
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 17776 7284 17828 7336
rect 32128 7327 32180 7336
rect 32128 7293 32137 7327
rect 32137 7293 32171 7327
rect 32171 7293 32180 7327
rect 32128 7284 32180 7293
rect 1492 7216 1544 7268
rect 2228 7216 2280 7268
rect 1768 7148 1820 7200
rect 2044 7148 2096 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 14096 7148 14148 7200
rect 14740 7148 14792 7200
rect 16580 7148 16632 7200
rect 17592 7191 17644 7200
rect 17592 7157 17601 7191
rect 17601 7157 17635 7191
rect 17635 7157 17644 7191
rect 17592 7148 17644 7157
rect 27436 7148 27488 7200
rect 28080 7148 28132 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1952 6944 2004 6996
rect 2320 6944 2372 6996
rect 2044 6808 2096 6860
rect 2320 6808 2372 6860
rect 2504 6808 2556 6860
rect 18880 6808 18932 6860
rect 19708 6808 19760 6860
rect 572 6740 624 6792
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 1952 6672 2004 6724
rect 17960 6672 18012 6724
rect 20536 6672 20588 6724
rect 21548 6672 21600 6724
rect 7472 6604 7524 6656
rect 8392 6604 8444 6656
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1676 6400 1728 6452
rect 16488 6400 16540 6452
rect 18880 6443 18932 6452
rect 18880 6409 18889 6443
rect 18889 6409 18923 6443
rect 18923 6409 18932 6443
rect 18880 6400 18932 6409
rect 19524 6400 19576 6452
rect 32496 6400 32548 6452
rect 17500 6264 17552 6316
rect 1676 6196 1728 6248
rect 2504 6196 2556 6248
rect 32128 6239 32180 6248
rect 32128 6205 32137 6239
rect 32137 6205 32171 6239
rect 32171 6205 32180 6239
rect 32128 6196 32180 6205
rect 15568 6128 15620 6180
rect 15936 6128 15988 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 16488 6103 16540 6112
rect 16488 6069 16497 6103
rect 16497 6069 16531 6103
rect 16531 6069 16540 6103
rect 16488 6060 16540 6069
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 1676 5899 1728 5908
rect 1676 5865 1685 5899
rect 1685 5865 1719 5899
rect 1719 5865 1728 5899
rect 1676 5856 1728 5865
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 6460 5899 6512 5908
rect 6460 5865 6469 5899
rect 6469 5865 6503 5899
rect 6503 5865 6512 5899
rect 6460 5856 6512 5865
rect 7564 5899 7616 5908
rect 7564 5865 7573 5899
rect 7573 5865 7607 5899
rect 7607 5865 7616 5899
rect 7564 5856 7616 5865
rect 16488 5856 16540 5908
rect 21456 5899 21508 5908
rect 21456 5865 21465 5899
rect 21465 5865 21499 5899
rect 21499 5865 21508 5899
rect 21456 5856 21508 5865
rect 29368 5856 29420 5908
rect 32404 5856 32456 5908
rect 20812 5788 20864 5840
rect 21272 5831 21324 5840
rect 21272 5797 21281 5831
rect 21281 5797 21315 5831
rect 21315 5797 21324 5831
rect 21272 5788 21324 5797
rect 4068 5763 4120 5772
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 7288 5720 7340 5772
rect 28908 5788 28960 5840
rect 28540 5763 28592 5772
rect 28540 5729 28574 5763
rect 28574 5729 28592 5763
rect 28540 5720 28592 5729
rect 32128 5763 32180 5772
rect 32128 5729 32137 5763
rect 32137 5729 32171 5763
rect 32171 5729 32180 5763
rect 32128 5720 32180 5729
rect 21732 5652 21784 5704
rect 28264 5695 28316 5704
rect 28264 5661 28273 5695
rect 28273 5661 28307 5695
rect 28307 5661 28316 5695
rect 28264 5652 28316 5661
rect 19708 5584 19760 5636
rect 16120 5516 16172 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1768 5312 1820 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 20812 5312 20864 5364
rect 21456 5312 21508 5364
rect 21732 5355 21784 5364
rect 21732 5321 21741 5355
rect 21741 5321 21775 5355
rect 21775 5321 21784 5355
rect 21732 5312 21784 5321
rect 28632 5355 28684 5364
rect 28632 5321 28641 5355
rect 28641 5321 28675 5355
rect 28675 5321 28684 5355
rect 28632 5312 28684 5321
rect 32128 5355 32180 5364
rect 32128 5321 32137 5355
rect 32137 5321 32171 5355
rect 32171 5321 32180 5355
rect 32128 5312 32180 5321
rect 21272 5287 21324 5296
rect 21272 5253 21281 5287
rect 21281 5253 21315 5287
rect 21315 5253 21324 5287
rect 21272 5244 21324 5253
rect 21824 5244 21876 5296
rect 4068 5108 4120 5160
rect 4252 5108 4304 5160
rect 4344 5040 4396 5092
rect 15476 5040 15528 5092
rect 16120 5083 16172 5092
rect 16120 5049 16129 5083
rect 16129 5049 16163 5083
rect 16163 5049 16172 5083
rect 16120 5040 16172 5049
rect 16948 5040 17000 5092
rect 4160 4972 4212 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 16028 5015 16080 5024
rect 15384 4972 15436 4981
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 28264 5015 28316 5024
rect 28264 4981 28273 5015
rect 28273 4981 28307 5015
rect 28307 4981 28316 5015
rect 28264 4972 28316 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1492 4768 1544 4820
rect 6828 4768 6880 4820
rect 8208 4768 8260 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 16948 4700 17000 4752
rect 17316 4700 17368 4752
rect 1676 4632 1728 4684
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 16488 4496 16540 4548
rect 20720 4428 20772 4480
rect 21364 4428 21416 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 16580 4267 16632 4276
rect 16580 4233 16589 4267
rect 16589 4233 16623 4267
rect 16623 4233 16632 4267
rect 16580 4224 16632 4233
rect 17868 4224 17920 4276
rect 14096 4088 14148 4140
rect 16672 4156 16724 4208
rect 16948 4199 17000 4208
rect 16948 4165 16957 4199
rect 16957 4165 16991 4199
rect 16991 4165 17000 4199
rect 16948 4156 17000 4165
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 2688 3884 2740 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 27436 3680 27488 3732
rect 28356 3680 28408 3732
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2596 3136 2648 3188
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 27528 3136 27580 3188
rect 2688 3111 2740 3120
rect 2688 3077 2697 3111
rect 2697 3077 2731 3111
rect 2731 3077 2740 3111
rect 2688 3068 2740 3077
rect 2780 2932 2832 2984
rect 26056 2975 26108 2984
rect 26056 2941 26065 2975
rect 26065 2941 26099 2975
rect 26099 2941 26108 2975
rect 26056 2932 26108 2941
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 25872 2839 25924 2848
rect 25872 2805 25881 2839
rect 25881 2805 25915 2839
rect 25915 2805 25924 2839
rect 25872 2796 25924 2805
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 3148 2592 3200 2644
rect 3608 2592 3660 2644
rect 26056 2635 26108 2644
rect 26056 2601 26065 2635
rect 26065 2601 26099 2635
rect 26099 2601 26108 2635
rect 26056 2592 26108 2601
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 3332 2456 3384 2508
rect 4712 2456 4764 2508
rect 18972 2499 19024 2508
rect 18972 2465 18981 2499
rect 18981 2465 19015 2499
rect 19015 2465 19024 2499
rect 18972 2456 19024 2465
rect 1584 2363 1636 2372
rect 1584 2329 1593 2363
rect 1593 2329 1627 2363
rect 1627 2329 1636 2363
rect 1584 2320 1636 2329
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 18512 2295 18564 2304
rect 18512 2261 18521 2295
rect 18521 2261 18555 2295
rect 18555 2261 18564 2295
rect 18512 2252 18564 2261
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 2686 15872 2742 15881
rect 2686 15807 2742 15816
rect 2318 15464 2374 15473
rect 2318 15399 2374 15408
rect 2226 15056 2282 15065
rect 2226 14991 2282 15000
rect 1768 14204 1820 14210
rect 1768 14146 1820 14152
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1490 13016 1546 13025
rect 1490 12951 1546 12960
rect 1504 10266 1532 12951
rect 1596 11898 1624 13874
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 9382 1440 10066
rect 1674 9752 1730 9761
rect 1674 9687 1730 9696
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8566 1440 8978
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1412 8242 1440 8502
rect 1492 8424 1544 8430
rect 1492 8366 1544 8372
rect 1320 8214 1440 8242
rect 1320 7041 1348 8214
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7546 1440 7890
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1504 7426 1532 8366
rect 1582 7848 1638 7857
rect 1582 7783 1584 7792
rect 1636 7783 1638 7792
rect 1584 7754 1636 7760
rect 1688 7478 1716 9687
rect 1780 9178 1808 14146
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1412 7398 1532 7426
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1306 7032 1362 7041
rect 1306 6967 1362 6976
rect 572 6792 624 6798
rect 572 6734 624 6740
rect 584 5817 612 6734
rect 1412 6225 1440 7398
rect 1780 7290 1808 8871
rect 1872 7993 1900 11630
rect 1964 8634 1992 12650
rect 2042 11792 2098 11801
rect 2042 11727 2098 11736
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1858 7984 1914 7993
rect 1858 7919 1914 7928
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1688 7262 1808 7290
rect 1398 6216 1454 6225
rect 1398 6151 1454 6160
rect 570 5808 626 5817
rect 570 5743 626 5752
rect 1504 4826 1532 7210
rect 1688 6458 1716 7262
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5914 1716 6190
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1780 5370 1808 7142
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1872 5001 1900 7482
rect 2056 7206 2084 11727
rect 2240 11354 2268 14991
rect 2332 12442 2360 15399
rect 2410 12608 2466 12617
rect 2410 12543 2466 12552
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2226 11248 2282 11257
rect 2136 11212 2188 11218
rect 2226 11183 2282 11192
rect 2136 11154 2188 11160
rect 2148 10470 2176 11154
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1964 6730 1992 6938
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 2056 6118 2084 6802
rect 2148 6361 2176 10406
rect 2240 7274 2268 11183
rect 2424 7426 2452 12543
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11558 2544 12242
rect 2700 11898 2728 15807
rect 19982 15520 20038 16000
rect 34886 15872 34942 15881
rect 34886 15807 34942 15816
rect 3422 14648 3478 14657
rect 3422 14583 3478 14592
rect 3330 14240 3386 14249
rect 3330 14175 3386 14184
rect 3344 14142 3372 14175
rect 3332 14136 3384 14142
rect 3332 14078 3384 14084
rect 3436 14074 3464 14583
rect 14096 14136 14148 14142
rect 14096 14078 14148 14084
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3054 13424 3110 13433
rect 3054 13359 3110 13368
rect 3068 12646 3096 13359
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2332 7398 2452 7426
rect 2228 7268 2280 7274
rect 2228 7210 2280 7216
rect 2332 7002 2360 7398
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2134 6352 2190 6361
rect 2134 6287 2190 6296
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1858 4992 1914 5001
rect 1858 4927 1914 4936
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 2056 4729 2084 6054
rect 2042 4720 2098 4729
rect 1676 4684 1728 4690
rect 2042 4655 2098 4664
rect 1676 4626 1728 4632
rect 1688 3534 1716 4626
rect 2332 4457 2360 6802
rect 2424 6089 2452 7278
rect 2516 7177 2544 11494
rect 2870 10976 2926 10985
rect 2870 10911 2926 10920
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2502 7168 2558 7177
rect 2502 7103 2558 7112
rect 2700 7018 2728 9318
rect 2516 6990 2728 7018
rect 2516 6866 2544 6990
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2516 6254 2544 6695
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2410 6080 2466 6089
rect 2410 6015 2466 6024
rect 2792 5930 2820 10503
rect 2608 5902 2820 5930
rect 2318 4448 2374 4457
rect 2318 4383 2374 4392
rect 2042 4040 2098 4049
rect 2042 3975 2044 3984
rect 2096 3975 2098 3984
rect 2044 3946 2096 3952
rect 1676 3528 1728 3534
rect 1674 3496 1676 3505
rect 1728 3496 1730 3505
rect 1674 3431 1730 3440
rect 2608 3194 2636 5902
rect 2884 5794 2912 10911
rect 3344 10810 3372 13942
rect 4068 13864 4120 13870
rect 4066 13832 4068 13841
rect 5724 13864 5776 13870
rect 4120 13832 4122 13841
rect 5724 13806 5776 13812
rect 4066 13767 4122 13776
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3160 7449 3188 10542
rect 3238 9344 3294 9353
rect 3238 9279 3294 9288
rect 3146 7440 3202 7449
rect 3146 7375 3202 7384
rect 3252 7324 3280 9279
rect 3436 7449 3464 11562
rect 3698 10160 3754 10169
rect 3698 10095 3754 10104
rect 3606 8528 3662 8537
rect 3606 8463 3662 8472
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 2700 5766 2912 5794
rect 3160 7296 3280 7324
rect 2700 3942 2728 5766
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2688 3120 2740 3126
rect 2686 3088 2688 3097
rect 2740 3088 2742 3097
rect 2686 3023 2742 3032
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 1329 1440 2450
rect 1582 2408 1638 2417
rect 1582 2343 1584 2352
rect 1636 2343 1638 2352
rect 1584 2314 1636 2320
rect 2056 1465 2084 2790
rect 2042 1456 2098 1465
rect 2042 1391 2098 1400
rect 1398 1320 1454 1329
rect 1398 1255 1454 1264
rect 2792 513 2820 2926
rect 3160 2650 3188 7296
rect 3238 5128 3294 5137
rect 3238 5063 3294 5072
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3252 921 3280 5063
rect 3422 3904 3478 3913
rect 3422 3839 3478 3848
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3344 2310 3372 2450
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3238 912 3294 921
rect 3238 847 3294 856
rect 2778 504 2834 513
rect 2778 439 2834 448
rect 3344 105 3372 2246
rect 3436 241 3464 3839
rect 3620 2650 3648 8463
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3712 1873 3740 10095
rect 4080 9625 4108 12135
rect 5736 9654 5764 13806
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 8312 10266 8340 12582
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 10010 8248 10066
rect 8220 9982 8340 10010
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 5724 9648 5776 9654
rect 4066 9616 4122 9625
rect 7472 9648 7524 9654
rect 5724 9590 5776 9596
rect 7470 9616 7472 9625
rect 7524 9616 7526 9625
rect 4066 9551 4122 9560
rect 7470 9551 7526 9560
rect 7930 9616 7986 9625
rect 7930 9551 7932 9560
rect 7984 9551 7986 9560
rect 7932 9522 7984 9528
rect 8312 9382 8340 9982
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 4066 8392 4122 8401
rect 4066 8327 4122 8336
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3790 6488 3846 6497
rect 3790 6423 3846 6432
rect 3804 4185 3832 6423
rect 3988 5409 4016 6831
rect 4080 6633 4108 8327
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 4264 5914 4292 8191
rect 6458 6216 6514 6225
rect 6458 6151 6514 6160
rect 6472 5914 6500 6151
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 5368 5817 5396 5850
rect 5354 5808 5410 5817
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 5172 5772 5224 5778
rect 5354 5743 5410 5752
rect 6276 5772 6328 5778
rect 5172 5714 5224 5720
rect 6276 5714 6328 5720
rect 3974 5400 4030 5409
rect 3974 5335 4030 5344
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3896 4593 3924 5199
rect 4080 5166 4108 5714
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4160 5024 4212 5030
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 4080 4972 4160 4978
rect 4080 4966 4212 4972
rect 4080 4950 4200 4966
rect 3882 4584 3938 4593
rect 3882 4519 3938 4528
rect 3882 4312 3938 4321
rect 3882 4247 3938 4256
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 3896 2961 3924 4247
rect 3988 3369 4016 4927
rect 4080 3777 4108 4950
rect 4264 4865 4292 5102
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4250 4856 4306 4865
rect 4250 4791 4306 4800
rect 4066 3768 4122 3777
rect 4066 3703 4122 3712
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 4356 2961 4384 5034
rect 5184 5030 5212 5714
rect 6288 5030 6316 5714
rect 5172 5024 5224 5030
rect 6276 5024 6328 5030
rect 5172 4966 5224 4972
rect 6274 4992 6276 5001
rect 6328 4992 6330 5001
rect 6274 4927 6330 4936
rect 6840 4826 6868 9318
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6497 7512 6598
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7470 6488 7526 6497
rect 7622 6480 7918 6500
rect 7470 6423 7526 6432
rect 7378 6352 7434 6361
rect 7378 6287 7434 6296
rect 7562 6352 7618 6361
rect 7562 6287 7618 6296
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7300 5522 7328 5714
rect 7392 5681 7420 6287
rect 7576 5914 7604 6287
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7378 5672 7434 5681
rect 7378 5607 7434 5616
rect 7300 5494 7420 5522
rect 7392 5030 7420 5494
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8312 5409 8340 9318
rect 8680 8090 8708 12718
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8496 7206 8524 7890
rect 9140 7546 9168 12786
rect 14108 11898 14136 14078
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 17224 12368 17276 12374
rect 17222 12336 17224 12345
rect 19996 12345 20024 15520
rect 34794 15464 34850 15473
rect 34794 15399 34850 15408
rect 34702 15056 34758 15065
rect 34702 14991 34758 15000
rect 34610 14648 34666 14657
rect 34610 14583 34666 14592
rect 34518 14240 34574 14249
rect 34518 14175 34520 14184
rect 34572 14175 34574 14184
rect 34520 14146 34572 14152
rect 28908 14136 28960 14142
rect 28908 14078 28960 14084
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 17276 12336 17278 12345
rect 17040 12300 17092 12306
rect 17222 12271 17278 12280
rect 19982 12336 20038 12345
rect 19982 12271 20038 12280
rect 17040 12242 17092 12248
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 17052 11558 17080 12242
rect 20456 11898 20484 14010
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9876 7993 9904 8026
rect 9862 7984 9918 7993
rect 9680 7948 9732 7954
rect 9862 7919 9918 7928
rect 9680 7890 9732 7896
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8496 6905 8524 7142
rect 8482 6896 8538 6905
rect 8482 6831 8538 6840
rect 8956 6798 8984 7278
rect 9692 7206 9720 7890
rect 9680 7200 9732 7206
rect 14096 7200 14148 7206
rect 9680 7142 9732 7148
rect 14094 7168 14096 7177
rect 14148 7168 14150 7177
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8392 6656 8444 6662
rect 8390 6624 8392 6633
rect 8444 6624 8446 6633
rect 8390 6559 8446 6568
rect 8298 5400 8354 5409
rect 8298 5335 8354 5344
rect 9692 5273 9720 7142
rect 14094 7103 14150 7112
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14094 6896 14150 6905
rect 14094 6831 14150 6840
rect 14108 6089 14136 6831
rect 14660 6769 14688 11494
rect 17052 11354 17080 11494
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 18050 11248 18106 11257
rect 17696 10470 17724 11222
rect 17776 11212 17828 11218
rect 18050 11183 18052 11192
rect 17776 11154 17828 11160
rect 18104 11183 18106 11192
rect 18052 11154 18104 11160
rect 17788 10810 17816 11154
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10826 17908 11086
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 17880 10810 18000 10826
rect 17776 10804 17828 10810
rect 17880 10804 18012 10810
rect 17880 10798 17960 10804
rect 17776 10746 17828 10752
rect 17960 10746 18012 10752
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17328 7818 17356 10406
rect 17972 9722 18000 10746
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 8424 17828 8430
rect 17774 8392 17776 8401
rect 17828 8392 17830 8401
rect 17500 8356 17552 8362
rect 17774 8327 17830 8336
rect 17500 8298 17552 8304
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 14740 7200 14792 7206
rect 14738 7168 14740 7177
rect 16580 7200 16632 7206
rect 14792 7168 14794 7177
rect 14738 7103 14794 7112
rect 16500 7148 16580 7154
rect 16500 7142 16632 7148
rect 16500 7126 16620 7142
rect 14646 6760 14702 6769
rect 14646 6695 14702 6704
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15474 6488 15530 6497
rect 15474 6423 15530 6432
rect 14094 6080 14150 6089
rect 14094 6015 14150 6024
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 14094 5264 14150 5273
rect 14094 5199 14150 5208
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 7392 4321 7420 4966
rect 14108 4865 14136 5199
rect 15382 5128 15438 5137
rect 15488 5098 15516 6423
rect 15948 6186 15976 6598
rect 16026 6488 16082 6497
rect 16500 6458 16528 7126
rect 16026 6423 16082 6432
rect 16488 6452 16540 6458
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15580 5370 15608 6122
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15382 5063 15438 5072
rect 15476 5092 15528 5098
rect 15396 5030 15424 5063
rect 15476 5034 15528 5040
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 8022 4856 8078 4865
rect 8022 4791 8078 4800
rect 8206 4856 8262 4865
rect 8206 4791 8208 4800
rect 7470 4720 7526 4729
rect 7470 4655 7526 4664
rect 7378 4312 7434 4321
rect 7378 4247 7434 4256
rect 7484 4185 7512 4655
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8036 4321 8064 4791
rect 8260 4791 8262 4800
rect 14094 4856 14150 4865
rect 14289 4848 14585 4868
rect 15488 4826 15516 5034
rect 16040 5030 16068 6423
rect 16488 6394 16540 6400
rect 17512 6322 17540 8298
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17604 7206 17632 8026
rect 17880 8022 17908 9318
rect 18418 8936 18474 8945
rect 18418 8871 18474 8880
rect 18432 8430 18460 8871
rect 18524 8838 18552 9551
rect 18616 9450 18644 9862
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8514 18552 8774
rect 18616 8634 18644 9386
rect 18708 9217 18736 9522
rect 18786 9480 18842 9489
rect 18786 9415 18788 9424
rect 18840 9415 18842 9424
rect 18788 9386 18840 9392
rect 18694 9208 18750 9217
rect 18694 9143 18750 9152
rect 20994 9208 21050 9217
rect 20994 9143 21050 9152
rect 21008 8906 21036 9143
rect 21284 9110 21312 11494
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 26976 11280 27028 11286
rect 26976 11222 27028 11228
rect 27894 11248 27950 11257
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26620 10470 26648 11154
rect 26988 10470 27016 11222
rect 28000 11234 28028 14010
rect 27950 11206 28028 11234
rect 27894 11183 27950 11192
rect 27908 11082 27936 11183
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 26620 10169 26648 10406
rect 26606 10160 26662 10169
rect 26606 10095 26662 10104
rect 26988 9489 27016 10406
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 28920 10169 28948 14078
rect 34624 14006 34652 14583
rect 34612 14000 34664 14006
rect 34518 13968 34574 13977
rect 34612 13942 34664 13948
rect 34716 13938 34744 14991
rect 34808 14074 34836 15399
rect 34900 14142 34928 15807
rect 34888 14136 34940 14142
rect 34888 14078 34940 14084
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34518 13903 34574 13912
rect 34704 13932 34756 13938
rect 34532 13870 34560 13903
rect 34704 13874 34756 13880
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 32324 10266 32352 13806
rect 34610 13560 34666 13569
rect 34610 13495 34666 13504
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34518 12744 34574 12753
rect 34518 12679 34520 12688
rect 34572 12679 34574 12688
rect 34520 12650 34572 12656
rect 34624 12646 34652 13495
rect 34702 13152 34758 13161
rect 34702 13087 34758 13096
rect 34716 12782 34744 13087
rect 34704 12776 34756 12782
rect 34704 12718 34756 12724
rect 34612 12640 34664 12646
rect 34612 12582 34664 12588
rect 34794 12336 34850 12345
rect 34794 12271 34850 12280
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 28906 10160 28962 10169
rect 28906 10095 28962 10104
rect 32128 10124 32180 10130
rect 26974 9480 27030 9489
rect 26974 9415 27030 9424
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21546 9072 21602 9081
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18524 8486 18644 8514
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18616 8294 18644 8486
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 7342 17816 7822
rect 17880 7546 17908 7958
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17776 7336 17828 7342
rect 17828 7284 18000 7290
rect 17776 7278 18000 7284
rect 17788 7262 18000 7278
rect 17788 7213 17816 7262
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17972 6730 18000 7262
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17590 6488 17646 6497
rect 17590 6423 17646 6432
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17604 6225 17632 6423
rect 17314 6216 17370 6225
rect 17314 6151 17370 6160
rect 17590 6216 17646 6225
rect 17590 6151 17646 6160
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 5914 16528 6054
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16132 5098 16160 5510
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 14094 4791 14150 4800
rect 15476 4820 15528 4826
rect 8208 4762 8260 4768
rect 15476 4762 15528 4768
rect 8022 4312 8078 4321
rect 8022 4247 8078 4256
rect 7470 4176 7526 4185
rect 7470 4111 7526 4120
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3913 14136 4082
rect 14094 3904 14150 3913
rect 14094 3839 14150 3848
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9876 3641 9904 3674
rect 9862 3632 9918 3641
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 9680 3596 9732 3602
rect 9862 3567 9918 3576
rect 9680 3538 9732 3544
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8404 3194 8432 3538
rect 8576 3392 8628 3398
rect 8574 3360 8576 3369
rect 8628 3360 8630 3369
rect 8574 3295 8630 3304
rect 9692 3194 9720 3538
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 3882 2952 3938 2961
rect 3882 2887 3938 2896
rect 4342 2952 4398 2961
rect 4342 2887 4398 2896
rect 8404 2553 8432 3130
rect 9692 2689 9720 3130
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 9678 2680 9734 2689
rect 14289 2672 14585 2692
rect 9678 2615 9734 2624
rect 7470 2544 7526 2553
rect 4712 2508 4764 2514
rect 7470 2479 7526 2488
rect 8390 2544 8446 2553
rect 8390 2479 8446 2488
rect 4712 2450 4764 2456
rect 4724 2310 4752 2450
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3698 1864 3754 1873
rect 3698 1799 3754 1808
rect 4724 241 4752 2246
rect 7484 2145 7512 2479
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7470 2136 7526 2145
rect 7622 2128 7918 2148
rect 7470 2071 7526 2080
rect 15488 377 15516 4762
rect 16500 4554 16528 5850
rect 17328 5817 17356 6151
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 17314 5264 17370 5273
rect 17314 5199 17370 5208
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16670 4992 16726 5001
rect 16670 4927 16726 4936
rect 16684 4826 16712 4927
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16592 4321 16620 4558
rect 16578 4312 16634 4321
rect 16578 4247 16580 4256
rect 16632 4247 16634 4256
rect 16580 4218 16632 4224
rect 16684 4214 16712 4762
rect 16960 4758 16988 5034
rect 17328 4758 17356 5199
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 16960 4214 16988 4694
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 17222 3768 17278 3777
rect 17222 3703 17278 3712
rect 17236 3369 17264 3703
rect 17222 3360 17278 3369
rect 17222 3295 17278 3304
rect 17880 513 17908 4218
rect 18616 3913 18644 8230
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18892 6633 18920 6802
rect 19536 6798 19564 8366
rect 21284 8362 21312 9046
rect 21546 9007 21548 9016
rect 21600 9007 21602 9016
rect 21548 8978 21600 8984
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21376 8634 21404 8910
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21560 8430 21588 8978
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 28920 8412 28948 10095
rect 32128 10066 32180 10072
rect 30654 9480 30710 9489
rect 30654 9415 30710 9424
rect 29366 9072 29422 9081
rect 29366 9007 29422 9016
rect 29380 8430 29408 9007
rect 30668 8634 30696 9415
rect 32140 9382 32168 10066
rect 32402 10024 32458 10033
rect 32402 9959 32458 9968
rect 32128 9376 32180 9382
rect 32128 9318 32180 9324
rect 32310 9344 32366 9353
rect 32140 8945 32168 9318
rect 32310 9279 32366 9288
rect 32126 8936 32182 8945
rect 32126 8871 32182 8880
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 29000 8424 29052 8430
rect 28920 8384 29000 8412
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 6905 21312 8298
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28078 8120 28134 8129
rect 28078 8055 28134 8064
rect 28092 7857 28120 8055
rect 28078 7848 28134 7857
rect 28078 7783 28134 7792
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 20810 6896 20866 6905
rect 19708 6860 19760 6866
rect 20810 6831 20866 6840
rect 21270 6896 21326 6905
rect 21270 6831 21326 6840
rect 19708 6802 19760 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 18878 6624 18934 6633
rect 18878 6559 18934 6568
rect 18892 6458 18920 6559
rect 19536 6458 19564 6734
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19720 6118 19748 6802
rect 20534 6760 20590 6769
rect 20534 6695 20536 6704
rect 20588 6695 20590 6704
rect 20536 6666 20588 6672
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19720 5642 19748 6054
rect 20824 5846 20852 6831
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21468 5914 21496 7511
rect 27436 7200 27488 7206
rect 27434 7168 27436 7177
rect 28080 7200 28132 7206
rect 27488 7168 27490 7177
rect 28078 7168 28080 7177
rect 28132 7168 28134 7177
rect 27434 7103 27490 7112
rect 27622 7100 27918 7120
rect 28078 7103 28134 7112
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 21546 6760 21602 6769
rect 21546 6695 21548 6704
rect 21600 6695 21602 6704
rect 28170 6760 28226 6769
rect 28170 6695 28226 6704
rect 21548 6666 21600 6672
rect 26790 6488 26846 6497
rect 26790 6423 26846 6432
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20720 4480 20772 4486
rect 20718 4448 20720 4457
rect 20772 4448 20774 4457
rect 20718 4383 20774 4392
rect 18602 3904 18658 3913
rect 18602 3839 18658 3848
rect 19982 2816 20038 2825
rect 19982 2751 20038 2760
rect 18970 2544 19026 2553
rect 18970 2479 18972 2488
rect 19024 2479 19026 2488
rect 18972 2450 19024 2456
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18524 1873 18552 2246
rect 18510 1864 18566 1873
rect 18510 1799 18566 1808
rect 17866 504 17922 513
rect 19996 480 20024 2751
rect 20824 2009 20852 5306
rect 21284 5302 21312 5782
rect 21468 5370 21496 5850
rect 26804 5817 26832 6423
rect 28078 6352 28134 6361
rect 28078 6287 28134 6296
rect 28092 6089 28120 6287
rect 28078 6080 28134 6089
rect 27622 6012 27918 6032
rect 28078 6015 28134 6024
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28184 5953 28212 6695
rect 28170 5944 28226 5953
rect 28170 5879 28226 5888
rect 28920 5846 28948 8384
rect 29000 8366 29052 8372
rect 29368 8424 29420 8430
rect 29368 8366 29420 8372
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 29380 8090 29408 8366
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29380 5914 29408 8026
rect 32048 6633 32076 8366
rect 32126 7576 32182 7585
rect 32324 7546 32352 9279
rect 32416 8634 32444 9959
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34610 8936 34666 8945
rect 34610 8871 34666 8880
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32494 8256 32550 8265
rect 32494 8191 32550 8200
rect 32402 7848 32458 7857
rect 32402 7783 32458 7792
rect 32126 7511 32182 7520
rect 32312 7540 32364 7546
rect 32140 7342 32168 7511
rect 32312 7482 32364 7488
rect 32128 7336 32180 7342
rect 32128 7278 32180 7284
rect 32034 6624 32090 6633
rect 32034 6559 32090 6568
rect 32128 6248 32180 6254
rect 32126 6216 32128 6225
rect 32180 6216 32182 6225
rect 32126 6151 32182 6160
rect 32416 5914 32444 7783
rect 32508 6458 32536 8191
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 32496 6452 32548 6458
rect 32496 6394 32548 6400
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 32404 5908 32456 5914
rect 32404 5850 32456 5856
rect 28908 5840 28960 5846
rect 26790 5808 26846 5817
rect 28908 5782 28960 5788
rect 26790 5743 26846 5752
rect 28540 5772 28592 5778
rect 28540 5714 28592 5720
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 21744 5409 21772 5646
rect 27526 5536 27582 5545
rect 27526 5471 27582 5480
rect 21730 5400 21786 5409
rect 21456 5364 21508 5370
rect 21730 5335 21732 5344
rect 21456 5306 21508 5312
rect 21784 5335 21786 5344
rect 21732 5306 21784 5312
rect 21272 5296 21324 5302
rect 21824 5296 21876 5302
rect 21272 5238 21324 5244
rect 21546 5264 21602 5273
rect 21824 5238 21876 5244
rect 27066 5264 27122 5273
rect 21546 5199 21602 5208
rect 21560 5001 21588 5199
rect 21546 4992 21602 5001
rect 21546 4927 21602 4936
rect 21364 4480 21416 4486
rect 21362 4448 21364 4457
rect 21416 4448 21418 4457
rect 20956 4380 21252 4400
rect 21362 4383 21418 4392
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21546 4040 21602 4049
rect 21546 3975 21602 3984
rect 21560 3641 21588 3975
rect 21362 3632 21418 3641
rect 21362 3567 21418 3576
rect 21546 3632 21602 3641
rect 21546 3567 21602 3576
rect 21376 3369 21404 3567
rect 21362 3360 21418 3369
rect 20956 3292 21252 3312
rect 21362 3295 21418 3304
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20810 2000 20866 2009
rect 20810 1935 20866 1944
rect 21836 1737 21864 5238
rect 27066 5199 27122 5208
rect 27080 4865 27108 5199
rect 27066 4856 27122 4865
rect 27066 4791 27122 4800
rect 26054 4720 26110 4729
rect 26054 4655 26110 4664
rect 26068 2990 26096 4655
rect 27434 3768 27490 3777
rect 27434 3703 27436 3712
rect 27488 3703 27490 3712
rect 27436 3674 27488 3680
rect 26698 3632 26754 3641
rect 26698 3567 26754 3576
rect 26882 3632 26938 3641
rect 26882 3567 26938 3576
rect 26712 3233 26740 3567
rect 26698 3224 26754 3233
rect 26698 3159 26754 3168
rect 26056 2984 26108 2990
rect 26896 2961 26924 3567
rect 27540 3194 27568 5471
rect 28276 5030 28304 5646
rect 28552 5522 28580 5714
rect 28630 5536 28686 5545
rect 28552 5494 28630 5522
rect 28630 5471 28686 5480
rect 28644 5370 28672 5471
rect 32140 5409 32168 5714
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 32126 5400 32182 5409
rect 28632 5364 28684 5370
rect 34289 5392 34585 5412
rect 32126 5335 32128 5344
rect 28632 5306 28684 5312
rect 32180 5335 32182 5344
rect 32128 5306 32180 5312
rect 28264 5024 28316 5030
rect 28264 4966 28316 4972
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28276 4729 28304 4966
rect 28262 4720 28318 4729
rect 28262 4655 28318 4664
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 28078 3904 28134 3913
rect 27622 3836 27918 3856
rect 28078 3839 28134 3848
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28092 3369 28120 3839
rect 28170 3768 28226 3777
rect 28170 3703 28226 3712
rect 28356 3732 28408 3738
rect 28078 3360 28134 3369
rect 28078 3295 28134 3304
rect 28078 3224 28134 3233
rect 27528 3188 27580 3194
rect 28078 3159 28134 3168
rect 27528 3130 27580 3136
rect 26056 2926 26108 2932
rect 26882 2952 26938 2961
rect 25872 2848 25924 2854
rect 25870 2816 25872 2825
rect 25924 2816 25926 2825
rect 25870 2751 25926 2760
rect 26068 2650 26096 2926
rect 26882 2887 26938 2896
rect 28092 2825 28120 3159
rect 28184 3097 28212 3703
rect 28356 3674 28408 3680
rect 28368 3097 28396 3674
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 28170 3088 28226 3097
rect 28170 3023 28226 3032
rect 28354 3088 28410 3097
rect 28354 3023 28410 3032
rect 28078 2816 28134 2825
rect 27622 2748 27918 2768
rect 28078 2751 28134 2760
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 26056 2644 26108 2650
rect 26056 2586 26108 2592
rect 34624 2417 34652 8871
rect 34808 8129 34836 12271
rect 34978 12064 35034 12073
rect 34978 11999 35034 12008
rect 34794 8120 34850 8129
rect 34794 8055 34850 8064
rect 34992 7993 35020 11999
rect 35438 11656 35494 11665
rect 35438 11591 35494 11600
rect 35346 10160 35402 10169
rect 35346 10095 35402 10104
rect 34978 7984 35034 7993
rect 34978 7919 35034 7928
rect 35360 3913 35388 10095
rect 35452 10033 35480 11591
rect 35714 11248 35770 11257
rect 35714 11183 35770 11192
rect 35530 10840 35586 10849
rect 35530 10775 35586 10784
rect 35438 10024 35494 10033
rect 35438 9959 35494 9968
rect 35438 9752 35494 9761
rect 35438 9687 35494 9696
rect 35346 3904 35402 3913
rect 35346 3839 35402 3848
rect 35452 3097 35480 9687
rect 35544 6769 35572 10775
rect 35622 10432 35678 10441
rect 35622 10367 35678 10376
rect 35530 6760 35586 6769
rect 35530 6695 35586 6704
rect 35636 6089 35664 10367
rect 35622 6080 35678 6089
rect 35622 6015 35678 6024
rect 35728 5817 35756 11183
rect 35806 8256 35862 8265
rect 35806 8191 35862 8200
rect 35714 5808 35770 5817
rect 35714 5743 35770 5752
rect 35820 3777 35848 8191
rect 39394 7168 39450 7177
rect 39394 7103 39450 7112
rect 39408 7041 39436 7103
rect 39394 7032 39450 7041
rect 39394 6967 39450 6976
rect 35898 6624 35954 6633
rect 35898 6559 35954 6568
rect 35912 5681 35940 6559
rect 35898 5672 35954 5681
rect 35898 5607 35954 5616
rect 35806 3768 35862 3777
rect 35806 3703 35862 3712
rect 35438 3088 35494 3097
rect 35438 3023 35494 3032
rect 34610 2408 34666 2417
rect 34610 2343 34666 2352
rect 35714 2408 35770 2417
rect 35714 2343 35770 2352
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 21822 1728 21878 1737
rect 21822 1663 21878 1672
rect 35728 1465 35756 2343
rect 35714 1456 35770 1465
rect 35714 1391 35770 1400
rect 30470 1320 30526 1329
rect 30470 1255 30526 1264
rect 17866 439 17922 448
rect 15474 368 15530 377
rect 15474 303 15530 312
rect 3422 232 3478 241
rect 3422 167 3478 176
rect 4710 232 4766 241
rect 4710 167 4766 176
rect 3330 96 3386 105
rect 3330 31 3386 40
rect 19982 0 20038 480
rect 30484 105 30512 1255
rect 30838 504 30894 513
rect 30838 439 30894 448
rect 31114 504 31170 513
rect 31114 439 31170 448
rect 30852 241 30880 439
rect 30838 232 30894 241
rect 30838 167 30894 176
rect 31128 105 31156 439
rect 30470 96 30526 105
rect 30470 31 30526 40
rect 31114 96 31170 105
rect 31114 31 31170 40
<< via2 >>
rect 2686 15816 2742 15872
rect 2318 15408 2374 15464
rect 2226 15000 2282 15056
rect 1490 12960 1546 13016
rect 1674 9696 1730 9752
rect 1582 7812 1638 7848
rect 1582 7792 1584 7812
rect 1584 7792 1636 7812
rect 1636 7792 1638 7812
rect 1766 8880 1822 8936
rect 1306 6976 1362 7032
rect 2042 11736 2098 11792
rect 1858 7928 1914 7984
rect 1398 6160 1454 6216
rect 570 5752 626 5808
rect 2410 12552 2466 12608
rect 2226 11192 2282 11248
rect 34886 15816 34942 15872
rect 3422 14592 3478 14648
rect 3330 14184 3386 14240
rect 3054 13368 3110 13424
rect 2134 6296 2190 6352
rect 1858 4936 1914 4992
rect 2042 4664 2098 4720
rect 2870 10920 2926 10976
rect 2778 10512 2834 10568
rect 2502 7112 2558 7168
rect 2502 6704 2558 6760
rect 2410 6024 2466 6080
rect 2318 4392 2374 4448
rect 2042 4004 2098 4040
rect 2042 3984 2044 4004
rect 2044 3984 2096 4004
rect 2096 3984 2098 4004
rect 1674 3476 1676 3496
rect 1676 3476 1728 3496
rect 1728 3476 1730 3496
rect 1674 3440 1730 3476
rect 4066 13812 4068 13832
rect 4068 13812 4120 13832
rect 4120 13812 4122 13832
rect 4066 13776 4122 13812
rect 4066 12144 4122 12200
rect 3238 9288 3294 9344
rect 3146 7384 3202 7440
rect 3698 10104 3754 10160
rect 3606 8472 3662 8528
rect 3422 7384 3478 7440
rect 2686 3068 2688 3088
rect 2688 3068 2740 3088
rect 2740 3068 2742 3088
rect 2686 3032 2742 3068
rect 1582 2372 1638 2408
rect 1582 2352 1584 2372
rect 1584 2352 1636 2372
rect 1636 2352 1638 2372
rect 2042 1400 2098 1456
rect 1398 1264 1454 1320
rect 3238 5072 3294 5128
rect 3422 3848 3478 3904
rect 3238 856 3294 912
rect 2778 448 2834 504
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 4066 9560 4122 9616
rect 7470 9596 7472 9616
rect 7472 9596 7524 9616
rect 7524 9596 7526 9616
rect 7470 9560 7526 9596
rect 7930 9580 7986 9616
rect 7930 9560 7932 9580
rect 7932 9560 7984 9580
rect 7984 9560 7986 9580
rect 4066 8336 4122 8392
rect 3974 6840 4030 6896
rect 3790 6432 3846 6488
rect 4250 8200 4306 8256
rect 4066 6568 4122 6624
rect 6458 6160 6514 6216
rect 5354 5752 5410 5808
rect 3974 5344 4030 5400
rect 3882 5208 3938 5264
rect 3974 4936 4030 4992
rect 3882 4528 3938 4584
rect 3882 4256 3938 4312
rect 3790 4120 3846 4176
rect 4250 4800 4306 4856
rect 4066 3712 4122 3768
rect 3974 3304 4030 3360
rect 6274 4972 6276 4992
rect 6276 4972 6328 4992
rect 6328 4972 6330 4992
rect 6274 4936 6330 4972
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7470 6432 7526 6488
rect 7378 6296 7434 6352
rect 7562 6296 7618 6352
rect 7378 5616 7434 5672
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 34794 15408 34850 15464
rect 34702 15000 34758 15056
rect 34610 14592 34666 14648
rect 34518 14204 34574 14240
rect 34518 14184 34520 14204
rect 34520 14184 34572 14204
rect 34572 14184 34574 14204
rect 17222 12316 17224 12336
rect 17224 12316 17276 12336
rect 17276 12316 17278 12336
rect 17222 12280 17278 12316
rect 19982 12280 20038 12336
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 9862 7928 9918 7984
rect 8482 6840 8538 6896
rect 14094 7148 14096 7168
rect 14096 7148 14148 7168
rect 14148 7148 14150 7168
rect 8390 6604 8392 6624
rect 8392 6604 8444 6624
rect 8444 6604 8446 6624
rect 8390 6568 8446 6604
rect 8298 5344 8354 5400
rect 14094 7112 14150 7148
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14094 6840 14150 6896
rect 18050 11212 18106 11248
rect 18050 11192 18052 11212
rect 18052 11192 18104 11212
rect 18104 11192 18106 11212
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 18510 9560 18566 9616
rect 17774 8372 17776 8392
rect 17776 8372 17828 8392
rect 17828 8372 17830 8392
rect 17774 8336 17830 8372
rect 14738 7148 14740 7168
rect 14740 7148 14792 7168
rect 14792 7148 14794 7168
rect 14738 7112 14794 7148
rect 14646 6704 14702 6760
rect 15474 6432 15530 6488
rect 14094 6024 14150 6080
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 9678 5208 9734 5264
rect 14094 5208 14150 5264
rect 15382 5072 15438 5128
rect 16026 6432 16082 6488
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 8022 4800 8078 4856
rect 8206 4820 8262 4856
rect 8206 4800 8208 4820
rect 8208 4800 8260 4820
rect 8260 4800 8262 4820
rect 7470 4664 7526 4720
rect 7378 4256 7434 4312
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 14094 4800 14150 4856
rect 18418 8880 18474 8936
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 18786 9444 18842 9480
rect 18786 9424 18788 9444
rect 18788 9424 18840 9444
rect 18840 9424 18842 9444
rect 18694 9152 18750 9208
rect 20994 9152 21050 9208
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 27894 11192 27950 11248
rect 26606 10104 26662 10160
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 34518 13912 34574 13968
rect 34610 13504 34666 13560
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34518 12708 34574 12744
rect 34518 12688 34520 12708
rect 34520 12688 34572 12708
rect 34572 12688 34574 12708
rect 34702 13096 34758 13152
rect 34794 12280 34850 12336
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 28906 10104 28962 10160
rect 26974 9424 27030 9480
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 17590 6432 17646 6488
rect 17314 6160 17370 6216
rect 17590 6160 17646 6216
rect 8022 4256 8078 4312
rect 7470 4120 7526 4176
rect 14094 3848 14150 3904
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 9862 3576 9918 3632
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 8574 3340 8576 3360
rect 8576 3340 8628 3360
rect 8628 3340 8630 3360
rect 8574 3304 8630 3340
rect 3882 2896 3938 2952
rect 4342 2896 4398 2952
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 9678 2624 9734 2680
rect 7470 2488 7526 2544
rect 8390 2488 8446 2544
rect 3698 1808 3754 1864
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 7470 2080 7526 2136
rect 17314 5752 17370 5808
rect 17314 5208 17370 5264
rect 16670 4936 16726 4992
rect 16578 4276 16634 4312
rect 16578 4256 16580 4276
rect 16580 4256 16632 4276
rect 16632 4256 16634 4276
rect 17222 3712 17278 3768
rect 17222 3304 17278 3360
rect 21546 9036 21602 9072
rect 21546 9016 21548 9036
rect 21548 9016 21600 9036
rect 21600 9016 21602 9036
rect 30654 9424 30710 9480
rect 29366 9016 29422 9072
rect 32402 9968 32458 10024
rect 32310 9288 32366 9344
rect 32126 8880 32182 8936
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 28078 8064 28134 8120
rect 28078 7792 28134 7848
rect 21454 7520 21510 7576
rect 20810 6840 20866 6896
rect 21270 6840 21326 6896
rect 18878 6568 18934 6624
rect 20534 6724 20590 6760
rect 20534 6704 20536 6724
rect 20536 6704 20588 6724
rect 20588 6704 20590 6724
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 27434 7148 27436 7168
rect 27436 7148 27488 7168
rect 27488 7148 27490 7168
rect 27434 7112 27490 7148
rect 28078 7148 28080 7168
rect 28080 7148 28132 7168
rect 28132 7148 28134 7168
rect 28078 7112 28134 7148
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 21546 6724 21602 6760
rect 21546 6704 21548 6724
rect 21548 6704 21600 6724
rect 21600 6704 21602 6724
rect 28170 6704 28226 6760
rect 26790 6432 26846 6488
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20718 4428 20720 4448
rect 20720 4428 20772 4448
rect 20772 4428 20774 4448
rect 20718 4392 20774 4428
rect 18602 3848 18658 3904
rect 19982 2760 20038 2816
rect 18970 2508 19026 2544
rect 18970 2488 18972 2508
rect 18972 2488 19024 2508
rect 19024 2488 19026 2508
rect 18510 1808 18566 1864
rect 17866 448 17922 504
rect 28078 6296 28134 6352
rect 28078 6024 28134 6080
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 28170 5888 28226 5944
rect 32126 7520 32182 7576
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34610 8880 34666 8936
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 32494 8200 32550 8256
rect 32402 7792 32458 7848
rect 32034 6568 32090 6624
rect 32126 6196 32128 6216
rect 32128 6196 32180 6216
rect 32180 6196 32182 6216
rect 32126 6160 32182 6196
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 26790 5752 26846 5808
rect 27526 5480 27582 5536
rect 21730 5364 21786 5400
rect 21730 5344 21732 5364
rect 21732 5344 21784 5364
rect 21784 5344 21786 5364
rect 21546 5208 21602 5264
rect 21546 4936 21602 4992
rect 21362 4428 21364 4448
rect 21364 4428 21416 4448
rect 21416 4428 21418 4448
rect 21362 4392 21418 4428
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 21546 3984 21602 4040
rect 21362 3576 21418 3632
rect 21546 3576 21602 3632
rect 21362 3304 21418 3360
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20810 1944 20866 2000
rect 27066 5208 27122 5264
rect 27066 4800 27122 4856
rect 26054 4664 26110 4720
rect 27434 3732 27490 3768
rect 27434 3712 27436 3732
rect 27436 3712 27488 3732
rect 27488 3712 27490 3732
rect 26698 3576 26754 3632
rect 26882 3576 26938 3632
rect 26698 3168 26754 3224
rect 28630 5480 28686 5536
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 32126 5364 32182 5400
rect 32126 5344 32128 5364
rect 32128 5344 32180 5364
rect 32180 5344 32182 5364
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 28262 4664 28318 4720
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 28078 3848 28134 3904
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 28170 3712 28226 3768
rect 28078 3304 28134 3360
rect 28078 3168 28134 3224
rect 25870 2796 25872 2816
rect 25872 2796 25924 2816
rect 25924 2796 25926 2816
rect 25870 2760 25926 2796
rect 26882 2896 26938 2952
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 28170 3032 28226 3088
rect 28354 3032 28410 3088
rect 28078 2760 28134 2816
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 34978 12008 35034 12064
rect 34794 8064 34850 8120
rect 35438 11600 35494 11656
rect 35346 10104 35402 10160
rect 34978 7928 35034 7984
rect 35714 11192 35770 11248
rect 35530 10784 35586 10840
rect 35438 9968 35494 10024
rect 35438 9696 35494 9752
rect 35346 3848 35402 3904
rect 35622 10376 35678 10432
rect 35530 6704 35586 6760
rect 35622 6024 35678 6080
rect 35806 8200 35862 8256
rect 35714 5752 35770 5808
rect 39394 7112 39450 7168
rect 39394 6976 39450 7032
rect 35898 6568 35954 6624
rect 35898 5616 35954 5672
rect 35806 3712 35862 3768
rect 35438 3032 35494 3088
rect 34610 2352 34666 2408
rect 35714 2352 35770 2408
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 21822 1672 21878 1728
rect 35714 1400 35770 1456
rect 30470 1264 30526 1320
rect 15474 312 15530 368
rect 3422 176 3478 232
rect 4710 176 4766 232
rect 3330 40 3386 96
rect 30838 448 30894 504
rect 31114 448 31170 504
rect 30838 176 30894 232
rect 30470 40 30526 96
rect 31114 40 31170 96
<< metal3 >>
rect 0 15874 480 15904
rect 2681 15874 2747 15877
rect 0 15872 2747 15874
rect 0 15816 2686 15872
rect 2742 15816 2747 15872
rect 0 15814 2747 15816
rect 0 15784 480 15814
rect 2681 15811 2747 15814
rect 34881 15874 34947 15877
rect 39520 15874 40000 15904
rect 34881 15872 40000 15874
rect 34881 15816 34886 15872
rect 34942 15816 40000 15872
rect 34881 15814 40000 15816
rect 34881 15811 34947 15814
rect 39520 15784 40000 15814
rect 0 15466 480 15496
rect 2313 15466 2379 15469
rect 0 15464 2379 15466
rect 0 15408 2318 15464
rect 2374 15408 2379 15464
rect 0 15406 2379 15408
rect 0 15376 480 15406
rect 2313 15403 2379 15406
rect 34789 15466 34855 15469
rect 39520 15466 40000 15496
rect 34789 15464 40000 15466
rect 34789 15408 34794 15464
rect 34850 15408 40000 15464
rect 34789 15406 40000 15408
rect 34789 15403 34855 15406
rect 39520 15376 40000 15406
rect 0 15058 480 15088
rect 2221 15058 2287 15061
rect 0 15056 2287 15058
rect 0 15000 2226 15056
rect 2282 15000 2287 15056
rect 0 14998 2287 15000
rect 0 14968 480 14998
rect 2221 14995 2287 14998
rect 34697 15058 34763 15061
rect 39520 15058 40000 15088
rect 34697 15056 40000 15058
rect 34697 15000 34702 15056
rect 34758 15000 40000 15056
rect 34697 14998 40000 15000
rect 34697 14995 34763 14998
rect 39520 14968 40000 14998
rect 0 14650 480 14680
rect 3417 14650 3483 14653
rect 0 14648 3483 14650
rect 0 14592 3422 14648
rect 3478 14592 3483 14648
rect 0 14590 3483 14592
rect 0 14560 480 14590
rect 3417 14587 3483 14590
rect 34605 14650 34671 14653
rect 39520 14650 40000 14680
rect 34605 14648 40000 14650
rect 34605 14592 34610 14648
rect 34666 14592 40000 14648
rect 34605 14590 40000 14592
rect 34605 14587 34671 14590
rect 39520 14560 40000 14590
rect 0 14242 480 14272
rect 3325 14242 3391 14245
rect 0 14240 3391 14242
rect 0 14184 3330 14240
rect 3386 14184 3391 14240
rect 0 14182 3391 14184
rect 0 14152 480 14182
rect 3325 14179 3391 14182
rect 34513 14242 34579 14245
rect 39520 14242 40000 14272
rect 34513 14240 40000 14242
rect 34513 14184 34518 14240
rect 34574 14184 40000 14240
rect 34513 14182 40000 14184
rect 34513 14179 34579 14182
rect 39520 14152 40000 14182
rect 34513 13970 34579 13973
rect 39520 13970 40000 14000
rect 34513 13968 40000 13970
rect 34513 13912 34518 13968
rect 34574 13912 40000 13968
rect 34513 13910 40000 13912
rect 34513 13907 34579 13910
rect 39520 13880 40000 13910
rect 0 13834 480 13864
rect 4061 13834 4127 13837
rect 0 13832 4127 13834
rect 0 13776 4066 13832
rect 4122 13776 4127 13832
rect 0 13774 4127 13776
rect 0 13744 480 13774
rect 4061 13771 4127 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 34605 13562 34671 13565
rect 39520 13562 40000 13592
rect 34605 13560 40000 13562
rect 34605 13504 34610 13560
rect 34666 13504 40000 13560
rect 34605 13502 40000 13504
rect 34605 13499 34671 13502
rect 39520 13472 40000 13502
rect 0 13426 480 13456
rect 3049 13426 3115 13429
rect 0 13424 3115 13426
rect 0 13368 3054 13424
rect 3110 13368 3115 13424
rect 0 13366 3115 13368
rect 0 13336 480 13366
rect 3049 13363 3115 13366
rect 34697 13154 34763 13157
rect 39520 13154 40000 13184
rect 34697 13152 40000 13154
rect 34697 13096 34702 13152
rect 34758 13096 40000 13152
rect 34697 13094 40000 13096
rect 34697 13091 34763 13094
rect 7610 13088 7930 13089
rect 0 13018 480 13048
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 39520 13064 40000 13094
rect 34277 13023 34597 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 480 12958
rect 1485 12955 1551 12958
rect 34513 12746 34579 12749
rect 39520 12746 40000 12776
rect 34513 12744 40000 12746
rect 34513 12688 34518 12744
rect 34574 12688 40000 12744
rect 34513 12686 40000 12688
rect 34513 12683 34579 12686
rect 39520 12656 40000 12686
rect 0 12610 480 12640
rect 2405 12610 2471 12613
rect 0 12608 2471 12610
rect 0 12552 2410 12608
rect 2466 12552 2471 12608
rect 0 12550 2471 12552
rect 0 12520 480 12550
rect 2405 12547 2471 12550
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 17217 12338 17283 12341
rect 19977 12338 20043 12341
rect 17217 12336 20043 12338
rect 17217 12280 17222 12336
rect 17278 12280 19982 12336
rect 20038 12280 20043 12336
rect 17217 12278 20043 12280
rect 17217 12275 17283 12278
rect 19977 12275 20043 12278
rect 34789 12338 34855 12341
rect 39520 12338 40000 12368
rect 34789 12336 40000 12338
rect 34789 12280 34794 12336
rect 34850 12280 40000 12336
rect 34789 12278 40000 12280
rect 34789 12275 34855 12278
rect 39520 12248 40000 12278
rect 0 12202 480 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 480 12142
rect 4061 12139 4127 12142
rect 34973 12066 35039 12069
rect 39520 12066 40000 12096
rect 34973 12064 40000 12066
rect 34973 12008 34978 12064
rect 35034 12008 40000 12064
rect 34973 12006 40000 12008
rect 34973 12003 35039 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12006
rect 34277 11935 34597 11936
rect 0 11794 480 11824
rect 2037 11794 2103 11797
rect 0 11792 2103 11794
rect 0 11736 2042 11792
rect 2098 11736 2103 11792
rect 0 11734 2103 11736
rect 0 11704 480 11734
rect 2037 11731 2103 11734
rect 35433 11658 35499 11661
rect 39520 11658 40000 11688
rect 35433 11656 40000 11658
rect 35433 11600 35438 11656
rect 35494 11600 40000 11656
rect 35433 11598 40000 11600
rect 35433 11595 35499 11598
rect 39520 11568 40000 11598
rect 14277 11456 14597 11457
rect 0 11386 480 11416
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 0 11326 2146 11386
rect 0 11296 480 11326
rect 2086 11250 2146 11326
rect 2221 11250 2287 11253
rect 2086 11248 2287 11250
rect 2086 11192 2226 11248
rect 2282 11192 2287 11248
rect 2086 11190 2287 11192
rect 2221 11187 2287 11190
rect 18045 11250 18111 11253
rect 27889 11250 27955 11253
rect 18045 11248 27955 11250
rect 18045 11192 18050 11248
rect 18106 11192 27894 11248
rect 27950 11192 27955 11248
rect 18045 11190 27955 11192
rect 18045 11187 18111 11190
rect 27889 11187 27955 11190
rect 35709 11250 35775 11253
rect 39520 11250 40000 11280
rect 35709 11248 40000 11250
rect 35709 11192 35714 11248
rect 35770 11192 40000 11248
rect 35709 11190 40000 11192
rect 35709 11187 35775 11190
rect 39520 11160 40000 11190
rect 0 10978 480 11008
rect 2865 10978 2931 10981
rect 0 10976 2931 10978
rect 0 10920 2870 10976
rect 2926 10920 2931 10976
rect 0 10918 2931 10920
rect 0 10888 480 10918
rect 2865 10915 2931 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 35525 10842 35591 10845
rect 39520 10842 40000 10872
rect 35525 10840 40000 10842
rect 35525 10784 35530 10840
rect 35586 10784 40000 10840
rect 35525 10782 40000 10784
rect 35525 10779 35591 10782
rect 39520 10752 40000 10782
rect 0 10570 480 10600
rect 2773 10570 2839 10573
rect 0 10568 2839 10570
rect 0 10512 2778 10568
rect 2834 10512 2839 10568
rect 0 10510 2839 10512
rect 0 10480 480 10510
rect 2773 10507 2839 10510
rect 35617 10434 35683 10437
rect 39520 10434 40000 10464
rect 35617 10432 40000 10434
rect 35617 10376 35622 10432
rect 35678 10376 40000 10432
rect 35617 10374 40000 10376
rect 35617 10371 35683 10374
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 39520 10344 40000 10374
rect 27610 10303 27930 10304
rect 0 10162 480 10192
rect 3693 10162 3759 10165
rect 0 10160 3759 10162
rect 0 10104 3698 10160
rect 3754 10104 3759 10160
rect 0 10102 3759 10104
rect 0 10072 480 10102
rect 3693 10099 3759 10102
rect 26601 10162 26667 10165
rect 28901 10162 28967 10165
rect 26601 10160 28967 10162
rect 26601 10104 26606 10160
rect 26662 10104 28906 10160
rect 28962 10104 28967 10160
rect 26601 10102 28967 10104
rect 26601 10099 26667 10102
rect 28901 10099 28967 10102
rect 35341 10162 35407 10165
rect 39520 10162 40000 10192
rect 35341 10160 40000 10162
rect 35341 10104 35346 10160
rect 35402 10104 40000 10160
rect 35341 10102 40000 10104
rect 35341 10099 35407 10102
rect 39520 10072 40000 10102
rect 32397 10026 32463 10029
rect 35433 10026 35499 10029
rect 32397 10024 35499 10026
rect 32397 9968 32402 10024
rect 32458 9968 35438 10024
rect 35494 9968 35499 10024
rect 32397 9966 35499 9968
rect 32397 9963 32463 9966
rect 35433 9963 35499 9966
rect 7610 9824 7930 9825
rect 0 9754 480 9784
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 1669 9754 1735 9757
rect 0 9752 1735 9754
rect 0 9696 1674 9752
rect 1730 9696 1735 9752
rect 0 9694 1735 9696
rect 0 9664 480 9694
rect 1669 9691 1735 9694
rect 35433 9754 35499 9757
rect 39520 9754 40000 9784
rect 35433 9752 40000 9754
rect 35433 9696 35438 9752
rect 35494 9696 40000 9752
rect 35433 9694 40000 9696
rect 35433 9691 35499 9694
rect 39520 9664 40000 9694
rect 4061 9618 4127 9621
rect 7465 9618 7531 9621
rect 4061 9616 7531 9618
rect 4061 9560 4066 9616
rect 4122 9560 7470 9616
rect 7526 9560 7531 9616
rect 4061 9558 7531 9560
rect 4061 9555 4127 9558
rect 7465 9555 7531 9558
rect 7925 9618 7991 9621
rect 18505 9618 18571 9621
rect 7925 9616 18571 9618
rect 7925 9560 7930 9616
rect 7986 9560 18510 9616
rect 18566 9560 18571 9616
rect 7925 9558 18571 9560
rect 7925 9555 7991 9558
rect 18505 9555 18571 9558
rect 18781 9482 18847 9485
rect 26969 9482 27035 9485
rect 30649 9482 30715 9485
rect 18781 9480 30715 9482
rect 18781 9424 18786 9480
rect 18842 9424 26974 9480
rect 27030 9424 30654 9480
rect 30710 9424 30715 9480
rect 18781 9422 30715 9424
rect 18781 9419 18847 9422
rect 26969 9419 27035 9422
rect 30649 9419 30715 9422
rect 0 9346 480 9376
rect 3233 9346 3299 9349
rect 0 9344 3299 9346
rect 0 9288 3238 9344
rect 3294 9288 3299 9344
rect 0 9286 3299 9288
rect 0 9256 480 9286
rect 3233 9283 3299 9286
rect 32305 9346 32371 9349
rect 39520 9346 40000 9376
rect 32305 9344 40000 9346
rect 32305 9288 32310 9344
rect 32366 9288 40000 9344
rect 32305 9286 40000 9288
rect 32305 9283 32371 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 18689 9210 18755 9213
rect 20989 9210 21055 9213
rect 18689 9208 21055 9210
rect 18689 9152 18694 9208
rect 18750 9152 20994 9208
rect 21050 9152 21055 9208
rect 18689 9150 21055 9152
rect 18689 9147 18755 9150
rect 20989 9147 21055 9150
rect 21541 9074 21607 9077
rect 29361 9074 29427 9077
rect 21541 9072 29427 9074
rect 21541 9016 21546 9072
rect 21602 9016 29366 9072
rect 29422 9016 29427 9072
rect 21541 9014 29427 9016
rect 21541 9011 21607 9014
rect 29361 9011 29427 9014
rect 0 8938 480 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 480 8878
rect 1761 8875 1827 8878
rect 18413 8938 18479 8941
rect 32121 8938 32187 8941
rect 18413 8936 32187 8938
rect 18413 8880 18418 8936
rect 18474 8880 32126 8936
rect 32182 8880 32187 8936
rect 18413 8878 32187 8880
rect 18413 8875 18479 8878
rect 32121 8875 32187 8878
rect 34605 8938 34671 8941
rect 39520 8938 40000 8968
rect 34605 8936 40000 8938
rect 34605 8880 34610 8936
rect 34666 8880 40000 8936
rect 34605 8878 40000 8880
rect 34605 8875 34671 8878
rect 39520 8848 40000 8878
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8530 480 8560
rect 3601 8530 3667 8533
rect 39520 8530 40000 8560
rect 0 8528 3667 8530
rect 0 8472 3606 8528
rect 3662 8472 3667 8528
rect 0 8470 3667 8472
rect 0 8440 480 8470
rect 3601 8467 3667 8470
rect 35390 8470 40000 8530
rect 4061 8394 4127 8397
rect 17769 8394 17835 8397
rect 4061 8392 17835 8394
rect 4061 8336 4066 8392
rect 4122 8336 17774 8392
rect 17830 8336 17835 8392
rect 4061 8334 17835 8336
rect 4061 8331 4127 8334
rect 17769 8331 17835 8334
rect 0 8258 480 8288
rect 4245 8258 4311 8261
rect 0 8256 4311 8258
rect 0 8200 4250 8256
rect 4306 8200 4311 8256
rect 0 8198 4311 8200
rect 0 8168 480 8198
rect 4245 8195 4311 8198
rect 32489 8258 32555 8261
rect 35390 8258 35450 8470
rect 39520 8440 40000 8470
rect 32489 8256 35450 8258
rect 32489 8200 32494 8256
rect 32550 8200 35450 8256
rect 32489 8198 35450 8200
rect 35801 8258 35867 8261
rect 39520 8258 40000 8288
rect 35801 8256 40000 8258
rect 35801 8200 35806 8256
rect 35862 8200 40000 8256
rect 35801 8198 40000 8200
rect 32489 8195 32555 8198
rect 35801 8195 35867 8198
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 39520 8168 40000 8198
rect 27610 8127 27930 8128
rect 28073 8122 28139 8125
rect 34789 8122 34855 8125
rect 28073 8120 34855 8122
rect 28073 8064 28078 8120
rect 28134 8064 34794 8120
rect 34850 8064 34855 8120
rect 28073 8062 34855 8064
rect 28073 8059 28139 8062
rect 34789 8059 34855 8062
rect 1853 7986 1919 7989
rect 1350 7984 1919 7986
rect 1350 7928 1858 7984
rect 1914 7928 1919 7984
rect 1350 7926 1919 7928
rect 0 7850 480 7880
rect 1350 7850 1410 7926
rect 1853 7923 1919 7926
rect 9857 7986 9923 7989
rect 34973 7986 35039 7989
rect 9857 7984 35039 7986
rect 9857 7928 9862 7984
rect 9918 7928 34978 7984
rect 35034 7928 35039 7984
rect 9857 7926 35039 7928
rect 9857 7923 9923 7926
rect 34973 7923 35039 7926
rect 0 7790 1410 7850
rect 1577 7850 1643 7853
rect 28073 7850 28139 7853
rect 1577 7848 28139 7850
rect 1577 7792 1582 7848
rect 1638 7792 28078 7848
rect 28134 7792 28139 7848
rect 1577 7790 28139 7792
rect 0 7760 480 7790
rect 1577 7787 1643 7790
rect 28073 7787 28139 7790
rect 32397 7850 32463 7853
rect 39520 7850 40000 7880
rect 32397 7848 40000 7850
rect 32397 7792 32402 7848
rect 32458 7792 40000 7848
rect 32397 7790 40000 7792
rect 32397 7787 32463 7790
rect 39520 7760 40000 7790
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 21449 7578 21515 7581
rect 32121 7578 32187 7581
rect 21449 7576 32187 7578
rect 21449 7520 21454 7576
rect 21510 7520 32126 7576
rect 32182 7520 32187 7576
rect 21449 7518 32187 7520
rect 21449 7515 21515 7518
rect 32121 7515 32187 7518
rect 0 7442 480 7472
rect 3141 7442 3207 7445
rect 0 7440 3207 7442
rect 0 7384 3146 7440
rect 3202 7384 3207 7440
rect 0 7382 3207 7384
rect 0 7352 480 7382
rect 3141 7379 3207 7382
rect 3417 7442 3483 7445
rect 39520 7442 40000 7472
rect 3417 7440 40000 7442
rect 3417 7384 3422 7440
rect 3478 7384 40000 7440
rect 3417 7382 40000 7384
rect 3417 7379 3483 7382
rect 39520 7352 40000 7382
rect 2497 7170 2563 7173
rect 14089 7170 14155 7173
rect 2497 7168 14155 7170
rect 2497 7112 2502 7168
rect 2558 7112 14094 7168
rect 14150 7112 14155 7168
rect 2497 7110 14155 7112
rect 2497 7107 2563 7110
rect 14089 7107 14155 7110
rect 14733 7170 14799 7173
rect 27429 7170 27495 7173
rect 14733 7168 27495 7170
rect 14733 7112 14738 7168
rect 14794 7112 27434 7168
rect 27490 7112 27495 7168
rect 14733 7110 27495 7112
rect 14733 7107 14799 7110
rect 27429 7107 27495 7110
rect 28073 7170 28139 7173
rect 39389 7170 39455 7173
rect 28073 7168 39455 7170
rect 28073 7112 28078 7168
rect 28134 7112 39394 7168
rect 39450 7112 39455 7168
rect 28073 7110 39455 7112
rect 28073 7107 28139 7110
rect 39389 7107 39455 7110
rect 14277 7104 14597 7105
rect 0 7034 480 7064
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 1301 7034 1367 7037
rect 0 7032 1367 7034
rect 0 6976 1306 7032
rect 1362 6976 1367 7032
rect 0 6974 1367 6976
rect 0 6944 480 6974
rect 1301 6971 1367 6974
rect 39389 7034 39455 7037
rect 39520 7034 40000 7064
rect 39389 7032 40000 7034
rect 39389 6976 39394 7032
rect 39450 6976 40000 7032
rect 39389 6974 40000 6976
rect 39389 6971 39455 6974
rect 39520 6944 40000 6974
rect 3969 6898 4035 6901
rect 8477 6898 8543 6901
rect 3969 6896 8543 6898
rect 3969 6840 3974 6896
rect 4030 6840 8482 6896
rect 8538 6840 8543 6896
rect 3969 6838 8543 6840
rect 3969 6835 4035 6838
rect 8477 6835 8543 6838
rect 14089 6898 14155 6901
rect 20805 6898 20871 6901
rect 14089 6896 20871 6898
rect 14089 6840 14094 6896
rect 14150 6840 20810 6896
rect 20866 6840 20871 6896
rect 14089 6838 20871 6840
rect 14089 6835 14155 6838
rect 20805 6835 20871 6838
rect 21265 6898 21331 6901
rect 21265 6896 35772 6898
rect 21265 6840 21270 6896
rect 21326 6840 35772 6896
rect 21265 6838 35772 6840
rect 21265 6835 21331 6838
rect 2497 6762 2563 6765
rect 14641 6762 14707 6765
rect 20529 6762 20595 6765
rect 21541 6762 21607 6765
rect 28165 6762 28231 6765
rect 35525 6762 35591 6765
rect 2497 6760 8218 6762
rect 2497 6704 2502 6760
rect 2558 6704 8218 6760
rect 2497 6702 8218 6704
rect 2497 6699 2563 6702
rect 0 6626 480 6656
rect 4061 6626 4127 6629
rect 0 6624 4127 6626
rect 0 6568 4066 6624
rect 4122 6568 4127 6624
rect 0 6566 4127 6568
rect 0 6536 480 6566
rect 4061 6563 4127 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 3785 6490 3851 6493
rect 7465 6490 7531 6493
rect 3785 6488 7531 6490
rect 3785 6432 3790 6488
rect 3846 6432 7470 6488
rect 7526 6432 7531 6488
rect 3785 6430 7531 6432
rect 8158 6490 8218 6702
rect 14641 6760 20595 6762
rect 14641 6704 14646 6760
rect 14702 6704 20534 6760
rect 20590 6704 20595 6760
rect 14641 6702 20595 6704
rect 14641 6699 14707 6702
rect 20529 6699 20595 6702
rect 20670 6702 21466 6762
rect 8385 6626 8451 6629
rect 18873 6626 18939 6629
rect 20670 6626 20730 6702
rect 8385 6624 20730 6626
rect 8385 6568 8390 6624
rect 8446 6568 18878 6624
rect 18934 6568 20730 6624
rect 8385 6566 20730 6568
rect 21406 6626 21466 6702
rect 21541 6760 28231 6762
rect 21541 6704 21546 6760
rect 21602 6704 28170 6760
rect 28226 6704 28231 6760
rect 21541 6702 28231 6704
rect 21541 6699 21607 6702
rect 28165 6699 28231 6702
rect 34102 6760 35591 6762
rect 34102 6704 35530 6760
rect 35586 6704 35591 6760
rect 34102 6702 35591 6704
rect 32029 6626 32095 6629
rect 21406 6624 32095 6626
rect 21406 6568 32034 6624
rect 32090 6568 32095 6624
rect 21406 6566 32095 6568
rect 8385 6563 8451 6566
rect 18873 6563 18939 6566
rect 32029 6563 32095 6566
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 15469 6490 15535 6493
rect 8158 6488 15535 6490
rect 8158 6432 15474 6488
rect 15530 6432 15535 6488
rect 8158 6430 15535 6432
rect 3785 6427 3851 6430
rect 7465 6427 7531 6430
rect 15469 6427 15535 6430
rect 16021 6490 16087 6493
rect 17585 6490 17651 6493
rect 16021 6488 17651 6490
rect 16021 6432 16026 6488
rect 16082 6432 17590 6488
rect 17646 6432 17651 6488
rect 16021 6430 17651 6432
rect 16021 6427 16087 6430
rect 17585 6427 17651 6430
rect 26785 6490 26851 6493
rect 34102 6490 34162 6702
rect 35525 6699 35591 6702
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 26785 6488 34162 6490
rect 26785 6432 26790 6488
rect 26846 6432 34162 6488
rect 26785 6430 34162 6432
rect 26785 6427 26851 6430
rect 2129 6354 2195 6357
rect 7373 6354 7439 6357
rect 2129 6352 7439 6354
rect 2129 6296 2134 6352
rect 2190 6296 7378 6352
rect 7434 6296 7439 6352
rect 2129 6294 7439 6296
rect 2129 6291 2195 6294
rect 7373 6291 7439 6294
rect 7557 6354 7623 6357
rect 28073 6354 28139 6357
rect 7557 6352 28139 6354
rect 7557 6296 7562 6352
rect 7618 6296 28078 6352
rect 28134 6296 28139 6352
rect 7557 6294 28139 6296
rect 7557 6291 7623 6294
rect 28073 6291 28139 6294
rect 0 6218 480 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 480 6158
rect 1393 6155 1459 6158
rect 6453 6218 6519 6221
rect 17309 6218 17375 6221
rect 6453 6216 17375 6218
rect 6453 6160 6458 6216
rect 6514 6160 17314 6216
rect 17370 6160 17375 6216
rect 6453 6158 17375 6160
rect 6453 6155 6519 6158
rect 17309 6155 17375 6158
rect 17585 6218 17651 6221
rect 32121 6218 32187 6221
rect 17585 6216 32187 6218
rect 17585 6160 17590 6216
rect 17646 6160 32126 6216
rect 32182 6160 32187 6216
rect 17585 6158 32187 6160
rect 35712 6218 35772 6838
rect 35893 6626 35959 6629
rect 39520 6626 40000 6656
rect 35893 6624 40000 6626
rect 35893 6568 35898 6624
rect 35954 6568 40000 6624
rect 35893 6566 40000 6568
rect 35893 6563 35959 6566
rect 39520 6536 40000 6566
rect 39520 6218 40000 6248
rect 35712 6158 40000 6218
rect 17585 6155 17651 6158
rect 32121 6155 32187 6158
rect 39520 6128 40000 6158
rect 2405 6082 2471 6085
rect 14089 6082 14155 6085
rect 2405 6080 14155 6082
rect 2405 6024 2410 6080
rect 2466 6024 14094 6080
rect 14150 6024 14155 6080
rect 2405 6022 14155 6024
rect 2405 6019 2471 6022
rect 14089 6019 14155 6022
rect 28073 6082 28139 6085
rect 35617 6082 35683 6085
rect 28073 6080 35683 6082
rect 28073 6024 28078 6080
rect 28134 6024 35622 6080
rect 35678 6024 35683 6080
rect 28073 6022 35683 6024
rect 28073 6019 28139 6022
rect 35617 6019 35683 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 28165 5946 28231 5949
rect 39520 5946 40000 5976
rect 17174 5886 26986 5946
rect 0 5810 480 5840
rect 565 5810 631 5813
rect 0 5808 631 5810
rect 0 5752 570 5808
rect 626 5752 631 5808
rect 0 5750 631 5752
rect 0 5720 480 5750
rect 565 5747 631 5750
rect 5349 5810 5415 5813
rect 17174 5810 17234 5886
rect 5349 5808 17234 5810
rect 5349 5752 5354 5808
rect 5410 5752 17234 5808
rect 5349 5750 17234 5752
rect 17309 5810 17375 5813
rect 26785 5810 26851 5813
rect 17309 5808 26851 5810
rect 17309 5752 17314 5808
rect 17370 5752 26790 5808
rect 26846 5752 26851 5808
rect 17309 5750 26851 5752
rect 26926 5810 26986 5886
rect 28165 5944 40000 5946
rect 28165 5888 28170 5944
rect 28226 5888 40000 5944
rect 28165 5886 40000 5888
rect 28165 5883 28231 5886
rect 39520 5856 40000 5886
rect 35709 5810 35775 5813
rect 26926 5808 35775 5810
rect 26926 5752 35714 5808
rect 35770 5752 35775 5808
rect 26926 5750 35775 5752
rect 5349 5747 5415 5750
rect 17309 5747 17375 5750
rect 26785 5747 26851 5750
rect 35709 5747 35775 5750
rect 7373 5674 7439 5677
rect 35893 5674 35959 5677
rect 7373 5672 35959 5674
rect 7373 5616 7378 5672
rect 7434 5616 35898 5672
rect 35954 5616 35959 5672
rect 7373 5614 35959 5616
rect 7373 5611 7439 5614
rect 35893 5611 35959 5614
rect 27521 5538 27587 5541
rect 28625 5538 28691 5541
rect 39520 5538 40000 5568
rect 26742 5536 28691 5538
rect 26742 5480 27526 5536
rect 27582 5480 28630 5536
rect 28686 5480 28691 5536
rect 26742 5478 28691 5480
rect 7610 5472 7930 5473
rect 0 5402 480 5432
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 3969 5402 4035 5405
rect 0 5400 4035 5402
rect 0 5344 3974 5400
rect 4030 5344 4035 5400
rect 0 5342 4035 5344
rect 0 5312 480 5342
rect 3969 5339 4035 5342
rect 8293 5402 8359 5405
rect 21725 5402 21791 5405
rect 26742 5402 26802 5478
rect 27521 5475 27587 5478
rect 28625 5475 28691 5478
rect 35712 5478 40000 5538
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 32121 5402 32187 5405
rect 8293 5400 17234 5402
rect 8293 5344 8298 5400
rect 8354 5344 17234 5400
rect 8293 5342 17234 5344
rect 8293 5339 8359 5342
rect 3877 5266 3943 5269
rect 9673 5266 9739 5269
rect 3877 5264 9739 5266
rect 3877 5208 3882 5264
rect 3938 5208 9678 5264
rect 9734 5208 9739 5264
rect 3877 5206 9739 5208
rect 3877 5203 3943 5206
rect 9673 5203 9739 5206
rect 14089 5266 14155 5269
rect 14089 5264 15578 5266
rect 14089 5208 14094 5264
rect 14150 5208 15578 5264
rect 14089 5206 15578 5208
rect 14089 5203 14155 5206
rect 3233 5130 3299 5133
rect 15377 5130 15443 5133
rect 3233 5128 15443 5130
rect 3233 5072 3238 5128
rect 3294 5072 15382 5128
rect 15438 5072 15443 5128
rect 3233 5070 15443 5072
rect 3233 5067 3299 5070
rect 15377 5067 15443 5070
rect 0 4994 480 5024
rect 1853 4994 1919 4997
rect 0 4992 1919 4994
rect 0 4936 1858 4992
rect 1914 4936 1919 4992
rect 0 4934 1919 4936
rect 0 4904 480 4934
rect 1853 4931 1919 4934
rect 3969 4994 4035 4997
rect 6269 4994 6335 4997
rect 3969 4992 6335 4994
rect 3969 4936 3974 4992
rect 4030 4936 6274 4992
rect 6330 4936 6335 4992
rect 3969 4934 6335 4936
rect 3969 4931 4035 4934
rect 6269 4931 6335 4934
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 4245 4858 4311 4861
rect 8017 4858 8083 4861
rect 4245 4856 8083 4858
rect 4245 4800 4250 4856
rect 4306 4800 8022 4856
rect 8078 4800 8083 4856
rect 4245 4798 8083 4800
rect 4245 4795 4311 4798
rect 8017 4795 8083 4798
rect 8201 4858 8267 4861
rect 14089 4858 14155 4861
rect 8201 4856 14155 4858
rect 8201 4800 8206 4856
rect 8262 4800 14094 4856
rect 14150 4800 14155 4856
rect 8201 4798 14155 4800
rect 15518 4858 15578 5206
rect 17174 5130 17234 5342
rect 21406 5400 26802 5402
rect 21406 5344 21730 5400
rect 21786 5344 26802 5400
rect 21406 5342 26802 5344
rect 26926 5400 32187 5402
rect 26926 5344 32126 5400
rect 32182 5344 32187 5400
rect 26926 5342 32187 5344
rect 17309 5266 17375 5269
rect 21406 5266 21466 5342
rect 21725 5339 21791 5342
rect 17309 5264 21466 5266
rect 17309 5208 17314 5264
rect 17370 5208 21466 5264
rect 17309 5206 21466 5208
rect 21541 5266 21607 5269
rect 26926 5266 26986 5342
rect 32121 5339 32187 5342
rect 21541 5264 26986 5266
rect 21541 5208 21546 5264
rect 21602 5208 26986 5264
rect 21541 5206 26986 5208
rect 27061 5266 27127 5269
rect 35712 5266 35772 5478
rect 39520 5448 40000 5478
rect 27061 5264 35772 5266
rect 27061 5208 27066 5264
rect 27122 5208 35772 5264
rect 27061 5206 35772 5208
rect 17309 5203 17375 5206
rect 21541 5203 21607 5206
rect 27061 5203 27127 5206
rect 39520 5130 40000 5160
rect 17174 5070 40000 5130
rect 39520 5040 40000 5070
rect 16665 4994 16731 4997
rect 21541 4994 21607 4997
rect 16665 4992 21607 4994
rect 16665 4936 16670 4992
rect 16726 4936 21546 4992
rect 21602 4936 21607 4992
rect 16665 4934 21607 4936
rect 16665 4931 16731 4934
rect 21541 4931 21607 4934
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 27061 4858 27127 4861
rect 15518 4856 27127 4858
rect 15518 4800 27066 4856
rect 27122 4800 27127 4856
rect 15518 4798 27127 4800
rect 8201 4795 8267 4798
rect 14089 4795 14155 4798
rect 27061 4795 27127 4798
rect 2037 4722 2103 4725
rect 7465 4722 7531 4725
rect 26049 4722 26115 4725
rect 28257 4722 28323 4725
rect 2037 4720 7531 4722
rect 2037 4664 2042 4720
rect 2098 4664 7470 4720
rect 7526 4664 7531 4720
rect 2037 4662 7531 4664
rect 2037 4659 2103 4662
rect 7465 4659 7531 4662
rect 7606 4662 8218 4722
rect 0 4586 480 4616
rect 3877 4586 3943 4589
rect 7606 4586 7666 4662
rect 0 4584 3943 4586
rect 0 4528 3882 4584
rect 3938 4528 3943 4584
rect 0 4526 3943 4528
rect 0 4496 480 4526
rect 3877 4523 3943 4526
rect 7422 4526 7666 4586
rect 2313 4450 2379 4453
rect 7422 4450 7482 4526
rect 2313 4448 7482 4450
rect 2313 4392 2318 4448
rect 2374 4392 7482 4448
rect 2313 4390 7482 4392
rect 8158 4450 8218 4662
rect 26049 4720 28323 4722
rect 26049 4664 26054 4720
rect 26110 4664 28262 4720
rect 28318 4664 28323 4720
rect 26049 4662 28323 4664
rect 26049 4659 26115 4662
rect 28257 4659 28323 4662
rect 28942 4660 28948 4724
rect 29012 4722 29018 4724
rect 39520 4722 40000 4752
rect 29012 4662 40000 4722
rect 29012 4660 29018 4662
rect 39520 4632 40000 4662
rect 20713 4450 20779 4453
rect 8158 4448 20779 4450
rect 8158 4392 20718 4448
rect 20774 4392 20779 4448
rect 8158 4390 20779 4392
rect 2313 4387 2379 4390
rect 20713 4387 20779 4390
rect 21357 4450 21423 4453
rect 28942 4450 28948 4452
rect 21357 4448 28948 4450
rect 21357 4392 21362 4448
rect 21418 4392 28948 4448
rect 21357 4390 28948 4392
rect 21357 4387 21423 4390
rect 28942 4388 28948 4390
rect 29012 4388 29018 4452
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 3877 4314 3943 4317
rect 7373 4314 7439 4317
rect 3877 4312 7439 4314
rect 3877 4256 3882 4312
rect 3938 4256 7378 4312
rect 7434 4256 7439 4312
rect 3877 4254 7439 4256
rect 3877 4251 3943 4254
rect 7373 4251 7439 4254
rect 8017 4314 8083 4317
rect 16573 4314 16639 4317
rect 39520 4314 40000 4344
rect 8017 4312 16639 4314
rect 8017 4256 8022 4312
rect 8078 4256 16578 4312
rect 16634 4256 16639 4312
rect 8017 4254 16639 4256
rect 8017 4251 8083 4254
rect 16573 4251 16639 4254
rect 35712 4254 40000 4314
rect 0 4178 480 4208
rect 3785 4178 3851 4181
rect 0 4176 3851 4178
rect 0 4120 3790 4176
rect 3846 4120 3851 4176
rect 0 4118 3851 4120
rect 0 4088 480 4118
rect 3785 4115 3851 4118
rect 7465 4178 7531 4181
rect 35712 4178 35772 4254
rect 39520 4224 40000 4254
rect 7465 4176 35772 4178
rect 7465 4120 7470 4176
rect 7526 4120 35772 4176
rect 7465 4118 35772 4120
rect 7465 4115 7531 4118
rect 2037 4042 2103 4045
rect 21541 4042 21607 4045
rect 39520 4042 40000 4072
rect 2037 4040 21607 4042
rect 2037 3984 2042 4040
rect 2098 3984 21546 4040
rect 21602 3984 21607 4040
rect 2037 3982 21607 3984
rect 2037 3979 2103 3982
rect 21541 3979 21607 3982
rect 21774 3982 40000 4042
rect 3417 3906 3483 3909
rect 14089 3906 14155 3909
rect 3417 3904 14155 3906
rect 3417 3848 3422 3904
rect 3478 3848 14094 3904
rect 14150 3848 14155 3904
rect 3417 3846 14155 3848
rect 3417 3843 3483 3846
rect 14089 3843 14155 3846
rect 18597 3906 18663 3909
rect 21774 3906 21834 3982
rect 39520 3952 40000 3982
rect 18597 3904 21834 3906
rect 18597 3848 18602 3904
rect 18658 3848 21834 3904
rect 18597 3846 21834 3848
rect 28073 3906 28139 3909
rect 35341 3906 35407 3909
rect 28073 3904 35407 3906
rect 28073 3848 28078 3904
rect 28134 3848 35346 3904
rect 35402 3848 35407 3904
rect 28073 3846 35407 3848
rect 18597 3843 18663 3846
rect 28073 3843 28139 3846
rect 35341 3843 35407 3846
rect 14277 3840 14597 3841
rect 0 3770 480 3800
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 4061 3770 4127 3773
rect 0 3768 4127 3770
rect 0 3712 4066 3768
rect 4122 3712 4127 3768
rect 0 3710 4127 3712
rect 0 3680 480 3710
rect 4061 3707 4127 3710
rect 17217 3770 17283 3773
rect 27429 3770 27495 3773
rect 17217 3768 27495 3770
rect 17217 3712 17222 3768
rect 17278 3712 27434 3768
rect 27490 3712 27495 3768
rect 17217 3710 27495 3712
rect 17217 3707 17283 3710
rect 27429 3707 27495 3710
rect 28165 3770 28231 3773
rect 35801 3770 35867 3773
rect 28165 3768 35867 3770
rect 28165 3712 28170 3768
rect 28226 3712 35806 3768
rect 35862 3712 35867 3768
rect 28165 3710 35867 3712
rect 28165 3707 28231 3710
rect 35801 3707 35867 3710
rect 9857 3634 9923 3637
rect 21357 3634 21423 3637
rect 9857 3632 21423 3634
rect 9857 3576 9862 3632
rect 9918 3576 21362 3632
rect 21418 3576 21423 3632
rect 9857 3574 21423 3576
rect 9857 3571 9923 3574
rect 21357 3571 21423 3574
rect 21541 3634 21607 3637
rect 26693 3634 26759 3637
rect 21541 3632 26759 3634
rect 21541 3576 21546 3632
rect 21602 3576 26698 3632
rect 26754 3576 26759 3632
rect 21541 3574 26759 3576
rect 21541 3571 21607 3574
rect 26693 3571 26759 3574
rect 26877 3634 26943 3637
rect 39520 3634 40000 3664
rect 26877 3632 40000 3634
rect 26877 3576 26882 3632
rect 26938 3576 40000 3632
rect 26877 3574 40000 3576
rect 26877 3571 26943 3574
rect 39520 3544 40000 3574
rect 1669 3498 1735 3501
rect 1669 3496 35772 3498
rect 1669 3440 1674 3496
rect 1730 3440 35772 3496
rect 1669 3438 35772 3440
rect 1669 3435 1735 3438
rect 0 3362 480 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 480 3302
rect 3969 3299 4035 3302
rect 8569 3362 8635 3365
rect 17217 3362 17283 3365
rect 8569 3360 17283 3362
rect 8569 3304 8574 3360
rect 8630 3304 17222 3360
rect 17278 3304 17283 3360
rect 8569 3302 17283 3304
rect 8569 3299 8635 3302
rect 17217 3299 17283 3302
rect 21357 3362 21423 3365
rect 28073 3362 28139 3365
rect 21357 3360 28139 3362
rect 21357 3304 21362 3360
rect 21418 3304 28078 3360
rect 28134 3304 28139 3360
rect 21357 3302 28139 3304
rect 21357 3299 21423 3302
rect 28073 3299 28139 3302
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 26693 3226 26759 3229
rect 28073 3226 28139 3229
rect 26693 3224 28139 3226
rect 26693 3168 26698 3224
rect 26754 3168 28078 3224
rect 28134 3168 28139 3224
rect 26693 3166 28139 3168
rect 35712 3226 35772 3438
rect 39520 3226 40000 3256
rect 35712 3166 40000 3226
rect 26693 3163 26759 3166
rect 28073 3163 28139 3166
rect 39520 3136 40000 3166
rect 2681 3090 2747 3093
rect 28165 3090 28231 3093
rect 2681 3088 28231 3090
rect 2681 3032 2686 3088
rect 2742 3032 28170 3088
rect 28226 3032 28231 3088
rect 2681 3030 28231 3032
rect 2681 3027 2747 3030
rect 28165 3027 28231 3030
rect 28349 3090 28415 3093
rect 35433 3090 35499 3093
rect 28349 3088 35499 3090
rect 28349 3032 28354 3088
rect 28410 3032 35438 3088
rect 35494 3032 35499 3088
rect 28349 3030 35499 3032
rect 28349 3027 28415 3030
rect 35433 3027 35499 3030
rect 0 2954 480 2984
rect 3877 2954 3943 2957
rect 0 2952 3943 2954
rect 0 2896 3882 2952
rect 3938 2896 3943 2952
rect 0 2894 3943 2896
rect 0 2864 480 2894
rect 3877 2891 3943 2894
rect 4337 2954 4403 2957
rect 26877 2954 26943 2957
rect 4337 2952 26943 2954
rect 4337 2896 4342 2952
rect 4398 2896 26882 2952
rect 26938 2896 26943 2952
rect 4337 2894 26943 2896
rect 4337 2891 4403 2894
rect 26877 2891 26943 2894
rect 19977 2818 20043 2821
rect 25865 2818 25931 2821
rect 19977 2816 25931 2818
rect 19977 2760 19982 2816
rect 20038 2760 25870 2816
rect 25926 2760 25931 2816
rect 19977 2758 25931 2760
rect 19977 2755 20043 2758
rect 25865 2755 25931 2758
rect 28073 2818 28139 2821
rect 39520 2818 40000 2848
rect 28073 2816 40000 2818
rect 28073 2760 28078 2816
rect 28134 2760 40000 2816
rect 28073 2758 40000 2760
rect 28073 2755 28139 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 39520 2728 40000 2758
rect 27610 2687 27930 2688
rect 9673 2682 9739 2685
rect 3374 2680 9739 2682
rect 3374 2624 9678 2680
rect 9734 2624 9739 2680
rect 3374 2622 9739 2624
rect 0 2546 480 2576
rect 3374 2546 3434 2622
rect 9673 2619 9739 2622
rect 0 2486 3434 2546
rect 7465 2546 7531 2549
rect 8385 2546 8451 2549
rect 7465 2544 8451 2546
rect 7465 2488 7470 2544
rect 7526 2488 8390 2544
rect 8446 2488 8451 2544
rect 7465 2486 8451 2488
rect 0 2456 480 2486
rect 7465 2483 7531 2486
rect 8385 2483 8451 2486
rect 18965 2546 19031 2549
rect 18965 2544 35634 2546
rect 18965 2488 18970 2544
rect 19026 2488 35634 2544
rect 18965 2486 35634 2488
rect 18965 2483 19031 2486
rect 1577 2410 1643 2413
rect 34605 2410 34671 2413
rect 1577 2408 34671 2410
rect 1577 2352 1582 2408
rect 1638 2352 34610 2408
rect 34666 2352 34671 2408
rect 1577 2350 34671 2352
rect 1577 2347 1643 2350
rect 34605 2347 34671 2350
rect 7610 2208 7930 2209
rect 0 2138 480 2168
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 7465 2138 7531 2141
rect 0 2136 7531 2138
rect 0 2080 7470 2136
rect 7526 2080 7531 2136
rect 0 2078 7531 2080
rect 35574 2138 35634 2486
rect 35709 2410 35775 2413
rect 39520 2410 40000 2440
rect 35709 2408 40000 2410
rect 35709 2352 35714 2408
rect 35770 2352 40000 2408
rect 35709 2350 40000 2352
rect 35709 2347 35775 2350
rect 39520 2320 40000 2350
rect 39520 2138 40000 2168
rect 35574 2078 40000 2138
rect 0 2048 480 2078
rect 7465 2075 7531 2078
rect 39520 2048 40000 2078
rect 20805 2002 20871 2005
rect 3374 2000 20871 2002
rect 3374 1944 20810 2000
rect 20866 1944 20871 2000
rect 3374 1942 20871 1944
rect 0 1730 480 1760
rect 3374 1730 3434 1942
rect 20805 1939 20871 1942
rect 3693 1866 3759 1869
rect 18505 1866 18571 1869
rect 3693 1864 18571 1866
rect 3693 1808 3698 1864
rect 3754 1808 18510 1864
rect 18566 1808 18571 1864
rect 3693 1806 18571 1808
rect 3693 1803 3759 1806
rect 18505 1803 18571 1806
rect 0 1670 3434 1730
rect 21817 1730 21883 1733
rect 39520 1730 40000 1760
rect 21817 1728 40000 1730
rect 21817 1672 21822 1728
rect 21878 1672 40000 1728
rect 21817 1670 40000 1672
rect 0 1640 480 1670
rect 21817 1667 21883 1670
rect 39520 1640 40000 1670
rect 2037 1458 2103 1461
rect 35709 1458 35775 1461
rect 2037 1456 35775 1458
rect 2037 1400 2042 1456
rect 2098 1400 35714 1456
rect 35770 1400 35775 1456
rect 2037 1398 35775 1400
rect 2037 1395 2103 1398
rect 35709 1395 35775 1398
rect 0 1322 480 1352
rect 1393 1322 1459 1325
rect 0 1320 1459 1322
rect 0 1264 1398 1320
rect 1454 1264 1459 1320
rect 0 1262 1459 1264
rect 0 1232 480 1262
rect 1393 1259 1459 1262
rect 30465 1322 30531 1325
rect 39520 1322 40000 1352
rect 30465 1320 40000 1322
rect 30465 1264 30470 1320
rect 30526 1264 40000 1320
rect 30465 1262 40000 1264
rect 30465 1259 30531 1262
rect 39520 1232 40000 1262
rect 0 914 480 944
rect 3233 914 3299 917
rect 39520 914 40000 944
rect 0 912 3299 914
rect 0 856 3238 912
rect 3294 856 3299 912
rect 0 854 3299 856
rect 0 824 480 854
rect 3233 851 3299 854
rect 30974 854 40000 914
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
rect 17861 506 17927 509
rect 30833 506 30899 509
rect 17861 504 30899 506
rect 17861 448 17866 504
rect 17922 448 30838 504
rect 30894 448 30899 504
rect 17861 446 30899 448
rect 17861 443 17927 446
rect 30833 443 30899 446
rect 15469 370 15535 373
rect 30974 370 31034 854
rect 39520 824 40000 854
rect 31109 506 31175 509
rect 39520 506 40000 536
rect 31109 504 40000 506
rect 31109 448 31114 504
rect 31170 448 40000 504
rect 31109 446 40000 448
rect 31109 443 31175 446
rect 39520 416 40000 446
rect 15469 368 31034 370
rect 15469 312 15474 368
rect 15530 312 31034 368
rect 15469 310 31034 312
rect 15469 307 15535 310
rect 0 234 480 264
rect 3417 234 3483 237
rect 0 232 3483 234
rect 0 176 3422 232
rect 3478 176 3483 232
rect 0 174 3483 176
rect 0 144 480 174
rect 3417 171 3483 174
rect 4705 234 4771 237
rect 30833 234 30899 237
rect 39520 234 40000 264
rect 4705 232 30666 234
rect 4705 176 4710 232
rect 4766 176 30666 232
rect 4705 174 30666 176
rect 4705 171 4771 174
rect 3325 98 3391 101
rect 30465 98 30531 101
rect 3325 96 30531 98
rect 3325 40 3330 96
rect 3386 40 30470 96
rect 30526 40 30531 96
rect 3325 38 30531 40
rect 30606 98 30666 174
rect 30833 232 40000 234
rect 30833 176 30838 232
rect 30894 176 40000 232
rect 30833 174 40000 176
rect 30833 171 30899 174
rect 39520 144 40000 174
rect 31109 98 31175 101
rect 30606 96 31175 98
rect 30606 40 31114 96
rect 31170 40 31175 96
rect 30606 38 31175 40
rect 3325 35 3391 38
rect 30465 35 30531 38
rect 31109 35 31175 38
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 28948 4660 29012 4724
rect 28948 4388 29012 4452
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 28947 4724 29013 4725
rect 28947 4660 28948 4724
rect 29012 4660 29013 4724
rect 28947 4659 29013 4660
rect 28950 4453 29010 4659
rect 28947 4452 29013 4453
rect 28947 4388 28948 4452
rect 29012 4388 29013 4452
rect 28947 4387 29013 4388
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _30_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _13_
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _15_
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_25
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_35 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_40
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_52 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_60
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_78 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_215
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_290
timestamp 1586364061
transform 1 0 27784 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_302
timestamp 1586364061
transform 1 0 28888 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _11_
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _10_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_109
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_133
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _29_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_165
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_169
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_181
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _28_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_172
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _27_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_54
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_165
timestamp 1586364061
transform 1 0 16284 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_297
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_301
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_336
timestamp 1586364061
transform 1 0 32016 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_339
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_351
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_363
timestamp 1586364061
transform 1 0 34500 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _07_
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use scs8hd_buf_2  _08_
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _09_
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_192
timestamp 1586364061
transform 1 0 18768 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 28244 0 -1 5984
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_294
timestamp 1586364061
transform 1 0 28152 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_314
timestamp 1586364061
transform 1 0 29992 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _14_
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_326
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_334
timestamp 1586364061
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_336
timestamp 1586364061
transform 1 0 32016 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_341
timestamp 1586364061
transform 1 0 32476 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_353
timestamp 1586364061
transform 1 0 33580 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_341
timestamp 1586364061
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_345
timestamp 1586364061
transform 1 0 32844 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_357
timestamp 1586364061
transform 1 0 33948 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_365
timestamp 1586364061
transform 1 0 34684 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_365
timestamp 1586364061
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_377
timestamp 1586364061
transform 1 0 35788 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_389
timestamp 1586364061
transform 1 0 36892 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _25_
timestamp 1586364061
transform 1 0 1472 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_8
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_20
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_28
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__02__A
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_160
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 590 592
use scs8hd_buf_2  _02_
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__03__A
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_89
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _12_
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_336
timestamp 1586364061
transform 1 0 32016 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_341
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_357
timestamp 1586364061
transform 1 0 33948 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_365
timestamp 1586364061
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _04_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _03_
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_2  _05_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_109
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 29256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_308
timestamp 1586364061
transform 1 0 29440 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_320
timestamp 1586364061
transform 1 0 30544 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_332
timestamp 1586364061
transform 1 0 31648 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_373
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_385
timestamp 1586364061
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _01_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_224
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _06_
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_325
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 32660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_341
timestamp 1586364061
transform 1 0 32476 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_345
timestamp 1586364061
transform 1 0 32844 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_357
timestamp 1586364061
transform 1 0 33948 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_365
timestamp 1586364061
transform 1 0 34684 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_8
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_236
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_248
timestamp 1586364061
transform 1 0 23920 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_260
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_385
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _24_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  _26_
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_339
timestamp 1586364061
transform 1 0 32292 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_351
timestamp 1586364061
transform 1 0 33396 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_341
timestamp 1586364061
transform 1 0 32476 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_353
timestamp 1586364061
transform 1 0 33580 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_363
timestamp 1586364061
transform 1 0 34500 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_365
timestamp 1586364061
transform 1 0 34684 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_377
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_200
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_212
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_224
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_278
timestamp 1586364061
transform 1 0 26680 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_282
timestamp 1586364061
transform 1 0 27048 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_294
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_302
timestamp 1586364061
transform 1 0 28888 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_mux2_2  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_295
timestamp 1586364061
transform 1 0 28244 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_307
timestamp 1586364061
transform 1 0 29348 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_319
timestamp 1586364061
transform 1 0 30452 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_331
timestamp 1586364061
transform 1 0 31556 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_335
timestamp 1586364061
transform 1 0 31924 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 19982 0 20038 480 6 ccff_head
port 0 nsew default input
rlabel metal3 s 39520 15376 40000 15496 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 144 480 264 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 3272 480 3392 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 12112 480 12232 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 12928 480 13048 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 9664 480 9784 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 10072 480 10192 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 11296 480 11416 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 11704 480 11824 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 39520 144 40000 264 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 39520 4224 40000 4344 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 39520 4632 40000 4752 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 39520 5040 40000 5160 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 39520 5448 40000 5568 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 39520 5856 40000 5976 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 39520 6128 40000 6248 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 39520 6944 40000 7064 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 39520 7352 40000 7472 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 39520 824 40000 944 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 39520 1640 40000 1760 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 39520 2048 40000 2168 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 39520 2320 40000 2440 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 39520 2728 40000 2848 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 39520 3136 40000 3256 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 39520 3544 40000 3664 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 39520 7760 40000 7880 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 39520 11568 40000 11688 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 39520 12248 40000 12368 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 39520 12656 40000 12776 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 39520 13064 40000 13184 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 39520 13472 40000 13592 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 39520 13880 40000 14000 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 39520 14152 40000 14272 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 39520 14968 40000 15088 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 39520 8168 40000 8288 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 39520 8848 40000 8968 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 39520 9664 40000 9784 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 39520 10072 40000 10192 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 39520 10344 40000 10464 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 39520 10752 40000 10872 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 39520 11160 40000 11280 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal3 s 39520 15784 40000 15904 6 prog_clk
port 82 nsew default input
rlabel metal2 s 19982 15520 20038 16000 6 top_grid_pin_0_
port 83 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 84 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 85 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
