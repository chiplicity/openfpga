VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__1_
  CLASS BLOCK ;
  FOREIGN sb_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN bottom_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END bottom_left_grid_pin_42_
  PIN bottom_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 2.400 ;
    END
  END bottom_left_grid_pin_43_
  PIN bottom_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 2.400 ;
    END
  END bottom_left_grid_pin_44_
  PIN bottom_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END bottom_left_grid_pin_45_
  PIN bottom_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END bottom_left_grid_pin_46_
  PIN bottom_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.400 ;
    END
  END bottom_left_grid_pin_47_
  PIN bottom_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END bottom_left_grid_pin_48_
  PIN bottom_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END bottom_left_grid_pin_49_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 2.400 67.960 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.400 82.240 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 2.400 84.280 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 2.400 89.040 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 19.760 114.000 20.360 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 43.560 114.000 44.160 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 45.600 114.000 46.200 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 48.320 114.000 48.920 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 50.360 114.000 50.960 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 53.080 114.000 53.680 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 55.120 114.000 55.720 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 57.840 114.000 58.440 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 59.880 114.000 60.480 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 62.600 114.000 63.200 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 64.640 114.000 65.240 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 21.800 114.000 22.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 24.520 114.000 25.120 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 26.560 114.000 27.160 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 29.280 114.000 29.880 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 31.320 114.000 31.920 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 34.040 114.000 34.640 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 36.080 114.000 36.680 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 38.800 114.000 39.400 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 40.840 114.000 41.440 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 67.360 114.000 67.960 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 91.160 114.000 91.760 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 93.200 114.000 93.800 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 95.920 114.000 96.520 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 97.960 114.000 98.560 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 100.680 114.000 101.280 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 102.720 114.000 103.320 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 105.440 114.000 106.040 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 107.480 114.000 108.080 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 110.200 114.000 110.800 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 112.240 114.000 112.840 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 69.400 114.000 70.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 72.120 114.000 72.720 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 74.160 114.000 74.760 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 76.880 114.000 77.480 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 78.920 114.000 79.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 81.640 114.000 82.240 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 83.680 114.000 84.280 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 86.400 114.000 87.000 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 88.440 114.000 89.040 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 111.600 20.150 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 111.600 44.070 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 111.600 46.370 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 111.600 48.670 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 111.600 50.970 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 111.600 53.270 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 111.600 55.570 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 111.600 58.330 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 111.600 60.630 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 111.600 62.930 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 111.600 65.230 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 111.600 22.450 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 111.600 24.750 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 111.600 27.050 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 111.600 29.810 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 111.600 32.110 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 111.600 34.410 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 111.600 36.710 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 111.600 39.010 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 111.600 41.310 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 111.600 67.530 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 111.600 91.450 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 111.600 93.750 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 111.600 96.050 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 111.600 98.350 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 111.600 101.110 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 111.600 103.410 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 111.600 105.710 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 111.600 108.010 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.030 111.600 110.310 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 111.600 112.610 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 111.600 69.830 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 111.600 72.590 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 111.600 74.890 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 111.600 77.190 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 111.600 79.490 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 111.600 81.790 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 111.600 84.090 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 111.600 86.850 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 111.600 89.150 114.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END left_bottom_grid_pin_34_
  PIN left_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END left_bottom_grid_pin_35_
  PIN left_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.400 6.080 ;
    END
  END left_bottom_grid_pin_36_
  PIN left_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END left_bottom_grid_pin_37_
  PIN left_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END left_bottom_grid_pin_38_
  PIN left_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END left_bottom_grid_pin_39_
  PIN left_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END left_bottom_grid_pin_40_
  PIN left_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_bottom_grid_pin_41_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 2.760 114.000 3.360 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 5.480 114.000 6.080 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 7.520 114.000 8.120 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 10.240 114.000 10.840 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 12.280 114.000 12.880 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 15.000 114.000 15.600 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 17.040 114.000 17.640 ;
    END
  END right_bottom_grid_pin_41_
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 111.600 1.290 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 111.600 3.590 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 111.600 5.890 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 111.600 8.190 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 111.600 10.490 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 111.600 12.790 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 111.600 15.550 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 111.600 17.850 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 2.760 113.090 111.140 ;
      LAYER met2 ;
        RECT 1.570 111.320 3.030 112.725 ;
        RECT 3.870 111.320 5.330 112.725 ;
        RECT 6.170 111.320 7.630 112.725 ;
        RECT 8.470 111.320 9.930 112.725 ;
        RECT 10.770 111.320 12.230 112.725 ;
        RECT 13.070 111.320 14.990 112.725 ;
        RECT 15.830 111.320 17.290 112.725 ;
        RECT 18.130 111.320 19.590 112.725 ;
        RECT 20.430 111.320 21.890 112.725 ;
        RECT 22.730 111.320 24.190 112.725 ;
        RECT 25.030 111.320 26.490 112.725 ;
        RECT 27.330 111.320 29.250 112.725 ;
        RECT 30.090 111.320 31.550 112.725 ;
        RECT 32.390 111.320 33.850 112.725 ;
        RECT 34.690 111.320 36.150 112.725 ;
        RECT 36.990 111.320 38.450 112.725 ;
        RECT 39.290 111.320 40.750 112.725 ;
        RECT 41.590 111.320 43.510 112.725 ;
        RECT 44.350 111.320 45.810 112.725 ;
        RECT 46.650 111.320 48.110 112.725 ;
        RECT 48.950 111.320 50.410 112.725 ;
        RECT 51.250 111.320 52.710 112.725 ;
        RECT 53.550 111.320 55.010 112.725 ;
        RECT 55.850 111.320 57.770 112.725 ;
        RECT 58.610 111.320 60.070 112.725 ;
        RECT 60.910 111.320 62.370 112.725 ;
        RECT 63.210 111.320 64.670 112.725 ;
        RECT 65.510 111.320 66.970 112.725 ;
        RECT 67.810 111.320 69.270 112.725 ;
        RECT 70.110 111.320 72.030 112.725 ;
        RECT 72.870 111.320 74.330 112.725 ;
        RECT 75.170 111.320 76.630 112.725 ;
        RECT 77.470 111.320 78.930 112.725 ;
        RECT 79.770 111.320 81.230 112.725 ;
        RECT 82.070 111.320 83.530 112.725 ;
        RECT 84.370 111.320 86.290 112.725 ;
        RECT 87.130 111.320 88.590 112.725 ;
        RECT 89.430 111.320 90.890 112.725 ;
        RECT 91.730 111.320 93.190 112.725 ;
        RECT 94.030 111.320 95.490 112.725 ;
        RECT 96.330 111.320 97.790 112.725 ;
        RECT 98.630 111.320 100.550 112.725 ;
        RECT 101.390 111.320 102.850 112.725 ;
        RECT 103.690 111.320 105.150 112.725 ;
        RECT 105.990 111.320 107.450 112.725 ;
        RECT 108.290 111.320 109.750 112.725 ;
        RECT 110.590 111.320 112.050 112.725 ;
        RECT 112.890 111.320 113.060 112.725 ;
        RECT 1.020 2.680 113.060 111.320 ;
        RECT 1.570 0.835 2.570 2.680 ;
        RECT 3.410 0.835 4.870 2.680 ;
        RECT 5.710 0.835 7.170 2.680 ;
        RECT 8.010 0.835 9.470 2.680 ;
        RECT 10.310 0.835 11.770 2.680 ;
        RECT 12.610 0.835 14.070 2.680 ;
        RECT 14.910 0.835 16.370 2.680 ;
        RECT 17.210 0.835 18.210 2.680 ;
        RECT 19.050 0.835 20.510 2.680 ;
        RECT 21.350 0.835 22.810 2.680 ;
        RECT 23.650 0.835 25.110 2.680 ;
        RECT 25.950 0.835 27.410 2.680 ;
        RECT 28.250 0.835 29.710 2.680 ;
        RECT 30.550 0.835 32.010 2.680 ;
        RECT 32.850 0.835 33.850 2.680 ;
        RECT 34.690 0.835 36.150 2.680 ;
        RECT 36.990 0.835 38.450 2.680 ;
        RECT 39.290 0.835 40.750 2.680 ;
        RECT 41.590 0.835 43.050 2.680 ;
        RECT 43.890 0.835 45.350 2.680 ;
        RECT 46.190 0.835 47.650 2.680 ;
        RECT 48.490 0.835 49.490 2.680 ;
        RECT 50.330 0.835 51.790 2.680 ;
        RECT 52.630 0.835 54.090 2.680 ;
        RECT 54.930 0.835 56.390 2.680 ;
        RECT 57.230 0.835 58.690 2.680 ;
        RECT 59.530 0.835 60.990 2.680 ;
        RECT 61.830 0.835 63.290 2.680 ;
        RECT 64.130 0.835 65.590 2.680 ;
        RECT 66.430 0.835 67.430 2.680 ;
        RECT 68.270 0.835 69.730 2.680 ;
        RECT 70.570 0.835 72.030 2.680 ;
        RECT 72.870 0.835 74.330 2.680 ;
        RECT 75.170 0.835 76.630 2.680 ;
        RECT 77.470 0.835 78.930 2.680 ;
        RECT 79.770 0.835 81.230 2.680 ;
        RECT 82.070 0.835 83.070 2.680 ;
        RECT 83.910 0.835 85.370 2.680 ;
        RECT 86.210 0.835 87.670 2.680 ;
        RECT 88.510 0.835 89.970 2.680 ;
        RECT 90.810 0.835 92.270 2.680 ;
        RECT 93.110 0.835 94.570 2.680 ;
        RECT 95.410 0.835 96.870 2.680 ;
        RECT 97.710 0.835 98.710 2.680 ;
        RECT 99.550 0.835 101.010 2.680 ;
        RECT 101.850 0.835 103.310 2.680 ;
        RECT 104.150 0.835 105.610 2.680 ;
        RECT 106.450 0.835 107.910 2.680 ;
        RECT 108.750 0.835 110.210 2.680 ;
        RECT 111.050 0.835 112.510 2.680 ;
      LAYER met3 ;
        RECT 2.800 111.840 111.200 112.705 ;
        RECT 2.400 111.200 111.600 111.840 ;
        RECT 2.800 109.800 111.200 111.200 ;
        RECT 2.400 108.480 111.600 109.800 ;
        RECT 2.800 107.080 111.200 108.480 ;
        RECT 2.400 106.440 111.600 107.080 ;
        RECT 2.800 105.040 111.200 106.440 ;
        RECT 2.400 103.720 111.600 105.040 ;
        RECT 2.800 102.320 111.200 103.720 ;
        RECT 2.400 101.680 111.600 102.320 ;
        RECT 2.800 100.280 111.200 101.680 ;
        RECT 2.400 98.960 111.600 100.280 ;
        RECT 2.800 97.560 111.200 98.960 ;
        RECT 2.400 96.920 111.600 97.560 ;
        RECT 2.800 95.520 111.200 96.920 ;
        RECT 2.400 94.200 111.600 95.520 ;
        RECT 2.800 92.800 111.200 94.200 ;
        RECT 2.400 92.160 111.600 92.800 ;
        RECT 2.800 90.760 111.200 92.160 ;
        RECT 2.400 89.440 111.600 90.760 ;
        RECT 2.800 88.040 111.200 89.440 ;
        RECT 2.400 87.400 111.600 88.040 ;
        RECT 2.800 86.000 111.200 87.400 ;
        RECT 2.400 84.680 111.600 86.000 ;
        RECT 2.800 83.280 111.200 84.680 ;
        RECT 2.400 82.640 111.600 83.280 ;
        RECT 2.800 81.240 111.200 82.640 ;
        RECT 2.400 79.920 111.600 81.240 ;
        RECT 2.800 78.520 111.200 79.920 ;
        RECT 2.400 77.880 111.600 78.520 ;
        RECT 2.800 76.480 111.200 77.880 ;
        RECT 2.400 75.160 111.600 76.480 ;
        RECT 2.800 73.760 111.200 75.160 ;
        RECT 2.400 73.120 111.600 73.760 ;
        RECT 2.800 71.720 111.200 73.120 ;
        RECT 2.400 70.400 111.600 71.720 ;
        RECT 2.800 69.000 111.200 70.400 ;
        RECT 2.400 68.360 111.600 69.000 ;
        RECT 2.800 66.960 111.200 68.360 ;
        RECT 2.400 65.640 111.600 66.960 ;
        RECT 2.800 64.240 111.200 65.640 ;
        RECT 2.400 63.600 111.600 64.240 ;
        RECT 2.800 62.200 111.200 63.600 ;
        RECT 2.400 60.880 111.600 62.200 ;
        RECT 2.800 59.480 111.200 60.880 ;
        RECT 2.400 58.840 111.600 59.480 ;
        RECT 2.800 57.440 111.200 58.840 ;
        RECT 2.400 56.120 111.600 57.440 ;
        RECT 2.800 54.720 111.200 56.120 ;
        RECT 2.400 54.080 111.600 54.720 ;
        RECT 2.800 52.680 111.200 54.080 ;
        RECT 2.400 51.360 111.600 52.680 ;
        RECT 2.800 49.960 111.200 51.360 ;
        RECT 2.400 49.320 111.600 49.960 ;
        RECT 2.800 47.920 111.200 49.320 ;
        RECT 2.400 46.600 111.600 47.920 ;
        RECT 2.800 45.200 111.200 46.600 ;
        RECT 2.400 44.560 111.600 45.200 ;
        RECT 2.800 43.160 111.200 44.560 ;
        RECT 2.400 41.840 111.600 43.160 ;
        RECT 2.800 40.440 111.200 41.840 ;
        RECT 2.400 39.800 111.600 40.440 ;
        RECT 2.800 38.400 111.200 39.800 ;
        RECT 2.400 37.080 111.600 38.400 ;
        RECT 2.800 35.680 111.200 37.080 ;
        RECT 2.400 35.040 111.600 35.680 ;
        RECT 2.800 33.640 111.200 35.040 ;
        RECT 2.400 32.320 111.600 33.640 ;
        RECT 2.800 30.920 111.200 32.320 ;
        RECT 2.400 30.280 111.600 30.920 ;
        RECT 2.800 28.880 111.200 30.280 ;
        RECT 2.400 27.560 111.600 28.880 ;
        RECT 2.800 26.160 111.200 27.560 ;
        RECT 2.400 25.520 111.600 26.160 ;
        RECT 2.800 24.120 111.200 25.520 ;
        RECT 2.400 22.800 111.600 24.120 ;
        RECT 2.800 21.400 111.200 22.800 ;
        RECT 2.400 20.760 111.600 21.400 ;
        RECT 2.800 19.360 111.200 20.760 ;
        RECT 2.400 18.040 111.600 19.360 ;
        RECT 2.800 16.640 111.200 18.040 ;
        RECT 2.400 16.000 111.600 16.640 ;
        RECT 2.800 14.600 111.200 16.000 ;
        RECT 2.400 13.280 111.600 14.600 ;
        RECT 2.800 11.880 111.200 13.280 ;
        RECT 2.400 11.240 111.600 11.880 ;
        RECT 2.800 9.840 111.200 11.240 ;
        RECT 2.400 8.520 111.600 9.840 ;
        RECT 2.800 7.120 111.200 8.520 ;
        RECT 2.400 6.480 111.600 7.120 ;
        RECT 2.800 5.080 111.200 6.480 ;
        RECT 2.400 3.760 111.600 5.080 ;
        RECT 2.800 2.360 111.200 3.760 ;
        RECT 2.400 1.720 111.600 2.360 ;
        RECT 2.800 0.855 111.200 1.720 ;
      LAYER met4 ;
        RECT 20.535 101.280 102.745 101.825 ;
        RECT 20.535 10.240 21.480 101.280 ;
        RECT 23.880 10.240 38.640 101.280 ;
        RECT 41.040 10.240 102.745 101.280 ;
        RECT 20.535 9.015 102.745 10.240 ;
  END
END sb_1__1_
END LIBRARY

