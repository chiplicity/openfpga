magic
tech EFS8A
magscale 1 2
timestamp 1604431043
<< viali >>
rect 3249 32521 3283 32555
rect 4353 32521 4387 32555
rect 7481 32521 7515 32555
rect 9597 32521 9631 32555
rect 10701 32521 10735 32555
rect 13093 32521 13127 32555
rect 3065 32317 3099 32351
rect 3617 32317 3651 32351
rect 4169 32317 4203 32351
rect 4721 32317 4755 32351
rect 6837 32317 6871 32351
rect 8953 32317 8987 32351
rect 10057 32317 10091 32351
rect 12449 32317 12483 32351
rect 7021 32181 7055 32215
rect 9137 32181 9171 32215
rect 10241 32181 10275 32215
rect 12633 32181 12667 32215
rect 1869 31977 1903 32011
rect 2973 31977 3007 32011
rect 4261 31977 4295 32011
rect 5549 31977 5583 32011
rect 6653 31977 6687 32011
rect 8033 31977 8067 32011
rect 9873 31977 9907 32011
rect 12541 31977 12575 32011
rect 1685 31841 1719 31875
rect 2789 31841 2823 31875
rect 4077 31841 4111 31875
rect 5365 31841 5399 31875
rect 6469 31841 6503 31875
rect 7849 31841 7883 31875
rect 9689 31841 9723 31875
rect 12357 31841 12391 31875
rect 13461 31841 13495 31875
rect 13645 31637 13679 31671
rect 2881 31433 2915 31467
rect 5089 31433 5123 31467
rect 6469 31433 6503 31467
rect 7021 31433 7055 31467
rect 13461 31433 13495 31467
rect 3985 31365 4019 31399
rect 9689 31365 9723 31399
rect 2697 31229 2731 31263
rect 3801 31229 3835 31263
rect 4905 31229 4939 31263
rect 6837 31229 6871 31263
rect 9505 31229 9539 31263
rect 12265 31229 12299 31263
rect 12449 31229 12483 31263
rect 1685 31093 1719 31127
rect 2513 31093 2547 31127
rect 3249 31093 3283 31127
rect 3617 31093 3651 31127
rect 4353 31093 4387 31127
rect 4721 31093 4755 31127
rect 5549 31093 5583 31127
rect 7389 31093 7423 31127
rect 7849 31093 7883 31127
rect 10057 31093 10091 31127
rect 10517 31093 10551 31127
rect 12633 31093 12667 31127
rect 13001 31093 13035 31127
rect 4077 30753 4111 30787
rect 9873 30753 9907 30787
rect 10057 30617 10091 30651
rect 4261 30549 4295 30583
rect 4077 30345 4111 30379
rect 9781 30277 9815 30311
rect 9873 30141 9907 30175
rect 11161 30141 11195 30175
rect 10057 30005 10091 30039
rect 10517 30005 10551 30039
rect 11345 30005 11379 30039
rect 11805 30005 11839 30039
rect 11161 29665 11195 29699
rect 11345 29461 11379 29495
rect 11161 29257 11195 29291
rect 10517 28713 10551 28747
rect 10333 28577 10367 28611
rect 10241 28169 10275 28203
rect 10333 27965 10367 27999
rect 6837 27829 6871 27863
rect 10517 27829 10551 27863
rect 10885 27829 10919 27863
rect 6929 27557 6963 27591
rect 7021 27421 7055 27455
rect 7205 27421 7239 27455
rect 6561 27285 6595 27319
rect 1593 27081 1627 27115
rect 5917 27081 5951 27115
rect 6285 27013 6319 27047
rect 7389 26945 7423 26979
rect 7849 26945 7883 26979
rect 1409 26877 1443 26911
rect 6653 26877 6687 26911
rect 7297 26877 7331 26911
rect 1961 26741 1995 26775
rect 6837 26741 6871 26775
rect 7205 26741 7239 26775
rect 5365 26537 5399 26571
rect 6929 26537 6963 26571
rect 5273 26469 5307 26503
rect 5457 26333 5491 26367
rect 4905 26265 4939 26299
rect 7205 26265 7239 26299
rect 4997 25993 5031 26027
rect 5365 25993 5399 26027
rect 5641 25993 5675 26027
rect 3249 25449 3283 25483
rect 12265 25449 12299 25483
rect 12081 25313 12115 25347
rect 3709 24769 3743 24803
rect 3617 24701 3651 24735
rect 2973 24565 3007 24599
rect 3157 24565 3191 24599
rect 3525 24565 3559 24599
rect 12081 24565 12115 24599
rect 3249 24021 3283 24055
rect 4537 21845 4571 21879
rect 4445 21641 4479 21675
rect 4997 21505 5031 21539
rect 4353 21369 4387 21403
rect 4813 21301 4847 21335
rect 4905 21301 4939 21335
rect 5917 21097 5951 21131
rect 6285 20961 6319 20995
rect 6377 20961 6411 20995
rect 6469 20893 6503 20927
rect 4537 20757 4571 20791
rect 6377 20553 6411 20587
rect 9597 20553 9631 20587
rect 8217 20349 8251 20383
rect 5641 20281 5675 20315
rect 8484 20281 8518 20315
rect 5917 20213 5951 20247
rect 8125 20213 8159 20247
rect 5641 20009 5675 20043
rect 7205 20009 7239 20043
rect 5549 19873 5583 19907
rect 6009 19873 6043 19907
rect 7573 19873 7607 19907
rect 7665 19873 7699 19907
rect 9781 19873 9815 19907
rect 10048 19873 10082 19907
rect 6101 19805 6135 19839
rect 6193 19805 6227 19839
rect 7849 19805 7883 19839
rect 6929 19669 6963 19703
rect 8309 19669 8343 19703
rect 11161 19669 11195 19703
rect 6837 19465 6871 19499
rect 10149 19465 10183 19499
rect 7481 19329 7515 19363
rect 3893 19261 3927 19295
rect 3985 19261 4019 19295
rect 4252 19261 4286 19295
rect 6285 19261 6319 19295
rect 3525 19193 3559 19227
rect 6653 19193 6687 19227
rect 7297 19193 7331 19227
rect 5365 19125 5399 19159
rect 7205 19125 7239 19159
rect 7849 19125 7883 19159
rect 9873 19125 9907 19159
rect 5733 18921 5767 18955
rect 6101 18921 6135 18955
rect 6285 18921 6319 18955
rect 7757 18921 7791 18955
rect 6653 18785 6687 18819
rect 6745 18717 6779 18751
rect 6929 18717 6963 18751
rect 7297 18581 7331 18615
rect 4537 18377 4571 18411
rect 6009 18377 6043 18411
rect 3065 18241 3099 18275
rect 3157 18241 3191 18275
rect 3402 18105 3436 18139
rect 7021 18105 7055 18139
rect 6377 18037 6411 18071
rect 3249 17833 3283 17867
rect 9965 14229 9999 14263
rect 9781 14025 9815 14059
rect 9873 13889 9907 13923
rect 10140 13821 10174 13855
rect 11253 13685 11287 13719
rect 9965 13481 9999 13515
rect 10333 13345 10367 13379
rect 10425 13277 10459 13311
rect 10517 13277 10551 13311
rect 10057 12937 10091 12971
rect 10701 12733 10735 12767
rect 10333 12597 10367 12631
rect 7757 12053 7791 12087
rect 9321 12053 9355 12087
rect 7757 11849 7791 11883
rect 9321 11849 9355 11883
rect 8309 11713 8343 11747
rect 9229 11713 9263 11747
rect 9965 11713 9999 11747
rect 9689 11645 9723 11679
rect 8217 11577 8251 11611
rect 7665 11509 7699 11543
rect 8125 11509 8159 11543
rect 9781 11509 9815 11543
rect 6929 11169 6963 11203
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 7757 11101 7791 11135
rect 6561 11033 6595 11067
rect 9321 11033 9355 11067
rect 6837 10761 6871 10795
rect 5917 10693 5951 10727
rect 7389 10625 7423 10659
rect 7849 10557 7883 10591
rect 8217 10489 8251 10523
rect 6193 10421 6227 10455
rect 6653 10421 6687 10455
rect 7205 10421 7239 10455
rect 7297 10421 7331 10455
rect 7297 10217 7331 10251
rect 7757 10217 7791 10251
rect 6101 10081 6135 10115
rect 7665 10081 7699 10115
rect 6193 10013 6227 10047
rect 6377 10013 6411 10047
rect 7849 10013 7883 10047
rect 5733 9945 5767 9979
rect 6929 9877 6963 9911
rect 6101 9673 6135 9707
rect 7665 9673 7699 9707
rect 8033 9673 8067 9707
rect 6469 9401 6503 9435
rect 5825 9333 5859 9367
rect 7389 9333 7423 9367
rect 4333 6817 4367 6851
rect 4077 6749 4111 6783
rect 5457 6613 5491 6647
rect 9965 6613 9999 6647
rect 4169 6409 4203 6443
rect 9873 6409 9907 6443
rect 9781 6341 9815 6375
rect 10333 6273 10367 6307
rect 10517 6273 10551 6307
rect 9413 6137 9447 6171
rect 10241 6137 10275 6171
rect 4537 6069 4571 6103
rect 9229 5865 9263 5899
rect 9873 5865 9907 5899
rect 10241 5797 10275 5831
rect 10333 5729 10367 5763
rect 10425 5661 10459 5695
rect 9137 5321 9171 5355
rect 10609 5321 10643 5355
rect 9229 5117 9263 5151
rect 9485 5117 9519 5151
rect 11161 4981 11195 5015
rect 7757 4777 7791 4811
rect 9321 4777 9355 4811
rect 10149 4777 10183 4811
rect 10609 4777 10643 4811
rect 6644 4709 6678 4743
rect 9965 4709 9999 4743
rect 6377 4641 6411 4675
rect 10517 4641 10551 4675
rect 10701 4573 10735 4607
rect 6469 4233 6503 4267
rect 9781 4233 9815 4267
rect 10793 4233 10827 4267
rect 7021 4097 7055 4131
rect 10333 4097 10367 4131
rect 10241 4029 10275 4063
rect 4077 3553 4111 3587
rect 5181 3553 5215 3587
rect 6285 3553 6319 3587
rect 4261 3417 4295 3451
rect 5365 3349 5399 3383
rect 6469 3349 6503 3383
rect 3433 3145 3467 3179
rect 3893 3145 3927 3179
rect 4169 3145 4203 3179
rect 4997 3145 5031 3179
rect 5733 3145 5767 3179
rect 6377 3145 6411 3179
rect 7941 3145 7975 3179
rect 5273 3077 5307 3111
rect 4629 3009 4663 3043
rect 2881 2941 2915 2975
rect 3985 2941 4019 2975
rect 5089 2941 5123 2975
rect 7297 2941 7331 2975
rect 3065 2805 3099 2839
rect 7481 2805 7515 2839
rect 3065 2601 3099 2635
rect 3433 2601 3467 2635
rect 4261 2601 4295 2635
rect 5825 2601 5859 2635
rect 7481 2601 7515 2635
rect 7941 2601 7975 2635
rect 1409 2465 1443 2499
rect 1961 2465 1995 2499
rect 2881 2465 2915 2499
rect 4077 2465 4111 2499
rect 4721 2465 4755 2499
rect 5181 2465 5215 2499
rect 7297 2465 7331 2499
rect 1593 2261 1627 2295
rect 5365 2261 5399 2295
<< metal1 >>
rect 13814 37748 13820 37800
rect 13872 37788 13878 37800
rect 14550 37788 14556 37800
rect 13872 37760 14556 37788
rect 13872 37748 13878 37760
rect 14550 37748 14556 37760
rect 14608 37748 14614 37800
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 198 34484 204 34536
rect 256 34524 262 34536
rect 1302 34524 1308 34536
rect 256 34496 1308 34524
rect 256 34484 262 34496
rect 1302 34484 1308 34496
rect 1360 34484 1366 34536
rect 1394 34484 1400 34536
rect 1452 34524 1458 34536
rect 2774 34524 2780 34536
rect 1452 34496 2780 34524
rect 1452 34484 1458 34496
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 2958 34484 2964 34536
rect 3016 34524 3022 34536
rect 4062 34524 4068 34536
rect 3016 34496 4068 34524
rect 3016 34484 3022 34496
rect 4062 34484 4068 34496
rect 4120 34484 4126 34536
rect 4154 34484 4160 34536
rect 4212 34524 4218 34536
rect 5534 34524 5540 34536
rect 4212 34496 5540 34524
rect 4212 34484 4218 34496
rect 5534 34484 5540 34496
rect 5592 34484 5598 34536
rect 7742 34484 7748 34536
rect 7800 34524 7806 34536
rect 8202 34524 8208 34536
rect 7800 34496 8208 34524
rect 7800 34484 7806 34496
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 2774 32512 2780 32564
rect 2832 32552 2838 32564
rect 3237 32555 3295 32561
rect 3237 32552 3249 32555
rect 2832 32524 3249 32552
rect 2832 32512 2838 32524
rect 3237 32521 3249 32524
rect 3283 32521 3295 32555
rect 3237 32515 3295 32521
rect 4154 32512 4160 32564
rect 4212 32552 4218 32564
rect 4341 32555 4399 32561
rect 4341 32552 4353 32555
rect 4212 32524 4353 32552
rect 4212 32512 4218 32524
rect 4341 32521 4353 32524
rect 4387 32521 4399 32555
rect 7466 32552 7472 32564
rect 7427 32524 7472 32552
rect 4341 32515 4399 32521
rect 7466 32512 7472 32524
rect 7524 32512 7530 32564
rect 9582 32552 9588 32564
rect 9543 32524 9588 32552
rect 9582 32512 9588 32524
rect 9640 32512 9646 32564
rect 10686 32552 10692 32564
rect 10647 32524 10692 32552
rect 10686 32512 10692 32524
rect 10744 32512 10750 32564
rect 13078 32552 13084 32564
rect 13039 32524 13084 32552
rect 13078 32512 13084 32524
rect 13136 32512 13142 32564
rect 3050 32348 3056 32360
rect 3011 32320 3056 32348
rect 3050 32308 3056 32320
rect 3108 32348 3114 32360
rect 3605 32351 3663 32357
rect 3605 32348 3617 32351
rect 3108 32320 3617 32348
rect 3108 32308 3114 32320
rect 3605 32317 3617 32320
rect 3651 32317 3663 32351
rect 3605 32311 3663 32317
rect 4157 32351 4215 32357
rect 4157 32317 4169 32351
rect 4203 32348 4215 32351
rect 4430 32348 4436 32360
rect 4203 32320 4436 32348
rect 4203 32317 4215 32320
rect 4157 32311 4215 32317
rect 4430 32308 4436 32320
rect 4488 32348 4494 32360
rect 4709 32351 4767 32357
rect 4709 32348 4721 32351
rect 4488 32320 4721 32348
rect 4488 32308 4494 32320
rect 4709 32317 4721 32320
rect 4755 32317 4767 32351
rect 4709 32311 4767 32317
rect 6825 32351 6883 32357
rect 6825 32317 6837 32351
rect 6871 32317 6883 32351
rect 6825 32311 6883 32317
rect 8941 32351 8999 32357
rect 8941 32317 8953 32351
rect 8987 32348 8999 32351
rect 9582 32348 9588 32360
rect 8987 32320 9588 32348
rect 8987 32317 8999 32320
rect 8941 32311 8999 32317
rect 6840 32280 6868 32311
rect 9582 32308 9588 32320
rect 9640 32308 9646 32360
rect 10045 32351 10103 32357
rect 10045 32317 10057 32351
rect 10091 32348 10103 32351
rect 10686 32348 10692 32360
rect 10091 32320 10692 32348
rect 10091 32317 10103 32320
rect 10045 32311 10103 32317
rect 10686 32308 10692 32320
rect 10744 32308 10750 32360
rect 12437 32351 12495 32357
rect 12437 32317 12449 32351
rect 12483 32348 12495 32351
rect 13078 32348 13084 32360
rect 12483 32320 13084 32348
rect 12483 32317 12495 32320
rect 12437 32311 12495 32317
rect 13078 32308 13084 32320
rect 13136 32308 13142 32360
rect 7466 32280 7472 32292
rect 6840 32252 7472 32280
rect 7466 32240 7472 32252
rect 7524 32240 7530 32292
rect 7009 32215 7067 32221
rect 7009 32181 7021 32215
rect 7055 32212 7067 32215
rect 7282 32212 7288 32224
rect 7055 32184 7288 32212
rect 7055 32181 7067 32184
rect 7009 32175 7067 32181
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 8846 32172 8852 32224
rect 8904 32212 8910 32224
rect 9125 32215 9183 32221
rect 9125 32212 9137 32215
rect 8904 32184 9137 32212
rect 8904 32172 8910 32184
rect 9125 32181 9137 32184
rect 9171 32181 9183 32215
rect 9125 32175 9183 32181
rect 9674 32172 9680 32224
rect 9732 32212 9738 32224
rect 10229 32215 10287 32221
rect 10229 32212 10241 32215
rect 9732 32184 10241 32212
rect 9732 32172 9738 32184
rect 10229 32181 10241 32184
rect 10275 32181 10287 32215
rect 12618 32212 12624 32224
rect 12579 32184 12624 32212
rect 10229 32175 10287 32181
rect 12618 32172 12624 32184
rect 12676 32172 12682 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1394 31968 1400 32020
rect 1452 32008 1458 32020
rect 1857 32011 1915 32017
rect 1857 32008 1869 32011
rect 1452 31980 1869 32008
rect 1452 31968 1458 31980
rect 1857 31977 1869 31980
rect 1903 31977 1915 32011
rect 1857 31971 1915 31977
rect 2866 31968 2872 32020
rect 2924 32008 2930 32020
rect 2961 32011 3019 32017
rect 2961 32008 2973 32011
rect 2924 31980 2973 32008
rect 2924 31968 2930 31980
rect 2961 31977 2973 31980
rect 3007 31977 3019 32011
rect 2961 31971 3019 31977
rect 4249 32011 4307 32017
rect 4249 31977 4261 32011
rect 4295 32008 4307 32011
rect 4338 32008 4344 32020
rect 4295 31980 4344 32008
rect 4295 31977 4307 31980
rect 4249 31971 4307 31977
rect 4338 31968 4344 31980
rect 4396 31968 4402 32020
rect 5534 32008 5540 32020
rect 5495 31980 5540 32008
rect 5534 31968 5540 31980
rect 5592 31968 5598 32020
rect 6641 32011 6699 32017
rect 6641 31977 6653 32011
rect 6687 32008 6699 32011
rect 6822 32008 6828 32020
rect 6687 31980 6828 32008
rect 6687 31977 6699 31980
rect 6641 31971 6699 31977
rect 6822 31968 6828 31980
rect 6880 31968 6886 32020
rect 8018 32008 8024 32020
rect 7979 31980 8024 32008
rect 8018 31968 8024 31980
rect 8076 31968 8082 32020
rect 9858 32008 9864 32020
rect 9819 31980 9864 32008
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 12526 32008 12532 32020
rect 12487 31980 12532 32008
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 1670 31872 1676 31884
rect 1631 31844 1676 31872
rect 1670 31832 1676 31844
rect 1728 31832 1734 31884
rect 2777 31875 2835 31881
rect 2777 31841 2789 31875
rect 2823 31872 2835 31875
rect 3234 31872 3240 31884
rect 2823 31844 3240 31872
rect 2823 31841 2835 31844
rect 2777 31835 2835 31841
rect 3234 31832 3240 31844
rect 3292 31832 3298 31884
rect 4065 31875 4123 31881
rect 4065 31841 4077 31875
rect 4111 31841 4123 31875
rect 4065 31835 4123 31841
rect 5353 31875 5411 31881
rect 5353 31841 5365 31875
rect 5399 31872 5411 31875
rect 5442 31872 5448 31884
rect 5399 31844 5448 31872
rect 5399 31841 5411 31844
rect 5353 31835 5411 31841
rect 4080 31736 4108 31835
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 6454 31872 6460 31884
rect 6415 31844 6460 31872
rect 6454 31832 6460 31844
rect 6512 31832 6518 31884
rect 7834 31872 7840 31884
rect 7795 31844 7840 31872
rect 7834 31832 7840 31844
rect 7892 31832 7898 31884
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31872 9735 31875
rect 10502 31872 10508 31884
rect 9723 31844 10508 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 10502 31832 10508 31844
rect 10560 31832 10566 31884
rect 12345 31875 12403 31881
rect 12345 31841 12357 31875
rect 12391 31841 12403 31875
rect 13446 31872 13452 31884
rect 13407 31844 13452 31872
rect 12345 31835 12403 31841
rect 7282 31764 7288 31816
rect 7340 31804 7346 31816
rect 7742 31804 7748 31816
rect 7340 31776 7748 31804
rect 7340 31764 7346 31776
rect 7742 31764 7748 31776
rect 7800 31764 7806 31816
rect 4338 31736 4344 31748
rect 4080 31708 4344 31736
rect 4338 31696 4344 31708
rect 4396 31696 4402 31748
rect 12360 31736 12388 31835
rect 13446 31832 13452 31844
rect 13504 31832 13510 31884
rect 12986 31736 12992 31748
rect 12360 31708 12992 31736
rect 12986 31696 12992 31708
rect 13044 31696 13050 31748
rect 13630 31668 13636 31680
rect 13591 31640 13636 31668
rect 13630 31628 13636 31640
rect 13688 31628 13694 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 2866 31464 2872 31476
rect 2827 31436 2872 31464
rect 2866 31424 2872 31436
rect 2924 31424 2930 31476
rect 4522 31424 4528 31476
rect 4580 31464 4586 31476
rect 5077 31467 5135 31473
rect 5077 31464 5089 31467
rect 4580 31436 5089 31464
rect 4580 31424 4586 31436
rect 5077 31433 5089 31436
rect 5123 31433 5135 31467
rect 6454 31464 6460 31476
rect 6415 31436 6460 31464
rect 5077 31427 5135 31433
rect 6454 31424 6460 31436
rect 6512 31424 6518 31476
rect 7006 31464 7012 31476
rect 6967 31436 7012 31464
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 13446 31464 13452 31476
rect 13407 31436 13452 31464
rect 13446 31424 13452 31436
rect 13504 31424 13510 31476
rect 2130 31356 2136 31408
rect 2188 31396 2194 31408
rect 3973 31399 4031 31405
rect 3973 31396 3985 31399
rect 2188 31368 3985 31396
rect 2188 31356 2194 31368
rect 3973 31365 3985 31368
rect 4019 31365 4031 31399
rect 9674 31396 9680 31408
rect 9635 31368 9680 31396
rect 3973 31359 4031 31365
rect 9674 31356 9680 31368
rect 9732 31356 9738 31408
rect 2685 31263 2743 31269
rect 2685 31260 2697 31263
rect 2516 31232 2697 31260
rect 2516 31136 2544 31232
rect 2685 31229 2697 31232
rect 2731 31229 2743 31263
rect 3789 31263 3847 31269
rect 3789 31260 3801 31263
rect 2685 31223 2743 31229
rect 3620 31232 3801 31260
rect 1670 31124 1676 31136
rect 1631 31096 1676 31124
rect 1670 31084 1676 31096
rect 1728 31084 1734 31136
rect 2498 31124 2504 31136
rect 2459 31096 2504 31124
rect 2498 31084 2504 31096
rect 2556 31084 2562 31136
rect 3234 31124 3240 31136
rect 3195 31096 3240 31124
rect 3234 31084 3240 31096
rect 3292 31084 3298 31136
rect 3418 31084 3424 31136
rect 3476 31124 3482 31136
rect 3620 31133 3648 31232
rect 3789 31229 3801 31232
rect 3835 31229 3847 31263
rect 4893 31263 4951 31269
rect 4893 31260 4905 31263
rect 3789 31223 3847 31229
rect 4724 31232 4905 31260
rect 4724 31136 4752 31232
rect 4893 31229 4905 31232
rect 4939 31229 4951 31263
rect 4893 31223 4951 31229
rect 6825 31263 6883 31269
rect 6825 31229 6837 31263
rect 6871 31260 6883 31263
rect 9493 31263 9551 31269
rect 6871 31232 7420 31260
rect 6871 31229 6883 31232
rect 6825 31223 6883 31229
rect 7392 31136 7420 31232
rect 9493 31229 9505 31263
rect 9539 31260 9551 31263
rect 12253 31263 12311 31269
rect 9539 31232 9996 31260
rect 9539 31229 9551 31232
rect 9493 31223 9551 31229
rect 9968 31136 9996 31232
rect 12253 31229 12265 31263
rect 12299 31260 12311 31263
rect 12437 31263 12495 31269
rect 12437 31260 12449 31263
rect 12299 31232 12449 31260
rect 12299 31229 12311 31232
rect 12253 31223 12311 31229
rect 12437 31229 12449 31232
rect 12483 31260 12495 31263
rect 13906 31260 13912 31272
rect 12483 31232 13912 31260
rect 12483 31229 12495 31232
rect 12437 31223 12495 31229
rect 13906 31220 13912 31232
rect 13964 31220 13970 31272
rect 3605 31127 3663 31133
rect 3605 31124 3617 31127
rect 3476 31096 3617 31124
rect 3476 31084 3482 31096
rect 3605 31093 3617 31096
rect 3651 31093 3663 31127
rect 4338 31124 4344 31136
rect 4299 31096 4344 31124
rect 3605 31087 3663 31093
rect 4338 31084 4344 31096
rect 4396 31084 4402 31136
rect 4706 31124 4712 31136
rect 4667 31096 4712 31124
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 5534 31124 5540 31136
rect 5495 31096 5540 31124
rect 5534 31084 5540 31096
rect 5592 31084 5598 31136
rect 7374 31124 7380 31136
rect 7335 31096 7380 31124
rect 7374 31084 7380 31096
rect 7432 31084 7438 31136
rect 7834 31124 7840 31136
rect 7795 31096 7840 31124
rect 7834 31084 7840 31096
rect 7892 31084 7898 31136
rect 9950 31084 9956 31136
rect 10008 31124 10014 31136
rect 10045 31127 10103 31133
rect 10045 31124 10057 31127
rect 10008 31096 10057 31124
rect 10008 31084 10014 31096
rect 10045 31093 10057 31096
rect 10091 31093 10103 31127
rect 10502 31124 10508 31136
rect 10415 31096 10508 31124
rect 10045 31087 10103 31093
rect 10502 31084 10508 31096
rect 10560 31124 10566 31136
rect 10962 31124 10968 31136
rect 10560 31096 10968 31124
rect 10560 31084 10566 31096
rect 10962 31084 10968 31096
rect 11020 31084 11026 31136
rect 12526 31084 12532 31136
rect 12584 31124 12590 31136
rect 12621 31127 12679 31133
rect 12621 31124 12633 31127
rect 12584 31096 12633 31124
rect 12584 31084 12590 31096
rect 12621 31093 12633 31096
rect 12667 31093 12679 31127
rect 12986 31124 12992 31136
rect 12947 31096 12992 31124
rect 12621 31087 12679 31093
rect 12986 31084 12992 31096
rect 13044 31084 13050 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 7466 30880 7472 30932
rect 7524 30920 7530 30932
rect 8110 30920 8116 30932
rect 7524 30892 8116 30920
rect 7524 30880 7530 30892
rect 8110 30880 8116 30892
rect 8168 30880 8174 30932
rect 4062 30784 4068 30796
rect 4023 30756 4068 30784
rect 4062 30744 4068 30756
rect 4120 30744 4126 30796
rect 9861 30787 9919 30793
rect 9861 30753 9873 30787
rect 9907 30784 9919 30787
rect 10134 30784 10140 30796
rect 9907 30756 10140 30784
rect 9907 30753 9919 30756
rect 9861 30747 9919 30753
rect 10134 30744 10140 30756
rect 10192 30744 10198 30796
rect 10042 30648 10048 30660
rect 10003 30620 10048 30648
rect 10042 30608 10048 30620
rect 10100 30608 10106 30660
rect 4154 30540 4160 30592
rect 4212 30580 4218 30592
rect 4249 30583 4307 30589
rect 4249 30580 4261 30583
rect 4212 30552 4261 30580
rect 4212 30540 4218 30552
rect 4249 30549 4261 30552
rect 4295 30549 4307 30583
rect 4249 30543 4307 30549
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 4062 30376 4068 30388
rect 4023 30348 4068 30376
rect 4062 30336 4068 30348
rect 4120 30336 4126 30388
rect 9769 30311 9827 30317
rect 9769 30277 9781 30311
rect 9815 30308 9827 30311
rect 10870 30308 10876 30320
rect 9815 30280 10876 30308
rect 9815 30277 9827 30280
rect 9769 30271 9827 30277
rect 9876 30181 9904 30280
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 9861 30175 9919 30181
rect 9861 30141 9873 30175
rect 9907 30141 9919 30175
rect 9861 30135 9919 30141
rect 11149 30175 11207 30181
rect 11149 30141 11161 30175
rect 11195 30172 11207 30175
rect 11195 30144 11836 30172
rect 11195 30141 11207 30144
rect 11149 30135 11207 30141
rect 10042 30036 10048 30048
rect 10003 30008 10048 30036
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 10134 29996 10140 30048
rect 10192 30036 10198 30048
rect 10505 30039 10563 30045
rect 10505 30036 10517 30039
rect 10192 30008 10517 30036
rect 10192 29996 10198 30008
rect 10505 30005 10517 30008
rect 10551 30036 10563 30039
rect 10962 30036 10968 30048
rect 10551 30008 10968 30036
rect 10551 30005 10563 30008
rect 10505 29999 10563 30005
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 11330 30036 11336 30048
rect 11291 30008 11336 30036
rect 11330 29996 11336 30008
rect 11388 29996 11394 30048
rect 11808 30045 11836 30144
rect 11793 30039 11851 30045
rect 11793 30005 11805 30039
rect 11839 30036 11851 30039
rect 11974 30036 11980 30048
rect 11839 30008 11980 30036
rect 11839 30005 11851 30008
rect 11793 29999 11851 30005
rect 11974 29996 11980 30008
rect 12032 29996 12038 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 11146 29696 11152 29708
rect 11107 29668 11152 29696
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 11330 29492 11336 29504
rect 11291 29464 11336 29492
rect 11330 29452 11336 29464
rect 11388 29452 11394 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 11146 29288 11152 29300
rect 11107 29260 11152 29288
rect 11146 29248 11152 29260
rect 11204 29248 11210 29300
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 10505 28747 10563 28753
rect 10505 28713 10517 28747
rect 10551 28744 10563 28747
rect 10778 28744 10784 28756
rect 10551 28716 10784 28744
rect 10551 28713 10563 28716
rect 10505 28707 10563 28713
rect 10778 28704 10784 28716
rect 10836 28704 10842 28756
rect 10321 28611 10379 28617
rect 10321 28577 10333 28611
rect 10367 28608 10379 28611
rect 10870 28608 10876 28620
rect 10367 28580 10876 28608
rect 10367 28577 10379 28580
rect 10321 28571 10379 28577
rect 10870 28568 10876 28580
rect 10928 28568 10934 28620
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 10229 28203 10287 28209
rect 10229 28169 10241 28203
rect 10275 28200 10287 28203
rect 10686 28200 10692 28212
rect 10275 28172 10692 28200
rect 10275 28169 10287 28172
rect 10229 28163 10287 28169
rect 10336 28005 10364 28172
rect 10686 28160 10692 28172
rect 10744 28160 10750 28212
rect 10321 27999 10379 28005
rect 10321 27965 10333 27999
rect 10367 27965 10379 27999
rect 10321 27959 10379 27965
rect 6822 27860 6828 27872
rect 6783 27832 6828 27860
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 10502 27860 10508 27872
rect 10463 27832 10508 27860
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 10870 27860 10876 27872
rect 10831 27832 10876 27860
rect 10870 27820 10876 27832
rect 10928 27820 10934 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 6914 27548 6920 27600
rect 6972 27588 6978 27600
rect 6972 27560 7017 27588
rect 6972 27548 6978 27560
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 4430 27452 4436 27464
rect 4212 27424 4436 27452
rect 4212 27412 4218 27424
rect 4430 27412 4436 27424
rect 4488 27412 4494 27464
rect 6822 27412 6828 27464
rect 6880 27452 6886 27464
rect 7009 27455 7067 27461
rect 7009 27452 7021 27455
rect 6880 27424 7021 27452
rect 6880 27412 6886 27424
rect 7009 27421 7021 27424
rect 7055 27421 7067 27455
rect 7190 27452 7196 27464
rect 7151 27424 7196 27452
rect 7009 27415 7067 27421
rect 7190 27412 7196 27424
rect 7248 27412 7254 27464
rect 5258 27276 5264 27328
rect 5316 27316 5322 27328
rect 6549 27319 6607 27325
rect 6549 27316 6561 27319
rect 5316 27288 6561 27316
rect 5316 27276 5322 27288
rect 6549 27285 6561 27288
rect 6595 27285 6607 27319
rect 6549 27279 6607 27285
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1578 27112 1584 27124
rect 1539 27084 1584 27112
rect 1578 27072 1584 27084
rect 1636 27072 1642 27124
rect 5905 27115 5963 27121
rect 5905 27081 5917 27115
rect 5951 27112 5963 27115
rect 6914 27112 6920 27124
rect 5951 27084 6920 27112
rect 5951 27081 5963 27084
rect 5905 27075 5963 27081
rect 6914 27072 6920 27084
rect 6972 27072 6978 27124
rect 6273 27047 6331 27053
rect 6273 27013 6285 27047
rect 6319 27044 6331 27047
rect 6546 27044 6552 27056
rect 6319 27016 6552 27044
rect 6319 27013 6331 27016
rect 6273 27007 6331 27013
rect 6546 27004 6552 27016
rect 6604 27044 6610 27056
rect 6822 27044 6828 27056
rect 6604 27016 6828 27044
rect 6604 27004 6610 27016
rect 6822 27004 6828 27016
rect 6880 27004 6886 27056
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7248 26948 7389 26976
rect 7248 26936 7254 26948
rect 7377 26945 7389 26948
rect 7423 26976 7435 26979
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7423 26948 7849 26976
rect 7423 26945 7435 26948
rect 7377 26939 7435 26945
rect 7837 26945 7849 26948
rect 7883 26945 7895 26979
rect 7837 26939 7895 26945
rect 1397 26911 1455 26917
rect 1397 26877 1409 26911
rect 1443 26908 1455 26911
rect 6638 26908 6644 26920
rect 1443 26880 1992 26908
rect 6599 26880 6644 26908
rect 1443 26877 1455 26880
rect 1397 26871 1455 26877
rect 1964 26781 1992 26880
rect 6638 26868 6644 26880
rect 6696 26908 6702 26920
rect 7285 26911 7343 26917
rect 6696 26880 7144 26908
rect 6696 26868 6702 26880
rect 1949 26775 2007 26781
rect 1949 26741 1961 26775
rect 1995 26772 2007 26775
rect 2682 26772 2688 26784
rect 1995 26744 2688 26772
rect 1995 26741 2007 26744
rect 1949 26735 2007 26741
rect 2682 26732 2688 26744
rect 2740 26732 2746 26784
rect 6822 26772 6828 26784
rect 6783 26744 6828 26772
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7116 26772 7144 26880
rect 7285 26877 7297 26911
rect 7331 26908 7343 26911
rect 7650 26908 7656 26920
rect 7331 26880 7656 26908
rect 7331 26877 7343 26880
rect 7285 26871 7343 26877
rect 7650 26868 7656 26880
rect 7708 26868 7714 26920
rect 7193 26775 7251 26781
rect 7193 26772 7205 26775
rect 7116 26744 7205 26772
rect 7193 26741 7205 26744
rect 7239 26772 7251 26775
rect 7926 26772 7932 26784
rect 7239 26744 7932 26772
rect 7239 26741 7251 26744
rect 7193 26735 7251 26741
rect 7926 26732 7932 26744
rect 7984 26732 7990 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 5350 26568 5356 26580
rect 5263 26540 5356 26568
rect 5350 26528 5356 26540
rect 5408 26568 5414 26580
rect 6822 26568 6828 26580
rect 5408 26540 6828 26568
rect 5408 26528 5414 26540
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7650 26568 7656 26580
rect 6972 26540 7656 26568
rect 6972 26528 6978 26540
rect 7650 26528 7656 26540
rect 7708 26528 7714 26580
rect 5258 26500 5264 26512
rect 5219 26472 5264 26500
rect 5258 26460 5264 26472
rect 5316 26500 5322 26512
rect 5626 26500 5632 26512
rect 5316 26472 5632 26500
rect 5316 26460 5322 26472
rect 5626 26460 5632 26472
rect 5684 26460 5690 26512
rect 5445 26367 5503 26373
rect 5445 26333 5457 26367
rect 5491 26333 5503 26367
rect 5445 26327 5503 26333
rect 4893 26299 4951 26305
rect 4893 26296 4905 26299
rect 4080 26268 4905 26296
rect 3326 26188 3332 26240
rect 3384 26228 3390 26240
rect 4080 26228 4108 26268
rect 4893 26265 4905 26268
rect 4939 26265 4951 26299
rect 4893 26259 4951 26265
rect 4982 26256 4988 26308
rect 5040 26296 5046 26308
rect 5460 26296 5488 26327
rect 7190 26296 7196 26308
rect 5040 26268 5488 26296
rect 7151 26268 7196 26296
rect 5040 26256 5046 26268
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 3384 26200 4108 26228
rect 3384 26188 3390 26200
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4982 26024 4988 26036
rect 4943 25996 4988 26024
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 5350 26024 5356 26036
rect 5311 25996 5356 26024
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 5626 26024 5632 26036
rect 5587 25996 5632 26024
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 3237 25483 3295 25489
rect 3237 25449 3249 25483
rect 3283 25480 3295 25483
rect 3326 25480 3332 25492
rect 3283 25452 3332 25480
rect 3283 25449 3295 25452
rect 3237 25443 3295 25449
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 12250 25480 12256 25492
rect 12211 25452 12256 25480
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 12066 25344 12072 25356
rect 12027 25316 12072 25344
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 2958 24760 2964 24812
rect 3016 24800 3022 24812
rect 3697 24803 3755 24809
rect 3697 24800 3709 24803
rect 3016 24772 3709 24800
rect 3016 24760 3022 24772
rect 3697 24769 3709 24772
rect 3743 24769 3755 24803
rect 3697 24763 3755 24769
rect 3510 24692 3516 24744
rect 3568 24732 3574 24744
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 3568 24704 3617 24732
rect 3568 24692 3574 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 2774 24624 2780 24676
rect 2832 24664 2838 24676
rect 2832 24636 3188 24664
rect 2832 24624 2838 24636
rect 2958 24596 2964 24608
rect 2919 24568 2964 24596
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 3160 24605 3188 24636
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24565 3203 24599
rect 3145 24559 3203 24565
rect 3326 24556 3332 24608
rect 3384 24596 3390 24608
rect 3513 24599 3571 24605
rect 3513 24596 3525 24599
rect 3384 24568 3525 24596
rect 3384 24556 3390 24568
rect 3513 24565 3525 24568
rect 3559 24565 3571 24599
rect 12066 24596 12072 24608
rect 12027 24568 12072 24596
rect 3513 24559 3571 24565
rect 12066 24556 12072 24568
rect 12124 24556 12130 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 3510 24052 3516 24064
rect 3283 24024 3516 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2406 22040 2412 22092
rect 2464 22080 2470 22092
rect 2590 22080 2596 22092
rect 2464 22052 2596 22080
rect 2464 22040 2470 22052
rect 2590 22040 2596 22052
rect 2648 22040 2654 22092
rect 12618 22040 12624 22092
rect 12676 22040 12682 22092
rect 12636 22012 12664 22040
rect 12802 22012 12808 22024
rect 12636 21984 12808 22012
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 4525 21879 4583 21885
rect 4525 21845 4537 21879
rect 4571 21876 4583 21879
rect 4798 21876 4804 21888
rect 4571 21848 4804 21876
rect 4571 21845 4583 21848
rect 4525 21839 4583 21845
rect 4798 21836 4804 21848
rect 4856 21836 4862 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 4433 21675 4491 21681
rect 4433 21672 4445 21675
rect 3568 21644 4445 21672
rect 3568 21632 3574 21644
rect 4433 21641 4445 21644
rect 4479 21641 4491 21675
rect 4433 21635 4491 21641
rect 4982 21536 4988 21548
rect 4895 21508 4988 21536
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 4341 21403 4399 21409
rect 4341 21369 4353 21403
rect 4387 21400 4399 21403
rect 5000 21400 5028 21496
rect 5350 21400 5356 21412
rect 4387 21372 5356 21400
rect 4387 21369 4399 21372
rect 4341 21363 4399 21369
rect 5350 21360 5356 21372
rect 5408 21360 5414 21412
rect 4798 21332 4804 21344
rect 4759 21304 4804 21332
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 4890 21292 4896 21344
rect 4948 21332 4954 21344
rect 4948 21304 4993 21332
rect 4948 21292 4954 21304
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 4798 21088 4804 21140
rect 4856 21128 4862 21140
rect 5905 21131 5963 21137
rect 5905 21128 5917 21131
rect 4856 21100 5917 21128
rect 4856 21088 4862 21100
rect 5905 21097 5917 21100
rect 5951 21097 5963 21131
rect 5905 21091 5963 21097
rect 7374 21088 7380 21140
rect 7432 21128 7438 21140
rect 7742 21128 7748 21140
rect 7432 21100 7748 21128
rect 7432 21088 7438 21100
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 5902 20952 5908 21004
rect 5960 20992 5966 21004
rect 6086 20992 6092 21004
rect 5960 20964 6092 20992
rect 5960 20952 5966 20964
rect 6086 20952 6092 20964
rect 6144 20992 6150 21004
rect 6273 20995 6331 21001
rect 6273 20992 6285 20995
rect 6144 20964 6285 20992
rect 6144 20952 6150 20964
rect 6273 20961 6285 20964
rect 6319 20961 6331 20995
rect 6273 20955 6331 20961
rect 6365 20995 6423 21001
rect 6365 20961 6377 20995
rect 6411 20992 6423 20995
rect 6730 20992 6736 21004
rect 6411 20964 6736 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 6454 20924 6460 20936
rect 6415 20896 6460 20924
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 4525 20791 4583 20797
rect 4525 20757 4537 20791
rect 4571 20788 4583 20791
rect 4890 20788 4896 20800
rect 4571 20760 4896 20788
rect 4571 20757 4583 20760
rect 4525 20751 4583 20757
rect 4890 20748 4896 20760
rect 4948 20788 4954 20800
rect 5626 20788 5632 20800
rect 4948 20760 5632 20788
rect 4948 20748 4954 20760
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 6144 20556 6377 20584
rect 6144 20544 6150 20556
rect 6365 20553 6377 20556
rect 6411 20584 6423 20587
rect 6454 20584 6460 20596
rect 6411 20556 6460 20584
rect 6411 20553 6423 20556
rect 6365 20547 6423 20553
rect 6454 20544 6460 20556
rect 6512 20584 6518 20596
rect 7190 20584 7196 20596
rect 6512 20556 7196 20584
rect 6512 20544 6518 20556
rect 7190 20544 7196 20556
rect 7248 20584 7254 20596
rect 9585 20587 9643 20593
rect 9585 20584 9597 20587
rect 7248 20556 9597 20584
rect 7248 20544 7254 20556
rect 9585 20553 9597 20556
rect 9631 20553 9643 20587
rect 9585 20547 9643 20553
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 8128 20352 8217 20380
rect 5629 20315 5687 20321
rect 5629 20281 5641 20315
rect 5675 20312 5687 20315
rect 6730 20312 6736 20324
rect 5675 20284 6736 20312
rect 5675 20281 5687 20284
rect 5629 20275 5687 20281
rect 6730 20272 6736 20284
rect 6788 20272 6794 20324
rect 8128 20256 8156 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 8205 20343 8263 20349
rect 8478 20321 8484 20324
rect 8472 20312 8484 20321
rect 8439 20284 8484 20312
rect 8472 20275 8484 20284
rect 8478 20272 8484 20275
rect 8536 20272 8542 20324
rect 5902 20244 5908 20256
rect 5863 20216 5908 20244
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 8110 20244 8116 20256
rect 8071 20216 8116 20244
rect 8110 20204 8116 20216
rect 8168 20204 8174 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 6788 20012 7205 20040
rect 6788 20000 6794 20012
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 5810 19932 5816 19984
rect 5868 19972 5874 19984
rect 6086 19972 6092 19984
rect 5868 19944 6092 19972
rect 5868 19932 5874 19944
rect 6086 19932 6092 19944
rect 6144 19932 6150 19984
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 5994 19904 6000 19916
rect 5583 19876 6000 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 5994 19864 6000 19876
rect 6052 19864 6058 19916
rect 6104 19904 6132 19932
rect 6104 19876 6224 19904
rect 6086 19836 6092 19848
rect 6047 19808 6092 19836
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6196 19845 6224 19876
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7558 19904 7564 19916
rect 7340 19876 7564 19904
rect 7340 19864 7346 19876
rect 7558 19864 7564 19876
rect 7616 19864 7622 19916
rect 7653 19907 7711 19913
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 7742 19904 7748 19916
rect 7699 19876 7748 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 9769 19907 9827 19913
rect 9769 19873 9781 19907
rect 9815 19904 9827 19907
rect 9858 19904 9864 19916
rect 9815 19876 9864 19904
rect 9815 19873 9827 19876
rect 9769 19867 9827 19873
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 10042 19913 10048 19916
rect 10036 19867 10048 19913
rect 10100 19904 10106 19916
rect 10100 19876 10136 19904
rect 10042 19864 10048 19867
rect 10100 19864 10106 19876
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 7834 19836 7840 19848
rect 7747 19808 7840 19836
rect 6181 19799 6239 19805
rect 7834 19796 7840 19808
rect 7892 19836 7898 19848
rect 7892 19808 8340 19836
rect 7892 19796 7898 19808
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7098 19700 7104 19712
rect 6963 19672 7104 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 8312 19709 8340 19808
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 8478 19700 8484 19712
rect 8343 19672 8484 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 8478 19660 8484 19672
rect 8536 19700 8542 19712
rect 11149 19703 11207 19709
rect 11149 19700 11161 19703
rect 8536 19672 11161 19700
rect 8536 19660 8542 19672
rect 11149 19669 11161 19672
rect 11195 19669 11207 19703
rect 11149 19663 11207 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6052 19468 6837 19496
rect 6052 19456 6058 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10137 19499 10195 19505
rect 10137 19496 10149 19499
rect 10100 19468 10149 19496
rect 10100 19456 10106 19468
rect 10137 19465 10149 19468
rect 10183 19465 10195 19499
rect 10137 19459 10195 19465
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7834 19360 7840 19372
rect 7515 19332 7840 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 2406 19252 2412 19304
rect 2464 19292 2470 19304
rect 2682 19292 2688 19304
rect 2464 19264 2688 19292
rect 2464 19252 2470 19264
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3878 19292 3884 19304
rect 3200 19264 3884 19292
rect 3200 19252 3206 19264
rect 3878 19252 3884 19264
rect 3936 19292 3942 19304
rect 3973 19295 4031 19301
rect 3973 19292 3985 19295
rect 3936 19264 3985 19292
rect 3936 19252 3942 19264
rect 3973 19261 3985 19264
rect 4019 19261 4031 19295
rect 4240 19295 4298 19301
rect 4240 19292 4252 19295
rect 3973 19255 4031 19261
rect 4172 19264 4252 19292
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 4172 19224 4200 19264
rect 4240 19261 4252 19264
rect 4286 19292 4298 19295
rect 5810 19292 5816 19304
rect 4286 19264 5816 19292
rect 4286 19261 4298 19264
rect 4240 19255 4298 19261
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6273 19295 6331 19301
rect 6273 19292 6285 19295
rect 6052 19264 6285 19292
rect 6052 19252 6058 19264
rect 6273 19261 6285 19264
rect 6319 19292 6331 19295
rect 7484 19292 7512 19323
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 6319 19264 7512 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 3559 19196 4200 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 6641 19227 6699 19233
rect 6641 19224 6653 19227
rect 5684 19196 6653 19224
rect 5684 19184 5690 19196
rect 6641 19193 6653 19196
rect 6687 19224 6699 19227
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 6687 19196 7297 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 7285 19193 7297 19196
rect 7331 19224 7343 19227
rect 8754 19224 8760 19236
rect 7331 19196 8760 19224
rect 7331 19193 7343 19196
rect 7285 19187 7343 19193
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 7098 19116 7104 19168
rect 7156 19156 7162 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 7156 19128 7205 19156
rect 7156 19116 7162 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7800 19128 7849 19156
rect 7800 19116 7806 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 9858 19156 9864 19168
rect 9819 19128 9864 19156
rect 7837 19119 7895 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 5810 18952 5816 18964
rect 5767 18924 5816 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 6086 18952 6092 18964
rect 6047 18924 6092 18952
rect 6086 18912 6092 18924
rect 6144 18952 6150 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 6144 18924 6285 18952
rect 6144 18912 6150 18924
rect 6273 18921 6285 18924
rect 6319 18921 6331 18955
rect 6273 18915 6331 18921
rect 7745 18955 7803 18961
rect 7745 18921 7757 18955
rect 7791 18952 7803 18955
rect 7834 18952 7840 18964
rect 7791 18924 7840 18952
rect 7791 18921 7803 18924
rect 7745 18915 7803 18921
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 6604 18788 6653 18816
rect 6604 18776 6610 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 6730 18748 6736 18760
rect 6691 18720 6736 18748
rect 6730 18708 6736 18720
rect 6788 18708 6794 18760
rect 6917 18751 6975 18757
rect 6917 18717 6929 18751
rect 6963 18748 6975 18751
rect 7760 18748 7788 18915
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 6963 18720 7788 18748
rect 6963 18717 6975 18720
rect 6917 18711 6975 18717
rect 7282 18612 7288 18624
rect 7243 18584 7288 18612
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 4525 18411 4583 18417
rect 4525 18408 4537 18411
rect 3568 18380 4537 18408
rect 3568 18368 3574 18380
rect 4525 18377 4537 18380
rect 4571 18377 4583 18411
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 4525 18371 4583 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18272 3111 18275
rect 3142 18272 3148 18284
rect 3099 18244 3148 18272
rect 3099 18241 3111 18244
rect 3053 18235 3111 18241
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 3234 18096 3240 18148
rect 3292 18136 3298 18148
rect 3390 18139 3448 18145
rect 3390 18136 3402 18139
rect 3292 18108 3402 18136
rect 3292 18096 3298 18108
rect 3390 18105 3402 18108
rect 3436 18136 3448 18139
rect 5350 18136 5356 18148
rect 3436 18108 5356 18136
rect 3436 18105 3448 18108
rect 3390 18099 3448 18105
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 6086 18096 6092 18148
rect 6144 18136 6150 18148
rect 6546 18136 6552 18148
rect 6144 18108 6552 18136
rect 6144 18096 6150 18108
rect 6546 18096 6552 18108
rect 6604 18136 6610 18148
rect 7009 18139 7067 18145
rect 7009 18136 7021 18139
rect 6604 18108 7021 18136
rect 6604 18096 6610 18108
rect 7009 18105 7021 18108
rect 7055 18136 7067 18139
rect 8386 18136 8392 18148
rect 7055 18108 8392 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 6365 18071 6423 18077
rect 6365 18037 6377 18071
rect 6411 18068 6423 18071
rect 6730 18068 6736 18080
rect 6411 18040 6736 18068
rect 6411 18037 6423 18040
rect 6365 18031 6423 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 3234 17864 3240 17876
rect 3195 17836 3240 17864
rect 3234 17824 3240 17836
rect 3292 17824 3298 17876
rect 6086 17824 6092 17876
rect 6144 17864 6150 17876
rect 6914 17864 6920 17876
rect 6144 17836 6920 17864
rect 6144 17824 6150 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 5810 17212 5816 17264
rect 5868 17252 5874 17264
rect 6178 17252 6184 17264
rect 5868 17224 6184 17252
rect 5868 17212 5874 17224
rect 6178 17212 6184 17224
rect 6236 17212 6242 17264
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 10134 14260 10140 14272
rect 9999 14232 10140 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14056 9922 14068
rect 10226 14056 10232 14068
rect 9916 14028 10232 14056
rect 9916 14016 9922 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 9876 13929 9904 14016
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10134 13861 10140 13864
rect 10128 13852 10140 13861
rect 10095 13824 10140 13852
rect 10128 13815 10140 13824
rect 10134 13812 10140 13815
rect 10192 13812 10198 13864
rect 10042 13676 10048 13728
rect 10100 13716 10106 13728
rect 11241 13719 11299 13725
rect 11241 13716 11253 13719
rect 10100 13688 11253 13716
rect 10100 13676 10106 13688
rect 11241 13685 11253 13688
rect 11287 13685 11299 13719
rect 11241 13679 11299 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 9950 13512 9956 13524
rect 9911 13484 9956 13512
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 10321 13379 10379 13385
rect 10321 13376 10333 13379
rect 9916 13348 10333 13376
rect 9916 13336 9922 13348
rect 10321 13345 10333 13348
rect 10367 13345 10379 13379
rect 10321 13339 10379 13345
rect 10410 13308 10416 13320
rect 10371 13280 10416 13308
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10520 13240 10548 13271
rect 10100 13212 10548 13240
rect 10100 13200 10106 13212
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 2498 12928 2504 12980
rect 2556 12968 2562 12980
rect 7374 12968 7380 12980
rect 2556 12940 7380 12968
rect 2556 12928 2562 12940
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10689 12767 10747 12773
rect 10689 12764 10701 12767
rect 9916 12736 10701 12764
rect 9916 12724 9922 12736
rect 10689 12733 10701 12736
rect 10735 12733 10747 12767
rect 10689 12727 10747 12733
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9640 12600 10333 12628
rect 9640 12588 9646 12600
rect 10321 12597 10333 12600
rect 10367 12628 10379 12631
rect 10410 12628 10416 12640
rect 10367 12600 10416 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 7742 12084 7748 12096
rect 7703 12056 7748 12084
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 9309 12087 9367 12093
rect 9309 12084 9321 12087
rect 8904 12056 9321 12084
rect 8904 12044 8910 12056
rect 9309 12053 9321 12056
rect 9355 12053 9367 12087
rect 9309 12047 9367 12053
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 8846 11880 8852 11892
rect 7791 11852 8852 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 9582 11880 9588 11892
rect 9355 11852 9588 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8168 11716 8309 11744
rect 8168 11704 8174 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9263 11716 9965 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9953 11713 9965 11716
rect 9999 11744 10011 11747
rect 10134 11744 10140 11756
rect 9999 11716 10140 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 8846 11636 8852 11688
rect 8904 11676 8910 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 8904 11648 9689 11676
rect 8904 11636 8910 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10962 11676 10968 11688
rect 9824 11648 10968 11676
rect 9824 11636 9830 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7742 11608 7748 11620
rect 6972 11580 7748 11608
rect 6972 11568 6978 11580
rect 7742 11568 7748 11580
rect 7800 11608 7806 11620
rect 8205 11611 8263 11617
rect 8205 11608 8217 11611
rect 7800 11580 8217 11608
rect 7800 11568 7806 11580
rect 8205 11577 8217 11580
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 8018 11540 8024 11552
rect 7699 11512 8024 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8018 11500 8024 11512
rect 8076 11540 8082 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 8076 11512 8125 11540
rect 8076 11500 8082 11512
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 8113 11503 8171 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7006 11132 7012 11144
rect 6967 11104 7012 11132
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7156 11104 7757 11132
rect 7156 11092 7162 11104
rect 7745 11101 7757 11104
rect 7791 11132 7803 11135
rect 8110 11132 8116 11144
rect 7791 11104 8116 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 6549 11067 6607 11073
rect 6549 11033 6561 11067
rect 6595 11064 6607 11067
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 6595 11036 9321 11064
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 9309 11033 9321 11036
rect 9355 11064 9367 11067
rect 9766 11064 9772 11076
rect 9355 11036 9772 11064
rect 9355 11033 9367 11036
rect 9309 11027 9367 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 6822 10792 6828 10804
rect 6783 10764 6828 10792
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 5905 10727 5963 10733
rect 5905 10693 5917 10727
rect 5951 10724 5963 10727
rect 7098 10724 7104 10736
rect 5951 10696 7104 10724
rect 5951 10693 5963 10696
rect 5905 10687 5963 10693
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6236 10628 7389 10656
rect 6236 10616 6242 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7064 10560 7849 10588
rect 7064 10548 7070 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 6972 10492 8217 10520
rect 6972 10480 6978 10492
rect 8205 10489 8217 10492
rect 8251 10489 8263 10523
rect 8205 10483 8263 10489
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 6730 10452 6736 10464
rect 6687 10424 6736 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 7156 10424 7205 10452
rect 7156 10412 7162 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7193 10415 7251 10421
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 7340 10424 7385 10452
rect 7340 10412 7346 10424
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 7432 10220 7757 10248
rect 7432 10208 7438 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 7745 10211 7803 10217
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 6052 10084 6101 10112
rect 6052 10072 6058 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 7650 10112 7656 10124
rect 7563 10084 7656 10112
rect 6089 10075 6147 10081
rect 7650 10072 7656 10084
rect 7708 10112 7714 10124
rect 8570 10112 8576 10124
rect 7708 10084 8576 10112
rect 7708 10072 7714 10084
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 6178 10044 6184 10056
rect 5684 10016 6184 10044
rect 5684 10004 5690 10016
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6362 10004 6368 10016
rect 6420 10044 6426 10056
rect 7837 10047 7895 10053
rect 6420 10016 7696 10044
rect 6420 10004 6426 10016
rect 5721 9979 5779 9985
rect 5721 9945 5733 9979
rect 5767 9976 5779 9979
rect 7006 9976 7012 9988
rect 5767 9948 7012 9976
rect 5767 9945 5779 9948
rect 5721 9939 5779 9945
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7668 9976 7696 10016
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 7852 9976 7880 10007
rect 8018 9976 8024 9988
rect 7668 9948 8024 9976
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7098 9908 7104 9920
rect 6963 9880 7104 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7098 9868 7104 9880
rect 7156 9908 7162 9920
rect 7282 9908 7288 9920
rect 7156 9880 7288 9908
rect 7156 9868 7162 9880
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6089 9707 6147 9713
rect 6089 9704 6101 9707
rect 6052 9676 6101 9704
rect 6052 9664 6058 9676
rect 6089 9673 6101 9676
rect 6135 9673 6147 9707
rect 7650 9704 7656 9716
rect 7611 9676 7656 9704
rect 6089 9667 6147 9673
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 8018 9704 8024 9716
rect 7979 9676 8024 9704
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 4798 9596 4804 9648
rect 4856 9636 4862 9648
rect 5166 9636 5172 9648
rect 4856 9608 5172 9636
rect 4856 9596 4862 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11514 9636 11520 9648
rect 11296 9608 11520 9636
rect 11296 9596 11302 9608
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 6362 9432 6368 9444
rect 5592 9404 6368 9432
rect 5592 9392 5598 9404
rect 6362 9392 6368 9404
rect 6420 9432 6426 9444
rect 6457 9435 6515 9441
rect 6457 9432 6469 9435
rect 6420 9404 6469 9432
rect 6420 9392 6426 9404
rect 6457 9401 6469 9404
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 5994 9364 6000 9376
rect 5859 9336 6000 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 5994 9324 6000 9336
rect 6052 9364 6058 9376
rect 6178 9364 6184 9376
rect 6052 9336 6184 9364
rect 6052 9324 6058 9336
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 7374 9364 7380 9376
rect 7335 9336 7380 9364
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13722 8276 13728 8288
rect 12768 8248 13728 8276
rect 12768 8236 12774 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 13354 8072 13360 8084
rect 12584 8044 13360 8072
rect 12584 8032 12590 8044
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14918 7732 14924 7744
rect 14056 7704 14924 7732
rect 14056 7692 14062 7704
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 15746 7528 15752 7540
rect 13964 7500 15752 7528
rect 13964 7488 13970 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 4212 6820 4333 6848
rect 4212 6808 4218 6820
rect 4321 6817 4333 6820
rect 4367 6817 4379 6851
rect 4321 6811 4379 6817
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4080 6644 4108 6743
rect 4246 6644 4252 6656
rect 4080 6616 4252 6644
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 5445 6647 5503 6653
rect 5445 6613 5457 6647
rect 5491 6644 5503 6647
rect 5534 6644 5540 6656
rect 5491 6616 5540 6644
rect 5491 6613 5503 6616
rect 5445 6607 5503 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10318 6644 10324 6656
rect 9999 6616 10324 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 9858 6440 9864 6452
rect 9819 6412 9864 6440
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 9769 6375 9827 6381
rect 9769 6341 9781 6375
rect 9815 6372 9827 6375
rect 10134 6372 10140 6384
rect 9815 6344 10140 6372
rect 9815 6341 9827 6344
rect 9769 6335 9827 6341
rect 10134 6332 10140 6344
rect 10192 6372 10198 6384
rect 10192 6344 10548 6372
rect 10192 6332 10198 6344
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10520 6313 10548 6344
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10594 6304 10600 6316
rect 10551 6276 10600 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 10134 6168 10140 6180
rect 9447 6140 10140 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10134 6128 10140 6140
rect 10192 6168 10198 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 10192 6140 10241 6168
rect 10192 6128 10198 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 4246 6060 4252 6112
rect 4304 6100 4310 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4304 6072 4537 6100
rect 4304 6060 4310 6072
rect 4525 6069 4537 6072
rect 4571 6100 4583 6103
rect 5626 6100 5632 6112
rect 4571 6072 5632 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 8352 5868 9229 5896
rect 8352 5856 8358 5868
rect 9217 5865 9229 5868
rect 9263 5896 9275 5899
rect 9306 5896 9312 5908
rect 9263 5868 9312 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9861 5899 9919 5905
rect 9861 5865 9873 5899
rect 9907 5896 9919 5899
rect 10318 5896 10324 5908
rect 9907 5868 10324 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10226 5828 10232 5840
rect 10187 5800 10232 5828
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 9640 5732 10333 5760
rect 9640 5720 9646 5732
rect 10321 5729 10333 5732
rect 10367 5760 10379 5763
rect 11422 5760 11428 5772
rect 10367 5732 11428 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 9364 5664 10425 5692
rect 9364 5652 9370 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8168 5324 9137 5352
rect 8168 5312 8174 5324
rect 9125 5321 9137 5324
rect 9171 5352 9183 5355
rect 9582 5352 9588 5364
rect 9171 5324 9588 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9232 5012 9260 5111
rect 9306 5108 9312 5160
rect 9364 5148 9370 5160
rect 9473 5151 9531 5157
rect 9473 5148 9485 5151
rect 9364 5120 9485 5148
rect 9364 5108 9370 5120
rect 9473 5117 9485 5120
rect 9519 5117 9531 5151
rect 9473 5111 9531 5117
rect 9490 5012 9496 5024
rect 9232 4984 9496 5012
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10744 4984 11161 5012
rect 10744 4972 10750 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8202 4808 8208 4820
rect 7791 4780 8208 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 9490 4808 9496 4820
rect 9355 4780 9496 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6632 4743 6690 4749
rect 6632 4740 6644 4743
rect 5592 4712 6644 4740
rect 5592 4700 5598 4712
rect 6632 4709 6644 4712
rect 6678 4740 6690 4743
rect 6822 4740 6828 4752
rect 6678 4712 6828 4740
rect 6678 4709 6690 4712
rect 6632 4703 6690 4709
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 5684 4644 6377 4672
rect 5684 4632 5690 4644
rect 6365 4641 6377 4644
rect 6411 4672 6423 4675
rect 6454 4672 6460 4684
rect 6411 4644 6460 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 6454 4632 6460 4644
rect 6512 4672 6518 4684
rect 9324 4672 9352 4771
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 9953 4743 10011 4749
rect 9953 4709 9965 4743
rect 9999 4740 10011 4743
rect 10226 4740 10232 4752
rect 9999 4712 10232 4740
rect 9999 4709 10011 4712
rect 9953 4703 10011 4709
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 10502 4672 10508 4684
rect 6512 4644 9352 4672
rect 10463 4644 10508 4672
rect 6512 4632 6518 4644
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 10686 4604 10692 4616
rect 9364 4576 10692 4604
rect 9364 4564 9370 4576
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 6454 4264 6460 4276
rect 6415 4236 6460 4264
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9364 4236 9781 4264
rect 9364 4224 9370 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 10502 4264 10508 4276
rect 9769 4227 9827 4233
rect 10336 4236 10508 4264
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 4062 4128 4068 4140
rect 3016 4100 4068 4128
rect 3016 4088 3022 4100
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5442 4128 5448 4140
rect 5040 4100 5448 4128
rect 5040 4088 5046 4100
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 10336 4137 10364 4236
rect 10502 4224 10508 4236
rect 10560 4264 10566 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10560 4236 10793 4264
rect 10560 4224 10566 4236
rect 10781 4233 10793 4236
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6880 4100 7021 4128
rect 6880 4088 6886 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10229 4063 10287 4069
rect 10229 4029 10241 4063
rect 10275 4060 10287 4063
rect 10594 4060 10600 4072
rect 10275 4032 10600 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12986 3720 12992 3732
rect 12492 3692 12992 3720
rect 12492 3680 12498 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 4028 3556 4077 3584
rect 4028 3544 4034 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 6086 3584 6092 3596
rect 5215 3556 6092 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6638 3584 6644 3596
rect 6319 3556 6644 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 4246 3448 4252 3460
rect 4207 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 4580 3352 5365 3380
rect 4580 3340 4586 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 6457 3383 6515 3389
rect 6457 3349 6469 3383
rect 6503 3380 6515 3383
rect 6914 3380 6920 3392
rect 6503 3352 6920 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 3384 3148 3433 3176
rect 3384 3136 3390 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 3881 3179 3939 3185
rect 3881 3145 3893 3179
rect 3927 3176 3939 3179
rect 3970 3176 3976 3188
rect 3927 3148 3976 3176
rect 3927 3145 3939 3148
rect 3881 3139 3939 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4154 3176 4160 3188
rect 4115 3148 4160 3176
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5074 3176 5080 3188
rect 5031 3148 5080 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6086 3176 6092 3188
rect 5767 3148 6092 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6638 3176 6644 3188
rect 6411 3148 6644 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7926 3176 7932 3188
rect 7887 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 2130 3068 2136 3120
rect 2188 3108 2194 3120
rect 5261 3111 5319 3117
rect 5261 3108 5273 3111
rect 2188 3080 5273 3108
rect 2188 3068 2194 3080
rect 5261 3077 5273 3080
rect 5307 3077 5319 3111
rect 5261 3071 5319 3077
rect 4614 3040 4620 3052
rect 3988 3012 4620 3040
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3326 2972 3332 2984
rect 2915 2944 3332 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3988 2981 4016 3012
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2941 4031 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 3973 2935 4031 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 7285 2975 7343 2981
rect 7285 2941 7297 2975
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2924 2808 3065 2836
rect 2924 2796 2930 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 7469 2839 7527 2845
rect 7469 2836 7481 2839
rect 6696 2808 7481 2836
rect 6696 2796 6702 2808
rect 7469 2805 7481 2808
rect 7515 2805 7527 2839
rect 7469 2799 7527 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 7282 2632 7288 2644
rect 5859 2604 7288 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2496 1458 2508
rect 1949 2499 2007 2505
rect 1949 2496 1961 2499
rect 1452 2468 1961 2496
rect 1452 2456 1458 2468
rect 1949 2465 1961 2468
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3436 2496 3464 2592
rect 2915 2468 3464 2496
rect 4065 2499 4123 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4706 2496 4712 2508
rect 4111 2468 4712 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5828 2496 5856 2595
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2632 7987 2635
rect 8110 2632 8116 2644
rect 7975 2604 8116 2632
rect 7975 2601 7987 2604
rect 7929 2595 7987 2601
rect 5215 2468 5856 2496
rect 7285 2499 7343 2505
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 7944 2496 7972 2595
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11790 2564 11796 2576
rect 11204 2536 11796 2564
rect 11204 2524 11210 2536
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 7331 2468 7972 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1762 2252 1768 2304
rect 1820 2292 1826 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 1820 2264 5365 2292
rect 1820 2252 1826 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 4798 552 4804 604
rect 4856 592 4862 604
rect 5350 592 5356 604
rect 4856 564 5356 592
rect 4856 552 4862 564
rect 5350 552 5356 564
rect 5408 552 5414 604
rect 11330 552 11336 604
rect 11388 592 11394 604
rect 11514 592 11520 604
rect 11388 564 11520 592
rect 11388 552 11394 564
rect 11514 552 11520 564
rect 11572 552 11578 604
<< via1 >>
rect 13820 37748 13872 37800
rect 14556 37748 14608 37800
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 204 34484 256 34536
rect 1308 34484 1360 34536
rect 1400 34484 1452 34536
rect 2780 34484 2832 34536
rect 2964 34484 3016 34536
rect 4068 34484 4120 34536
rect 4160 34484 4212 34536
rect 5540 34484 5592 34536
rect 7748 34484 7800 34536
rect 8208 34484 8260 34536
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 2780 32512 2832 32564
rect 4160 32512 4212 32564
rect 7472 32555 7524 32564
rect 7472 32521 7481 32555
rect 7481 32521 7515 32555
rect 7515 32521 7524 32555
rect 7472 32512 7524 32521
rect 9588 32555 9640 32564
rect 9588 32521 9597 32555
rect 9597 32521 9631 32555
rect 9631 32521 9640 32555
rect 9588 32512 9640 32521
rect 10692 32555 10744 32564
rect 10692 32521 10701 32555
rect 10701 32521 10735 32555
rect 10735 32521 10744 32555
rect 10692 32512 10744 32521
rect 13084 32555 13136 32564
rect 13084 32521 13093 32555
rect 13093 32521 13127 32555
rect 13127 32521 13136 32555
rect 13084 32512 13136 32521
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 3056 32308 3108 32317
rect 4436 32308 4488 32360
rect 9588 32308 9640 32360
rect 10692 32308 10744 32360
rect 13084 32308 13136 32360
rect 7472 32240 7524 32292
rect 7288 32172 7340 32224
rect 8852 32172 8904 32224
rect 9680 32172 9732 32224
rect 12624 32215 12676 32224
rect 12624 32181 12633 32215
rect 12633 32181 12667 32215
rect 12667 32181 12676 32215
rect 12624 32172 12676 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 1400 31968 1452 32020
rect 2872 31968 2924 32020
rect 4344 31968 4396 32020
rect 5540 32011 5592 32020
rect 5540 31977 5549 32011
rect 5549 31977 5583 32011
rect 5583 31977 5592 32011
rect 5540 31968 5592 31977
rect 6828 31968 6880 32020
rect 8024 32011 8076 32020
rect 8024 31977 8033 32011
rect 8033 31977 8067 32011
rect 8067 31977 8076 32011
rect 8024 31968 8076 31977
rect 9864 32011 9916 32020
rect 9864 31977 9873 32011
rect 9873 31977 9907 32011
rect 9907 31977 9916 32011
rect 9864 31968 9916 31977
rect 12532 32011 12584 32020
rect 12532 31977 12541 32011
rect 12541 31977 12575 32011
rect 12575 31977 12584 32011
rect 12532 31968 12584 31977
rect 1676 31875 1728 31884
rect 1676 31841 1685 31875
rect 1685 31841 1719 31875
rect 1719 31841 1728 31875
rect 1676 31832 1728 31841
rect 3240 31832 3292 31884
rect 5448 31832 5500 31884
rect 6460 31875 6512 31884
rect 6460 31841 6469 31875
rect 6469 31841 6503 31875
rect 6503 31841 6512 31875
rect 6460 31832 6512 31841
rect 7840 31875 7892 31884
rect 7840 31841 7849 31875
rect 7849 31841 7883 31875
rect 7883 31841 7892 31875
rect 7840 31832 7892 31841
rect 10508 31832 10560 31884
rect 13452 31875 13504 31884
rect 7288 31764 7340 31816
rect 7748 31764 7800 31816
rect 4344 31696 4396 31748
rect 13452 31841 13461 31875
rect 13461 31841 13495 31875
rect 13495 31841 13504 31875
rect 13452 31832 13504 31841
rect 12992 31696 13044 31748
rect 13636 31671 13688 31680
rect 13636 31637 13645 31671
rect 13645 31637 13679 31671
rect 13679 31637 13688 31671
rect 13636 31628 13688 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 2872 31467 2924 31476
rect 2872 31433 2881 31467
rect 2881 31433 2915 31467
rect 2915 31433 2924 31467
rect 2872 31424 2924 31433
rect 4528 31424 4580 31476
rect 6460 31467 6512 31476
rect 6460 31433 6469 31467
rect 6469 31433 6503 31467
rect 6503 31433 6512 31467
rect 6460 31424 6512 31433
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 13452 31467 13504 31476
rect 13452 31433 13461 31467
rect 13461 31433 13495 31467
rect 13495 31433 13504 31467
rect 13452 31424 13504 31433
rect 2136 31356 2188 31408
rect 9680 31399 9732 31408
rect 9680 31365 9689 31399
rect 9689 31365 9723 31399
rect 9723 31365 9732 31399
rect 9680 31356 9732 31365
rect 1676 31127 1728 31136
rect 1676 31093 1685 31127
rect 1685 31093 1719 31127
rect 1719 31093 1728 31127
rect 1676 31084 1728 31093
rect 2504 31127 2556 31136
rect 2504 31093 2513 31127
rect 2513 31093 2547 31127
rect 2547 31093 2556 31127
rect 2504 31084 2556 31093
rect 3240 31127 3292 31136
rect 3240 31093 3249 31127
rect 3249 31093 3283 31127
rect 3283 31093 3292 31127
rect 3240 31084 3292 31093
rect 3424 31084 3476 31136
rect 13912 31220 13964 31272
rect 4344 31127 4396 31136
rect 4344 31093 4353 31127
rect 4353 31093 4387 31127
rect 4387 31093 4396 31127
rect 4344 31084 4396 31093
rect 4712 31127 4764 31136
rect 4712 31093 4721 31127
rect 4721 31093 4755 31127
rect 4755 31093 4764 31127
rect 4712 31084 4764 31093
rect 5540 31127 5592 31136
rect 5540 31093 5549 31127
rect 5549 31093 5583 31127
rect 5583 31093 5592 31127
rect 5540 31084 5592 31093
rect 7380 31127 7432 31136
rect 7380 31093 7389 31127
rect 7389 31093 7423 31127
rect 7423 31093 7432 31127
rect 7380 31084 7432 31093
rect 7840 31127 7892 31136
rect 7840 31093 7849 31127
rect 7849 31093 7883 31127
rect 7883 31093 7892 31127
rect 7840 31084 7892 31093
rect 9956 31084 10008 31136
rect 10508 31127 10560 31136
rect 10508 31093 10517 31127
rect 10517 31093 10551 31127
rect 10551 31093 10560 31127
rect 10508 31084 10560 31093
rect 10968 31084 11020 31136
rect 12532 31084 12584 31136
rect 12992 31127 13044 31136
rect 12992 31093 13001 31127
rect 13001 31093 13035 31127
rect 13035 31093 13044 31127
rect 12992 31084 13044 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 7472 30880 7524 30932
rect 8116 30880 8168 30932
rect 4068 30787 4120 30796
rect 4068 30753 4077 30787
rect 4077 30753 4111 30787
rect 4111 30753 4120 30787
rect 4068 30744 4120 30753
rect 10140 30744 10192 30796
rect 10048 30651 10100 30660
rect 10048 30617 10057 30651
rect 10057 30617 10091 30651
rect 10091 30617 10100 30651
rect 10048 30608 10100 30617
rect 4160 30540 4212 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 4068 30379 4120 30388
rect 4068 30345 4077 30379
rect 4077 30345 4111 30379
rect 4111 30345 4120 30379
rect 4068 30336 4120 30345
rect 10876 30268 10928 30320
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 10140 29996 10192 30048
rect 10968 29996 11020 30048
rect 11336 30039 11388 30048
rect 11336 30005 11345 30039
rect 11345 30005 11379 30039
rect 11379 30005 11388 30039
rect 11336 29996 11388 30005
rect 11980 29996 12032 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 11152 29699 11204 29708
rect 11152 29665 11161 29699
rect 11161 29665 11195 29699
rect 11195 29665 11204 29699
rect 11152 29656 11204 29665
rect 11336 29495 11388 29504
rect 11336 29461 11345 29495
rect 11345 29461 11379 29495
rect 11379 29461 11388 29495
rect 11336 29452 11388 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 11152 29291 11204 29300
rect 11152 29257 11161 29291
rect 11161 29257 11195 29291
rect 11195 29257 11204 29291
rect 11152 29248 11204 29257
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 10784 28704 10836 28756
rect 10876 28568 10928 28620
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 10692 28160 10744 28212
rect 6828 27863 6880 27872
rect 6828 27829 6837 27863
rect 6837 27829 6871 27863
rect 6871 27829 6880 27863
rect 6828 27820 6880 27829
rect 10508 27863 10560 27872
rect 10508 27829 10517 27863
rect 10517 27829 10551 27863
rect 10551 27829 10560 27863
rect 10508 27820 10560 27829
rect 10876 27863 10928 27872
rect 10876 27829 10885 27863
rect 10885 27829 10919 27863
rect 10919 27829 10928 27863
rect 10876 27820 10928 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 6920 27591 6972 27600
rect 6920 27557 6929 27591
rect 6929 27557 6963 27591
rect 6963 27557 6972 27591
rect 6920 27548 6972 27557
rect 4160 27412 4212 27464
rect 4436 27412 4488 27464
rect 6828 27412 6880 27464
rect 7196 27455 7248 27464
rect 7196 27421 7205 27455
rect 7205 27421 7239 27455
rect 7239 27421 7248 27455
rect 7196 27412 7248 27421
rect 5264 27276 5316 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 1584 27115 1636 27124
rect 1584 27081 1593 27115
rect 1593 27081 1627 27115
rect 1627 27081 1636 27115
rect 1584 27072 1636 27081
rect 6920 27072 6972 27124
rect 6552 27004 6604 27056
rect 6828 27004 6880 27056
rect 7196 26936 7248 26988
rect 6644 26911 6696 26920
rect 6644 26877 6653 26911
rect 6653 26877 6687 26911
rect 6687 26877 6696 26911
rect 6644 26868 6696 26877
rect 2688 26732 2740 26784
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 7656 26868 7708 26920
rect 7932 26732 7984 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 5356 26571 5408 26580
rect 5356 26537 5365 26571
rect 5365 26537 5399 26571
rect 5399 26537 5408 26571
rect 5356 26528 5408 26537
rect 6828 26528 6880 26580
rect 6920 26571 6972 26580
rect 6920 26537 6929 26571
rect 6929 26537 6963 26571
rect 6963 26537 6972 26571
rect 6920 26528 6972 26537
rect 7656 26528 7708 26580
rect 5264 26503 5316 26512
rect 5264 26469 5273 26503
rect 5273 26469 5307 26503
rect 5307 26469 5316 26503
rect 5264 26460 5316 26469
rect 5632 26460 5684 26512
rect 3332 26188 3384 26240
rect 4988 26256 5040 26308
rect 7196 26299 7248 26308
rect 7196 26265 7205 26299
rect 7205 26265 7239 26299
rect 7239 26265 7248 26299
rect 7196 26256 7248 26265
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4988 26027 5040 26036
rect 4988 25993 4997 26027
rect 4997 25993 5031 26027
rect 5031 25993 5040 26027
rect 4988 25984 5040 25993
rect 5356 26027 5408 26036
rect 5356 25993 5365 26027
rect 5365 25993 5399 26027
rect 5399 25993 5408 26027
rect 5356 25984 5408 25993
rect 5632 26027 5684 26036
rect 5632 25993 5641 26027
rect 5641 25993 5675 26027
rect 5675 25993 5684 26027
rect 5632 25984 5684 25993
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 3332 25440 3384 25492
rect 12256 25483 12308 25492
rect 12256 25449 12265 25483
rect 12265 25449 12299 25483
rect 12299 25449 12308 25483
rect 12256 25440 12308 25449
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2964 24760 3016 24812
rect 3516 24692 3568 24744
rect 2780 24624 2832 24676
rect 2964 24599 3016 24608
rect 2964 24565 2973 24599
rect 2973 24565 3007 24599
rect 3007 24565 3016 24599
rect 2964 24556 3016 24565
rect 3332 24556 3384 24608
rect 12072 24599 12124 24608
rect 12072 24565 12081 24599
rect 12081 24565 12115 24599
rect 12115 24565 12124 24599
rect 12072 24556 12124 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 3516 24012 3568 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2412 22040 2464 22092
rect 2596 22040 2648 22092
rect 12624 22040 12676 22092
rect 12808 21972 12860 22024
rect 4804 21836 4856 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 3516 21632 3568 21684
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 5356 21360 5408 21412
rect 4804 21335 4856 21344
rect 4804 21301 4813 21335
rect 4813 21301 4847 21335
rect 4847 21301 4856 21335
rect 4804 21292 4856 21301
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 4804 21088 4856 21140
rect 7380 21088 7432 21140
rect 7748 21088 7800 21140
rect 5908 20952 5960 21004
rect 6092 20952 6144 21004
rect 6736 20952 6788 21004
rect 6460 20927 6512 20936
rect 6460 20893 6469 20927
rect 6469 20893 6503 20927
rect 6503 20893 6512 20927
rect 6460 20884 6512 20893
rect 4896 20748 4948 20800
rect 5632 20748 5684 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 6092 20544 6144 20596
rect 6460 20544 6512 20596
rect 7196 20544 7248 20596
rect 6736 20272 6788 20324
rect 8484 20315 8536 20324
rect 8484 20281 8518 20315
rect 8518 20281 8536 20315
rect 8484 20272 8536 20281
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 8116 20247 8168 20256
rect 8116 20213 8125 20247
rect 8125 20213 8159 20247
rect 8159 20213 8168 20247
rect 8116 20204 8168 20213
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 6736 20000 6788 20052
rect 5816 19932 5868 19984
rect 6092 19932 6144 19984
rect 6000 19907 6052 19916
rect 6000 19873 6009 19907
rect 6009 19873 6043 19907
rect 6043 19873 6052 19907
rect 6000 19864 6052 19873
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 7288 19864 7340 19916
rect 7564 19907 7616 19916
rect 7564 19873 7573 19907
rect 7573 19873 7607 19907
rect 7607 19873 7616 19907
rect 7564 19864 7616 19873
rect 7748 19864 7800 19916
rect 9864 19864 9916 19916
rect 10048 19907 10100 19916
rect 10048 19873 10082 19907
rect 10082 19873 10100 19907
rect 10048 19864 10100 19873
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 7104 19660 7156 19712
rect 8484 19660 8536 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 6000 19456 6052 19508
rect 10048 19456 10100 19508
rect 2412 19252 2464 19304
rect 2688 19252 2740 19304
rect 3148 19252 3200 19304
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 5816 19252 5868 19304
rect 6000 19252 6052 19304
rect 7840 19320 7892 19372
rect 5632 19184 5684 19236
rect 8760 19184 8812 19236
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 7104 19116 7156 19168
rect 7748 19116 7800 19168
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 9864 19116 9916 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 5816 18912 5868 18964
rect 6092 18955 6144 18964
rect 6092 18921 6101 18955
rect 6101 18921 6135 18955
rect 6135 18921 6144 18955
rect 6092 18912 6144 18921
rect 6552 18776 6604 18828
rect 6736 18751 6788 18760
rect 6736 18717 6745 18751
rect 6745 18717 6779 18751
rect 6779 18717 6788 18751
rect 6736 18708 6788 18717
rect 7840 18912 7892 18964
rect 7288 18615 7340 18624
rect 7288 18581 7297 18615
rect 7297 18581 7331 18615
rect 7331 18581 7340 18615
rect 7288 18572 7340 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 3516 18368 3568 18420
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 3240 18096 3292 18148
rect 5356 18096 5408 18148
rect 6092 18096 6144 18148
rect 6552 18096 6604 18148
rect 8392 18096 8444 18148
rect 6736 18028 6788 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3240 17867 3292 17876
rect 3240 17833 3249 17867
rect 3249 17833 3283 17867
rect 3283 17833 3292 17867
rect 3240 17824 3292 17833
rect 6092 17824 6144 17876
rect 6920 17824 6972 17876
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 5816 17212 5868 17264
rect 6184 17212 6236 17264
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 10140 14220 10192 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 9864 14016 9916 14068
rect 10232 14016 10284 14068
rect 10140 13855 10192 13864
rect 10140 13821 10174 13855
rect 10174 13821 10192 13855
rect 10140 13812 10192 13821
rect 10048 13676 10100 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 9956 13515 10008 13524
rect 9956 13481 9965 13515
rect 9965 13481 9999 13515
rect 9999 13481 10008 13515
rect 9956 13472 10008 13481
rect 9864 13336 9916 13388
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10048 13200 10100 13252
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 2504 12928 2556 12980
rect 7380 12928 7432 12980
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 9864 12724 9916 12776
rect 9588 12588 9640 12640
rect 10416 12588 10468 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 8852 12044 8904 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 8852 11840 8904 11892
rect 9588 11840 9640 11892
rect 8116 11704 8168 11756
rect 10140 11704 10192 11756
rect 8852 11636 8904 11688
rect 9772 11636 9824 11688
rect 10968 11636 11020 11688
rect 6920 11568 6972 11620
rect 7748 11568 7800 11620
rect 8024 11500 8076 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 8116 11092 8168 11144
rect 9772 11024 9824 11076
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 7104 10684 7156 10736
rect 6184 10616 6236 10668
rect 7012 10548 7064 10600
rect 6920 10480 6972 10532
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 6736 10412 6788 10464
rect 7104 10412 7156 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 6920 10208 6972 10260
rect 7380 10208 7432 10260
rect 6000 10072 6052 10124
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 8576 10072 8628 10124
rect 5632 10004 5684 10056
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 7012 9936 7064 9988
rect 8024 9936 8076 9988
rect 7104 9868 7156 9920
rect 7288 9868 7340 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 6000 9664 6052 9716
rect 7656 9707 7708 9716
rect 7656 9673 7665 9707
rect 7665 9673 7699 9707
rect 7699 9673 7708 9707
rect 7656 9664 7708 9673
rect 8024 9707 8076 9716
rect 8024 9673 8033 9707
rect 8033 9673 8067 9707
rect 8067 9673 8076 9707
rect 8024 9664 8076 9673
rect 4804 9596 4856 9648
rect 5172 9596 5224 9648
rect 11244 9596 11296 9648
rect 11520 9596 11572 9648
rect 5540 9392 5592 9444
rect 6368 9392 6420 9444
rect 6000 9324 6052 9376
rect 6184 9324 6236 9376
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 12716 8236 12768 8288
rect 13728 8236 13780 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 12532 8032 12584 8084
rect 13360 8032 13412 8084
rect 14004 7692 14056 7744
rect 14924 7692 14976 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 13912 7488 13964 7540
rect 15752 7488 15804 7540
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 4160 6808 4212 6860
rect 4252 6604 4304 6656
rect 5540 6604 5592 6656
rect 10324 6604 10376 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10140 6332 10192 6384
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10600 6264 10652 6316
rect 10140 6128 10192 6180
rect 4252 6060 4304 6112
rect 5632 6060 5684 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 8300 5856 8352 5908
rect 9312 5856 9364 5908
rect 10324 5856 10376 5908
rect 10232 5831 10284 5840
rect 10232 5797 10241 5831
rect 10241 5797 10275 5831
rect 10275 5797 10284 5831
rect 10232 5788 10284 5797
rect 9588 5720 9640 5772
rect 11428 5720 11480 5772
rect 9312 5652 9364 5704
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 8116 5312 8168 5364
rect 9588 5312 9640 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 9312 5108 9364 5160
rect 9496 4972 9548 5024
rect 10692 4972 10744 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 8208 4768 8260 4820
rect 5540 4700 5592 4752
rect 6828 4700 6880 4752
rect 5632 4632 5684 4684
rect 6460 4632 6512 4684
rect 9496 4768 9548 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 10232 4700 10284 4752
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 9312 4564 9364 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 9312 4224 9364 4276
rect 2964 4088 3016 4140
rect 4068 4088 4120 4140
rect 4988 4088 5040 4140
rect 5448 4088 5500 4140
rect 6828 4088 6880 4140
rect 10508 4224 10560 4276
rect 10600 4020 10652 4072
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 12440 3680 12492 3732
rect 12992 3680 13044 3732
rect 3976 3544 4028 3596
rect 6092 3544 6144 3596
rect 6644 3544 6696 3596
rect 4252 3451 4304 3460
rect 4252 3417 4261 3451
rect 4261 3417 4295 3451
rect 4295 3417 4304 3451
rect 4252 3408 4304 3417
rect 4528 3340 4580 3392
rect 6920 3340 6972 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 3332 3136 3384 3188
rect 3976 3136 4028 3188
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 5080 3136 5132 3188
rect 6092 3136 6144 3188
rect 6644 3136 6696 3188
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 2136 3068 2188 3120
rect 4620 3043 4672 3052
rect 3332 2932 3384 2984
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 7932 2932 7984 2984
rect 2872 2796 2924 2848
rect 6644 2796 6696 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 7288 2592 7340 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 8116 2592 8168 2644
rect 11152 2524 11204 2576
rect 11796 2524 11848 2576
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 1768 2252 1820 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 4804 552 4856 604
rect 5356 552 5408 604
rect 11336 552 11388 604
rect 11520 552 11572 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39522 2650 40000
rect 2516 39520 2650 39522
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39522 14978 40000
rect 14922 39520 15056 39522
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34542 244 39520
rect 584 34649 612 39520
rect 570 34640 626 34649
rect 570 34575 626 34584
rect 204 34536 256 34542
rect 204 34478 256 34484
rect 952 31521 980 39520
rect 1412 34542 1440 39520
rect 1780 35057 1808 39520
rect 1766 35048 1822 35057
rect 1766 34983 1822 34992
rect 1308 34536 1360 34542
rect 1308 34478 1360 34484
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 1320 33266 1348 34478
rect 1582 33416 1638 33425
rect 1582 33351 1638 33360
rect 1320 33238 1440 33266
rect 1412 32026 1440 33238
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 938 31512 994 31521
rect 938 31447 994 31456
rect 1596 27130 1624 33351
rect 1676 31884 1728 31890
rect 1676 31826 1728 31832
rect 1688 31142 1716 31826
rect 2148 31414 2176 39520
rect 2516 39494 2636 39520
rect 2136 31408 2188 31414
rect 2136 31350 2188 31356
rect 2516 31226 2544 39494
rect 2870 34640 2926 34649
rect 2870 34575 2926 34584
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2792 32570 2820 34478
rect 2780 32564 2832 32570
rect 2780 32506 2832 32512
rect 2884 32026 2912 34575
rect 2976 34542 3004 39520
rect 3344 35193 3372 39520
rect 3804 37754 3832 39520
rect 3804 37726 4016 37754
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3330 35184 3386 35193
rect 3330 35119 3386 35128
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 2964 34536 3016 34542
rect 2964 34478 3016 34484
rect 3988 34105 4016 37726
rect 4172 34542 4200 39520
rect 4342 35048 4398 35057
rect 4342 34983 4398 34992
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 4160 34536 4212 34542
rect 4160 34478 4212 34484
rect 3974 34096 4030 34105
rect 3974 34031 4030 34040
rect 3974 33960 4030 33969
rect 3974 33895 4030 33904
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 2870 31512 2926 31521
rect 2870 31447 2872 31456
rect 2924 31447 2926 31456
rect 2872 31418 2924 31424
rect 2516 31198 2636 31226
rect 1676 31136 1728 31142
rect 1676 31078 1728 31084
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 1584 27124 1636 27130
rect 1584 27066 1636 27072
rect 1688 10305 1716 31078
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2424 19310 2452 22034
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2516 12986 2544 31078
rect 2608 22098 2636 31198
rect 2688 26784 2740 26790
rect 2740 26744 2820 26772
rect 2688 26726 2740 26732
rect 2792 24682 2820 26744
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2780 24676 2832 24682
rect 2780 24618 2832 24624
rect 2976 24614 3004 24754
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2596 22092 2648 22098
rect 2596 22034 2648 22040
rect 2976 20097 3004 24550
rect 2962 20088 3018 20097
rect 2962 20023 3018 20032
rect 2688 19304 2740 19310
rect 3068 19281 3096 32302
rect 3240 31884 3292 31890
rect 3240 31826 3292 31832
rect 3252 31142 3280 31826
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 3424 31136 3476 31142
rect 3424 31078 3476 31084
rect 3148 19304 3200 19310
rect 2688 19246 2740 19252
rect 3054 19272 3110 19281
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1398 10024 1454 10033
rect 1398 9959 1454 9968
rect 938 2952 994 2961
rect 938 2887 994 2896
rect 570 2816 626 2825
rect 570 2751 626 2760
rect 202 1456 258 1465
rect 202 1391 258 1400
rect 216 480 244 1391
rect 584 480 612 2751
rect 952 480 980 2887
rect 1412 2514 1440 9959
rect 2700 9704 2728 19246
rect 3148 19246 3200 19252
rect 3054 19207 3110 19216
rect 3160 18290 3188 19246
rect 3252 18873 3280 31078
rect 3332 26240 3384 26246
rect 3332 26182 3384 26188
rect 3344 25498 3372 26182
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3344 24614 3372 25434
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 3436 21049 3464 31078
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3528 24070 3556 24686
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3528 21690 3556 24006
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3422 21040 3478 21049
rect 3422 20975 3478 20984
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3514 20088 3570 20097
rect 3514 20023 3570 20032
rect 3238 18864 3294 18873
rect 3238 18799 3294 18808
rect 3528 18426 3556 20023
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3882 19408 3938 19417
rect 3882 19343 3938 19352
rect 3896 19310 3924 19343
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3240 18148 3292 18154
rect 3240 18090 3292 18096
rect 3252 17882 3280 18090
rect 3422 18048 3478 18057
rect 3422 17983 3478 17992
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3238 16552 3294 16561
rect 3238 16487 3294 16496
rect 2424 9676 2728 9704
rect 2424 4185 2452 9676
rect 2410 4176 2466 4185
rect 2410 4111 2466 4120
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2594 3496 2650 3505
rect 2594 3431 2650 3440
rect 2136 3120 2188 3126
rect 1490 3088 1546 3097
rect 2136 3062 2188 3068
rect 1490 3023 1546 3032
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1504 1170 1532 3023
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1596 1465 1624 2246
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 1412 1142 1532 1170
rect 1412 480 1440 1142
rect 1780 480 1808 2246
rect 2148 480 2176 3062
rect 2608 480 2636 3431
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 2884 2854 2912 2887
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2976 480 3004 4082
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 3068 2650 3096 2751
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3252 1578 3280 16487
rect 3330 5672 3386 5681
rect 3330 5607 3386 5616
rect 3344 3194 3372 5607
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3344 2990 3372 3130
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3436 2650 3464 17983
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3514 17232 3570 17241
rect 3514 17167 3570 17176
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3528 1986 3556 17167
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3988 3602 4016 33895
rect 4080 32586 4108 34478
rect 4080 32570 4200 32586
rect 4080 32564 4212 32570
rect 4080 32558 4160 32564
rect 4160 32506 4212 32512
rect 4356 32026 4384 34983
rect 4436 32360 4488 32366
rect 4436 32302 4488 32308
rect 4344 32020 4396 32026
rect 4344 31962 4396 31968
rect 4344 31748 4396 31754
rect 4344 31690 4396 31696
rect 4356 31142 4384 31690
rect 4344 31136 4396 31142
rect 4344 31078 4396 31084
rect 4066 30832 4122 30841
rect 4066 30767 4068 30776
rect 4120 30767 4122 30776
rect 4068 30738 4120 30744
rect 4080 30394 4108 30738
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4172 27554 4200 30534
rect 4080 27526 4200 27554
rect 4080 4146 4108 27526
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 4172 22681 4200 27406
rect 4158 22672 4214 22681
rect 4158 22607 4214 22616
rect 4356 10577 4384 31078
rect 4448 27470 4476 32302
rect 4540 31482 4568 39520
rect 4528 31476 4580 31482
rect 4528 31418 4580 31424
rect 5000 31385 5028 39520
rect 4986 31376 5042 31385
rect 4986 31311 5042 31320
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4724 22137 4752 31078
rect 5368 30705 5396 39520
rect 5540 34536 5592 34542
rect 5540 34478 5592 34484
rect 5552 32026 5580 34478
rect 5736 32609 5764 39520
rect 5722 32600 5778 32609
rect 5722 32535 5778 32544
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 5460 31770 5488 31826
rect 5460 31742 5580 31770
rect 5552 31142 5580 31742
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5354 30696 5410 30705
rect 5354 30631 5410 30640
rect 5446 29608 5502 29617
rect 5446 29543 5502 29552
rect 5170 28520 5226 28529
rect 5170 28455 5226 28464
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 5000 26042 5028 26250
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4710 22128 4766 22137
rect 4710 22063 4766 22072
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4816 21350 4844 21830
rect 5000 21554 5028 25978
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4816 21146 4844 21286
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4908 20806 4936 21286
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 5078 17776 5134 17785
rect 5078 17711 5134 17720
rect 4342 10568 4398 10577
rect 4342 10503 4398 10512
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 6769 4200 6802
rect 4158 6760 4214 6769
rect 4158 6695 4214 6704
rect 4172 6458 4200 6695
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4264 6118 4292 6598
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4158 4176 4214 4185
rect 4068 4140 4120 4146
rect 4158 4111 4214 4120
rect 4068 4082 4120 4088
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3988 3194 4016 3538
rect 4172 3194 4200 4111
rect 4250 3496 4306 3505
rect 4250 3431 4252 3440
rect 4304 3431 4306 3440
rect 4252 3402 4304 3408
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4250 3088 4306 3097
rect 4250 3023 4306 3032
rect 4264 2650 4292 3023
rect 4342 2952 4398 2961
rect 4342 2887 4398 2896
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3528 1958 3832 1986
rect 3252 1550 3372 1578
rect 3344 480 3372 1550
rect 3804 480 3832 1958
rect 4356 1714 4384 2887
rect 4172 1686 4384 1714
rect 4172 480 4200 1686
rect 4540 480 4568 3334
rect 4618 3088 4674 3097
rect 4618 3023 4620 3032
rect 4672 3023 4674 3032
rect 4620 2994 4672 3000
rect 4710 2544 4766 2553
rect 4710 2479 4712 2488
rect 4764 2479 4766 2488
rect 4712 2450 4764 2456
rect 4816 610 4844 9590
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 604 4856 610
rect 4804 546 4856 552
rect 5000 480 5028 4082
rect 5092 3194 5120 17711
rect 5184 9654 5212 28455
rect 5264 27328 5316 27334
rect 5264 27270 5316 27276
rect 5276 26518 5304 27270
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5264 26512 5316 26518
rect 5264 26454 5316 26460
rect 5368 26042 5396 26522
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5368 19174 5396 21354
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5368 18154 5396 19110
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5460 4146 5488 29543
rect 5552 11257 5580 31078
rect 6196 30161 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6656 32473 6684 37726
rect 6932 34626 6960 39520
rect 7010 35184 7066 35193
rect 7010 35119 7066 35128
rect 6840 34598 6960 34626
rect 6642 32464 6698 32473
rect 6642 32399 6698 32408
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6840 32026 6868 34598
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6460 31884 6512 31890
rect 6460 31826 6512 31832
rect 6472 31482 6500 31826
rect 7024 31482 7052 35119
rect 7102 34640 7158 34649
rect 7102 34575 7158 34584
rect 6460 31476 6512 31482
rect 7012 31476 7064 31482
rect 6512 31436 6684 31464
rect 6460 31418 6512 31424
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6182 30152 6238 30161
rect 6182 30087 6238 30096
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6552 27056 6604 27062
rect 6552 26998 6604 27004
rect 6564 26772 6592 26998
rect 6656 26926 6684 31436
rect 7012 31418 7064 31424
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6840 27554 6868 27814
rect 6920 27600 6972 27606
rect 6840 27548 6920 27554
rect 6840 27542 6972 27548
rect 6840 27526 6960 27542
rect 6828 27464 6880 27470
rect 6826 27432 6828 27441
rect 6880 27432 6882 27441
rect 6826 27367 6882 27376
rect 6840 27062 6868 27367
rect 6932 27130 6960 27526
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6644 26920 6696 26926
rect 6644 26862 6696 26868
rect 6828 26784 6880 26790
rect 6564 26744 6684 26772
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 5632 26512 5684 26518
rect 5632 26454 5684 26460
rect 5644 26042 5672 26454
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 6182 25936 6238 25945
rect 6182 25871 6238 25880
rect 5722 24168 5778 24177
rect 5722 24103 5778 24112
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 20058 5672 20742
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5630 19272 5686 19281
rect 5630 19207 5632 19216
rect 5684 19207 5686 19216
rect 5632 19178 5684 19184
rect 5538 11248 5594 11257
rect 5538 11183 5594 11192
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5644 10062 5672 10231
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 6662 5580 9386
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 4758 5580 6598
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5644 4690 5672 6054
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5092 2990 5120 3130
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5356 604 5408 610
rect 5356 546 5408 552
rect 5368 480 5396 546
rect 5736 480 5764 24103
rect 6090 22128 6146 22137
rect 6090 22063 6146 22072
rect 6104 21010 6132 22063
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 5920 20262 5948 20946
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5828 19310 5856 19926
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5828 18970 5856 19246
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5828 3074 5856 17206
rect 5920 7857 5948 20198
rect 6104 19990 6132 20538
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 6012 19514 6040 19858
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 18426 6040 19246
rect 6104 18970 6132 19790
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6104 18057 6132 18090
rect 6090 18048 6146 18057
rect 6090 17983 6146 17992
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 10033 6040 10066
rect 5998 10024 6054 10033
rect 5998 9959 6054 9968
rect 6012 9722 6040 9959
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5906 7848 5962 7857
rect 5906 7783 5962 7792
rect 6012 4729 6040 9318
rect 5998 4720 6054 4729
rect 5998 4655 6054 4664
rect 6104 3602 6132 17818
rect 6196 17270 6224 25871
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20602 6500 20878
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6564 18154 6592 18770
rect 6552 18148 6604 18154
rect 6552 18090 6604 18096
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6196 10470 6224 10610
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10146 6224 10406
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6196 10118 6408 10146
rect 6380 10062 6408 10118
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6196 9382 6224 9998
rect 6380 9450 6408 9998
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 4282 6500 4626
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6656 3602 6684 26744
rect 6828 26726 6880 26732
rect 6840 26586 6868 26726
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6748 20330 6776 20946
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6748 20058 6776 20266
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6734 18864 6790 18873
rect 6734 18799 6790 18808
rect 6748 18766 6776 18799
rect 6736 18760 6788 18766
rect 6736 18702 6788 18708
rect 6748 18086 6776 18702
rect 6736 18080 6788 18086
rect 6734 18048 6736 18057
rect 6788 18048 6790 18057
rect 6734 17983 6790 17992
rect 6932 17882 6960 26522
rect 7116 19718 7144 34575
rect 7392 32337 7420 39520
rect 7760 34542 7788 39520
rect 8220 34626 8248 39520
rect 8128 34598 8248 34626
rect 7748 34536 7800 34542
rect 7748 34478 7800 34484
rect 7654 33552 7710 33561
rect 7654 33487 7710 33496
rect 7562 33280 7618 33289
rect 7562 33215 7618 33224
rect 7470 32872 7526 32881
rect 7470 32807 7526 32816
rect 7484 32570 7512 32807
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7378 32328 7434 32337
rect 7484 32298 7512 32506
rect 7378 32263 7434 32272
rect 7472 32292 7524 32298
rect 7472 32234 7524 32240
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7300 31822 7328 32166
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 7380 31136 7432 31142
rect 7378 31104 7380 31113
rect 7432 31104 7434 31113
rect 7378 31039 7434 31048
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 7208 26994 7236 27406
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7208 26314 7236 26930
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 20602 7236 26250
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7116 19174 7144 19654
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 11506 6960 11562
rect 6840 11478 6960 11506
rect 6840 10810 6868 11478
rect 7116 11234 7144 19110
rect 7300 18630 7328 19858
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 17785 7328 18566
rect 7286 17776 7342 17785
rect 7286 17711 7342 17720
rect 7392 16561 7420 21082
rect 7378 16552 7434 16561
rect 7378 16487 7434 16496
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6920 11212 6972 11218
rect 7116 11206 7236 11234
rect 6920 11154 6972 11160
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6932 10538 6960 11154
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7024 10606 7052 11086
rect 7116 10742 7144 11086
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7102 10568 7158 10577
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6736 10464 6788 10470
rect 6734 10432 6736 10441
rect 6788 10432 6790 10441
rect 6734 10367 6790 10376
rect 6932 10266 6960 10474
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7024 9994 7052 10542
rect 7102 10503 7158 10512
rect 7116 10470 7144 10503
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7116 9926 7144 10406
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6840 4146 6868 4694
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6104 3194 6132 3538
rect 6656 3194 6684 3538
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 5828 3046 6224 3074
rect 6196 480 6224 3046
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 1442 6684 2790
rect 6564 1414 6684 1442
rect 6564 480 6592 1414
rect 6932 480 6960 3334
rect 7208 2553 7236 11206
rect 7288 10464 7340 10470
rect 7286 10432 7288 10441
rect 7340 10432 7342 10441
rect 7286 10367 7342 10376
rect 7392 10266 7420 12922
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 3890 7328 9862
rect 7392 9382 7420 10202
rect 7484 10033 7512 30874
rect 7576 19922 7604 33215
rect 7668 26926 7696 33487
rect 8022 32464 8078 32473
rect 8022 32399 8078 32408
rect 8036 32026 8064 32399
rect 8024 32020 8076 32026
rect 8024 31962 8076 31968
rect 7840 31884 7892 31890
rect 7840 31826 7892 31832
rect 7748 31816 7800 31822
rect 7748 31758 7800 31764
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 26586 7696 26862
rect 7656 26580 7708 26586
rect 7656 26522 7708 26528
rect 7760 21146 7788 31758
rect 7852 31142 7880 31826
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7746 21040 7802 21049
rect 7746 20975 7802 20984
rect 7760 19922 7788 20975
rect 7852 20913 7880 31078
rect 8128 30938 8156 34598
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8220 31249 8248 34478
rect 8206 31240 8262 31249
rect 8588 31226 8616 39520
rect 8956 37890 8984 39520
rect 8206 31175 8262 31184
rect 8404 31198 8616 31226
rect 8680 37862 8984 37890
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 7932 26784 7984 26790
rect 7932 26726 7984 26732
rect 7838 20904 7894 20913
rect 7838 20839 7894 20848
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7760 19174 7788 19858
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7852 19378 7880 19790
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 12186 7788 19110
rect 7852 18970 7880 19314
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7944 17785 7972 26726
rect 8116 20256 8168 20262
rect 8114 20224 8116 20233
rect 8168 20224 8170 20233
rect 8114 20159 8170 20168
rect 8128 19417 8156 20159
rect 8114 19408 8170 19417
rect 8114 19343 8170 19352
rect 8404 18154 8432 31198
rect 8680 31090 8708 37862
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9416 34649 9444 39520
rect 9402 34640 9458 34649
rect 9402 34575 9458 34584
rect 9586 34640 9642 34649
rect 9586 34575 9642 34584
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 9600 32570 9628 34575
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 9600 32366 9628 32506
rect 9588 32360 9640 32366
rect 9588 32302 9640 32308
rect 8852 32224 8904 32230
rect 8852 32166 8904 32172
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 8588 31062 8708 31090
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8496 19718 8524 20266
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8482 18048 8538 18057
rect 8482 17983 8538 17992
rect 7930 17776 7986 17785
rect 7930 17711 7986 17720
rect 7760 12158 7880 12186
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11626 7788 12038
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7668 9722 7696 10066
rect 7852 10033 7880 12158
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 11257 8064 11494
rect 8022 11248 8078 11257
rect 8022 11183 8078 11192
rect 8128 11150 8156 11698
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7838 10024 7894 10033
rect 7838 9959 7894 9968
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9722 8064 9930
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 4049 7420 9318
rect 7668 5681 7696 9658
rect 8128 5930 8156 11086
rect 8496 7562 8524 17983
rect 8588 10130 8616 31062
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8496 7534 8616 7562
rect 8128 5914 8340 5930
rect 8128 5908 8352 5914
rect 8128 5902 8300 5908
rect 7654 5672 7710 5681
rect 7654 5607 7710 5616
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7378 4040 7434 4049
rect 7378 3975 7434 3984
rect 7300 3862 7420 3890
rect 7392 2666 7420 3862
rect 7746 3632 7802 3641
rect 7746 3567 7802 3576
rect 7470 2952 7526 2961
rect 7654 2952 7710 2961
rect 7470 2887 7526 2896
rect 7576 2910 7654 2938
rect 7300 2650 7420 2666
rect 7484 2650 7512 2887
rect 7288 2644 7420 2650
rect 7340 2638 7420 2644
rect 7472 2644 7524 2650
rect 7288 2586 7340 2592
rect 7472 2586 7524 2592
rect 7194 2544 7250 2553
rect 7576 2530 7604 2910
rect 7654 2887 7710 2896
rect 7194 2479 7250 2488
rect 7392 2502 7604 2530
rect 7392 480 7420 2502
rect 7760 480 7788 3567
rect 7930 3496 7986 3505
rect 7930 3431 7986 3440
rect 7944 3194 7972 3431
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7944 2990 7972 3130
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8128 2650 8156 5306
rect 8220 4826 8248 5902
rect 8300 5850 8352 5856
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8206 4720 8262 4729
rect 8206 4655 8262 4664
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8220 480 8248 4655
rect 8588 480 8616 7534
rect 8772 7426 8800 19178
rect 8864 17241 8892 32166
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9692 31498 9720 32166
rect 9600 31470 9720 31498
rect 9600 31226 9628 31470
rect 9680 31408 9732 31414
rect 9678 31376 9680 31385
rect 9732 31376 9734 31385
rect 9678 31311 9734 31320
rect 9784 31226 9812 39520
rect 9862 34096 9918 34105
rect 9862 34031 9918 34040
rect 9876 32026 9904 34031
rect 10152 33289 10180 39520
rect 10612 33969 10640 39520
rect 10690 34912 10746 34921
rect 10690 34847 10746 34856
rect 10598 33960 10654 33969
rect 10598 33895 10654 33904
rect 10704 33538 10732 34847
rect 10874 34776 10930 34785
rect 10874 34711 10930 34720
rect 10612 33510 10732 33538
rect 10138 33280 10194 33289
rect 10138 33215 10194 33224
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 10322 31376 10378 31385
rect 10322 31311 10378 31320
rect 9600 31198 9720 31226
rect 9784 31198 10272 31226
rect 9310 31104 9366 31113
rect 9310 31039 9366 31048
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8850 17232 8906 17241
rect 8850 17167 8906 17176
rect 9324 16561 9352 31039
rect 9692 29617 9720 31198
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9678 29608 9734 29617
rect 9678 29543 9734 29552
rect 9968 24993 9996 31078
rect 10140 30796 10192 30802
rect 10140 30738 10192 30744
rect 10046 30696 10102 30705
rect 10046 30631 10048 30640
rect 10100 30631 10102 30640
rect 10048 30602 10100 30608
rect 10152 30054 10180 30738
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10060 28529 10088 29990
rect 10046 28520 10102 28529
rect 10046 28455 10102 28464
rect 10244 28098 10272 31198
rect 10336 30841 10364 31311
rect 10520 31142 10548 31826
rect 10612 31362 10640 33510
rect 10690 33416 10746 33425
rect 10690 33351 10746 33360
rect 10704 32570 10732 33351
rect 10692 32564 10744 32570
rect 10692 32506 10744 32512
rect 10704 32366 10732 32506
rect 10782 32464 10838 32473
rect 10782 32399 10838 32408
rect 10692 32360 10744 32366
rect 10692 32302 10744 32308
rect 10612 31334 10732 31362
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10322 30832 10378 30841
rect 10322 30767 10378 30776
rect 10704 28218 10732 31334
rect 10796 28762 10824 32399
rect 10888 30326 10916 34711
rect 10980 31385 11008 39520
rect 11150 35184 11206 35193
rect 11150 35119 11206 35128
rect 10966 31376 11022 31385
rect 10966 31311 11022 31320
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10980 30954 11008 31078
rect 10980 30926 11100 30954
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10244 28070 10732 28098
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 9954 24984 10010 24993
rect 9954 24919 10010 24928
rect 10520 24177 10548 27814
rect 10506 24168 10562 24177
rect 10506 24103 10562 24112
rect 9678 22672 9734 22681
rect 9678 22607 9734 22616
rect 9310 16552 9366 16561
rect 9310 16487 9366 16496
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9692 12730 9720 22607
rect 10322 20904 10378 20913
rect 10322 20839 10378 20848
rect 9862 20224 9918 20233
rect 9862 20159 9918 20168
rect 9876 19922 9904 20159
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9876 19174 9904 19858
rect 10060 19514 10088 19858
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9954 19408 10010 19417
rect 9954 19343 10010 19352
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 14074 9904 19110
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9968 13530 9996 19343
rect 10060 13734 10088 19450
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 13870 10180 14214
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 12782 9904 13330
rect 10060 13258 10088 13670
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10060 12986 10088 13194
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9864 12776 9916 12782
rect 9692 12702 9812 12730
rect 9864 12718 9916 12724
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11898 8892 12038
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9600 11898 9628 12582
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 8864 11694 8892 11834
rect 9784 11694 9812 12702
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11082 9812 11494
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9770 10432 9826 10441
rect 9770 10367 9826 10376
rect 9494 9888 9550 9897
rect 8956 9820 9252 9840
rect 9494 9823 9550 9832
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8772 7398 9444 7426
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5710 9352 5850
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5166 9352 5646
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9324 4622 9352 5102
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9324 4282 9352 4558
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 8850 4040 8906 4049
rect 8850 3975 8906 3984
rect 8864 1986 8892 3975
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1958 8984 1986
rect 8956 480 8984 1958
rect 9416 480 9444 7398
rect 9508 5030 9536 9823
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5370 9628 5714
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4826 9536 4966
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9784 480 9812 10367
rect 9876 6458 9904 12718
rect 10152 11762 10180 13806
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10046 10024 10102 10033
rect 10046 9959 10102 9968
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10060 4706 10088 9959
rect 10152 6390 10180 11698
rect 10244 10033 10272 14010
rect 10230 10024 10286 10033
rect 10230 9959 10286 9968
rect 10336 6746 10364 20839
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12646 10456 13262
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10704 10577 10732 28070
rect 10888 27878 10916 28562
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 10888 22137 10916 27814
rect 10980 23633 11008 29990
rect 11072 29186 11100 30926
rect 11164 29714 11192 35119
rect 11348 32881 11376 39520
rect 11808 37754 11836 39520
rect 11440 37726 11836 37754
rect 11440 34649 11468 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11426 34640 11482 34649
rect 11426 34575 11482 34584
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11334 32872 11390 32881
rect 11334 32807 11390 32816
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 12176 31226 12204 39520
rect 12544 33561 12572 39520
rect 12530 33552 12586 33561
rect 12530 33487 12586 33496
rect 13004 33425 13032 39520
rect 13082 35048 13138 35057
rect 13082 34983 13138 34992
rect 12990 33416 13046 33425
rect 12990 33351 13046 33360
rect 13096 32570 13124 34983
rect 13372 34785 13400 39520
rect 13740 34921 13768 39520
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 13726 34912 13782 34921
rect 13726 34847 13782 34856
rect 13358 34776 13414 34785
rect 13358 34711 13414 34720
rect 13450 34640 13506 34649
rect 13450 34575 13506 34584
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 13096 32366 13124 32506
rect 13084 32360 13136 32366
rect 12530 32328 12586 32337
rect 13084 32302 13136 32308
rect 12530 32263 12586 32272
rect 12544 32026 12572 32263
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 11440 31198 12204 31226
rect 12530 31240 12586 31249
rect 11334 30152 11390 30161
rect 11334 30087 11390 30096
rect 11348 30054 11376 30087
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 11164 29306 11192 29650
rect 11336 29504 11388 29510
rect 11336 29446 11388 29452
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 11072 29158 11192 29186
rect 10966 23624 11022 23633
rect 10966 23559 11022 23568
rect 10874 22128 10930 22137
rect 10874 22063 10930 22072
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10244 6718 10364 6746
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10152 4826 10180 6122
rect 10244 5846 10272 6718
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6322 10364 6598
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10336 5914 10364 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10244 4758 10272 5782
rect 10612 5370 10640 6258
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10598 5128 10654 5137
rect 10598 5063 10654 5072
rect 10612 4826 10640 5063
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10232 4752 10284 4758
rect 10060 4678 10180 4706
rect 10232 4694 10284 4700
rect 10152 480 10180 4678
rect 10244 4049 10272 4694
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10520 4282 10548 4626
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10612 4078 10640 4762
rect 10704 4622 10732 4966
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10600 4072 10652 4078
rect 10230 4040 10286 4049
rect 10600 4014 10652 4020
rect 10230 3975 10286 3984
rect 10612 3505 10640 4014
rect 10598 3496 10654 3505
rect 10598 3431 10654 3440
rect 10598 3088 10654 3097
rect 10598 3023 10654 3032
rect 10612 480 10640 3023
rect 10980 480 11008 11630
rect 11164 2582 11192 29158
rect 11348 25945 11376 29446
rect 11334 25936 11390 25945
rect 11334 25871 11390 25880
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 11256 9654 11284 16487
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11440 5778 11468 31198
rect 12530 31175 12586 31184
rect 12544 31142 12572 31175
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 12254 30016 12310 30025
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11532 610 11560 9590
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11992 3505 12020 29990
rect 12254 29951 12310 29960
rect 12268 25498 12296 29951
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12084 24614 12112 25298
rect 12438 24984 12494 24993
rect 12438 24919 12494 24928
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 12084 19417 12112 24550
rect 12070 19408 12126 19417
rect 12070 19343 12126 19352
rect 12162 11248 12218 11257
rect 12162 11183 12218 11192
rect 11978 3496 12034 3505
rect 11978 3431 12034 3440
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11336 604 11388 610
rect 11336 546 11388 552
rect 11520 604 11572 610
rect 11520 546 11572 552
rect 11348 480 11376 546
rect 11808 480 11836 2518
rect 12176 480 12204 11183
rect 12452 3738 12480 24919
rect 12530 23624 12586 23633
rect 12530 23559 12586 23568
rect 12544 8090 12572 23559
rect 12636 22098 12664 32166
rect 13464 31890 13492 34575
rect 13452 31884 13504 31890
rect 13452 31826 13504 31832
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 13004 31142 13032 31690
rect 13464 31482 13492 31826
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 12714 22128 12770 22137
rect 12624 22092 12676 22098
rect 12714 22063 12770 22072
rect 12624 22034 12676 22040
rect 12728 8294 12756 22063
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12530 7848 12586 7857
rect 12530 7783 12586 7792
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 480 12572 7783
rect 12820 3641 12848 21966
rect 13004 3913 13032 31078
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 12990 3904 13046 3913
rect 12990 3839 13046 3848
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12806 3632 12862 3641
rect 12806 3567 12862 3576
rect 13004 480 13032 3674
rect 13372 480 13400 8026
rect 13648 2961 13676 31622
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13634 2952 13690 2961
rect 13634 2887 13690 2896
rect 13740 480 13768 8230
rect 13832 5137 13860 37742
rect 14200 35193 14228 39520
rect 14568 37806 14596 39520
rect 14936 39494 15056 39520
rect 14556 37800 14608 37806
rect 14556 37742 14608 37748
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14186 35184 14242 35193
rect 14186 35119 14242 35128
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 13912 31272 13964 31278
rect 13912 31214 13964 31220
rect 13924 7546 13952 31214
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 15028 27441 15056 39494
rect 15396 34649 15424 39520
rect 15764 35057 15792 39520
rect 15750 35048 15806 35057
rect 15750 34983 15806 34992
rect 15382 34640 15438 34649
rect 15382 34575 15438 34584
rect 15014 27432 15070 27441
rect 15014 27367 15070 27376
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14002 17776 14058 17785
rect 14002 17711 14058 17720
rect 14016 7750 14044 17711
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 13818 5128 13874 5137
rect 13818 5063 13874 5072
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14186 3496 14242 3505
rect 14186 3431 14242 3440
rect 14200 480 14228 3431
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 3975
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 7686
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15396 480 15424 3839
rect 15764 480 15792 7482
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 570 34584 626 34640
rect 1766 34992 1822 35048
rect 1582 33360 1638 33416
rect 938 31456 994 31512
rect 2870 34584 2926 34640
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3330 35128 3386 35184
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4342 34992 4398 35048
rect 3974 34040 4030 34096
rect 3974 33904 4030 33960
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 2870 31476 2926 31512
rect 2870 31456 2872 31476
rect 2872 31456 2924 31476
rect 2924 31456 2926 31476
rect 2962 20032 3018 20088
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 1674 10240 1730 10296
rect 1398 9968 1454 10024
rect 938 2896 994 2952
rect 570 2760 626 2816
rect 202 1400 258 1456
rect 3054 19216 3110 19272
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3422 20984 3478 21040
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3514 20032 3570 20088
rect 3238 18808 3294 18864
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3882 19352 3938 19408
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3422 17992 3478 18048
rect 3238 16496 3294 16552
rect 2410 4120 2466 4176
rect 2594 3440 2650 3496
rect 1490 3032 1546 3088
rect 1582 1400 1638 1456
rect 2870 2896 2926 2952
rect 3054 2760 3110 2816
rect 3330 5616 3386 5672
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3514 17176 3570 17232
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4066 30796 4122 30832
rect 4066 30776 4068 30796
rect 4068 30776 4120 30796
rect 4120 30776 4122 30796
rect 4158 22616 4214 22672
rect 4986 31320 5042 31376
rect 5722 32544 5778 32600
rect 5354 30640 5410 30696
rect 5446 29552 5502 29608
rect 5170 28464 5226 28520
rect 4710 22072 4766 22128
rect 5078 17720 5134 17776
rect 4342 10512 4398 10568
rect 4158 6704 4214 6760
rect 4158 4120 4214 4176
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4250 3460 4306 3496
rect 4250 3440 4252 3460
rect 4252 3440 4304 3460
rect 4304 3440 4306 3460
rect 4250 3032 4306 3088
rect 4342 2896 4398 2952
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4618 3052 4674 3088
rect 4618 3032 4620 3052
rect 4620 3032 4672 3052
rect 4672 3032 4674 3052
rect 4710 2508 4766 2544
rect 4710 2488 4712 2508
rect 4712 2488 4764 2508
rect 4764 2488 4766 2508
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 7010 35128 7066 35184
rect 6642 32408 6698 32464
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 7102 34584 7158 34640
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6182 30096 6238 30152
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6826 27412 6828 27432
rect 6828 27412 6880 27432
rect 6880 27412 6882 27432
rect 6826 27376 6882 27412
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6182 25880 6238 25936
rect 5722 24112 5778 24168
rect 5630 19236 5686 19272
rect 5630 19216 5632 19236
rect 5632 19216 5684 19236
rect 5684 19216 5686 19236
rect 5538 11192 5594 11248
rect 5630 10240 5686 10296
rect 6090 22072 6146 22128
rect 6090 17992 6146 18048
rect 5998 9968 6054 10024
rect 5906 7792 5962 7848
rect 5998 4664 6054 4720
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6734 18808 6790 18864
rect 6734 18028 6736 18048
rect 6736 18028 6788 18048
rect 6788 18028 6790 18048
rect 6734 17992 6790 18028
rect 7654 33496 7710 33552
rect 7562 33224 7618 33280
rect 7470 32816 7526 32872
rect 7378 32272 7434 32328
rect 7378 31084 7380 31104
rect 7380 31084 7432 31104
rect 7432 31084 7434 31104
rect 7378 31048 7434 31084
rect 7286 17720 7342 17776
rect 7378 16496 7434 16552
rect 6734 10412 6736 10432
rect 6736 10412 6788 10432
rect 6788 10412 6790 10432
rect 6734 10376 6790 10412
rect 7102 10512 7158 10568
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7286 10412 7288 10432
rect 7288 10412 7340 10432
rect 7340 10412 7342 10432
rect 7286 10376 7342 10412
rect 8022 32408 8078 32464
rect 7746 20984 7802 21040
rect 8206 31184 8262 31240
rect 7838 20848 7894 20904
rect 8114 20204 8116 20224
rect 8116 20204 8168 20224
rect 8168 20204 8170 20224
rect 8114 20168 8170 20204
rect 8114 19352 8170 19408
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 9402 34584 9458 34640
rect 9586 34584 9642 34640
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8482 17992 8538 18048
rect 7930 17720 7986 17776
rect 7470 9968 7526 10024
rect 8022 11192 8078 11248
rect 7838 9968 7894 10024
rect 7654 5616 7710 5672
rect 7378 3984 7434 4040
rect 7746 3576 7802 3632
rect 7470 2896 7526 2952
rect 7194 2488 7250 2544
rect 7654 2896 7710 2952
rect 7930 3440 7986 3496
rect 8206 4664 8262 4720
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 9678 31356 9680 31376
rect 9680 31356 9732 31376
rect 9732 31356 9734 31376
rect 9678 31320 9734 31356
rect 9862 34040 9918 34096
rect 10690 34856 10746 34912
rect 10598 33904 10654 33960
rect 10874 34720 10930 34776
rect 10138 33224 10194 33280
rect 10322 31320 10378 31376
rect 9310 31048 9366 31104
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8850 17176 8906 17232
rect 9678 29552 9734 29608
rect 10046 30660 10102 30696
rect 10046 30640 10048 30660
rect 10048 30640 10100 30660
rect 10100 30640 10102 30660
rect 10046 28464 10102 28520
rect 10690 33360 10746 33416
rect 10782 32408 10838 32464
rect 10322 30776 10378 30832
rect 11150 35128 11206 35184
rect 10966 31320 11022 31376
rect 9954 24928 10010 24984
rect 10506 24112 10562 24168
rect 9678 22616 9734 22672
rect 9310 16496 9366 16552
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 10322 20848 10378 20904
rect 9862 20168 9918 20224
rect 9954 19352 10010 19408
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 9770 10376 9826 10432
rect 9494 9832 9550 9888
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8850 3984 8906 4040
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10046 9968 10102 10024
rect 10230 9968 10286 10024
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11426 34584 11482 34640
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11334 32816 11390 32872
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 12530 33496 12586 33552
rect 13082 34992 13138 35048
rect 12990 33360 13046 33416
rect 13726 34856 13782 34912
rect 13358 34720 13414 34776
rect 13450 34584 13506 34640
rect 12530 32272 12586 32328
rect 11334 30096 11390 30152
rect 10966 23568 11022 23624
rect 10874 22072 10930 22128
rect 10690 10512 10746 10568
rect 10598 5072 10654 5128
rect 10230 3984 10286 4040
rect 10598 3440 10654 3496
rect 10598 3032 10654 3088
rect 11334 25880 11390 25936
rect 11242 16496 11298 16552
rect 12530 31184 12586 31240
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 12254 29960 12310 30016
rect 12438 24928 12494 24984
rect 12070 19352 12126 19408
rect 12162 11192 12218 11248
rect 11978 3440 12034 3496
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12530 23568 12586 23624
rect 12714 22072 12770 22128
rect 12530 7792 12586 7848
rect 12990 3848 13046 3904
rect 12806 3576 12862 3632
rect 13634 2896 13690 2952
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14186 35128 14242 35184
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 15750 34992 15806 35048
rect 15382 34584 15438 34640
rect 15014 27376 15070 27432
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14002 17720 14058 17776
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 13818 5072 13874 5128
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14646 3984 14702 4040
rect 14186 3440 14242 3496
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15382 3848 15438 3904
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3325 35186 3391 35189
rect 7005 35186 7071 35189
rect 3325 35184 7071 35186
rect 3325 35128 3330 35184
rect 3386 35128 7010 35184
rect 7066 35128 7071 35184
rect 3325 35126 7071 35128
rect 3325 35123 3391 35126
rect 7005 35123 7071 35126
rect 11145 35186 11211 35189
rect 14181 35186 14247 35189
rect 11145 35184 14247 35186
rect 11145 35128 11150 35184
rect 11206 35128 14186 35184
rect 14242 35128 14247 35184
rect 11145 35126 14247 35128
rect 11145 35123 11211 35126
rect 14181 35123 14247 35126
rect 1761 35050 1827 35053
rect 4337 35050 4403 35053
rect 1761 35048 4403 35050
rect 1761 34992 1766 35048
rect 1822 34992 4342 35048
rect 4398 34992 4403 35048
rect 1761 34990 4403 34992
rect 1761 34987 1827 34990
rect 4337 34987 4403 34990
rect 13077 35050 13143 35053
rect 15745 35050 15811 35053
rect 13077 35048 15811 35050
rect 13077 34992 13082 35048
rect 13138 34992 15750 35048
rect 15806 34992 15811 35048
rect 13077 34990 15811 34992
rect 13077 34987 13143 34990
rect 15745 34987 15811 34990
rect 10685 34914 10751 34917
rect 13721 34914 13787 34917
rect 10685 34912 13787 34914
rect 10685 34856 10690 34912
rect 10746 34856 13726 34912
rect 13782 34856 13787 34912
rect 10685 34854 13787 34856
rect 10685 34851 10751 34854
rect 13721 34851 13787 34854
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 10869 34778 10935 34781
rect 13353 34778 13419 34781
rect 10869 34776 13419 34778
rect 10869 34720 10874 34776
rect 10930 34720 13358 34776
rect 13414 34720 13419 34776
rect 10869 34718 13419 34720
rect 10869 34715 10935 34718
rect 13353 34715 13419 34718
rect 565 34642 631 34645
rect 2865 34642 2931 34645
rect 565 34640 2931 34642
rect 565 34584 570 34640
rect 626 34584 2870 34640
rect 2926 34584 2931 34640
rect 565 34582 2931 34584
rect 565 34579 631 34582
rect 2865 34579 2931 34582
rect 7097 34642 7163 34645
rect 9397 34642 9463 34645
rect 7097 34640 9463 34642
rect 7097 34584 7102 34640
rect 7158 34584 9402 34640
rect 9458 34584 9463 34640
rect 7097 34582 9463 34584
rect 7097 34579 7163 34582
rect 9397 34579 9463 34582
rect 9581 34642 9647 34645
rect 11421 34642 11487 34645
rect 9581 34640 11487 34642
rect 9581 34584 9586 34640
rect 9642 34584 11426 34640
rect 11482 34584 11487 34640
rect 9581 34582 11487 34584
rect 9581 34579 9647 34582
rect 11421 34579 11487 34582
rect 13445 34642 13511 34645
rect 15377 34642 15443 34645
rect 13445 34640 15443 34642
rect 13445 34584 13450 34640
rect 13506 34584 15382 34640
rect 15438 34584 15443 34640
rect 13445 34582 15443 34584
rect 13445 34579 13511 34582
rect 15377 34579 15443 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3969 34098 4035 34101
rect 9857 34098 9923 34101
rect 3969 34096 9923 34098
rect 3969 34040 3974 34096
rect 4030 34040 9862 34096
rect 9918 34040 9923 34096
rect 3969 34038 9923 34040
rect 3969 34035 4035 34038
rect 9857 34035 9923 34038
rect 3969 33962 4035 33965
rect 10593 33962 10659 33965
rect 3969 33960 10659 33962
rect 3969 33904 3974 33960
rect 4030 33904 10598 33960
rect 10654 33904 10659 33960
rect 3969 33902 10659 33904
rect 3969 33899 4035 33902
rect 10593 33899 10659 33902
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 7649 33554 7715 33557
rect 12525 33554 12591 33557
rect 7649 33552 12591 33554
rect 7649 33496 7654 33552
rect 7710 33496 12530 33552
rect 12586 33496 12591 33552
rect 7649 33494 12591 33496
rect 7649 33491 7715 33494
rect 12525 33491 12591 33494
rect 0 33418 480 33448
rect 1577 33418 1643 33421
rect 0 33416 1643 33418
rect 0 33360 1582 33416
rect 1638 33360 1643 33416
rect 0 33358 1643 33360
rect 0 33328 480 33358
rect 1577 33355 1643 33358
rect 10685 33418 10751 33421
rect 12985 33418 13051 33421
rect 10685 33416 13051 33418
rect 10685 33360 10690 33416
rect 10746 33360 12990 33416
rect 13046 33360 13051 33416
rect 10685 33358 13051 33360
rect 10685 33355 10751 33358
rect 12985 33355 13051 33358
rect 7557 33282 7623 33285
rect 10133 33282 10199 33285
rect 7557 33280 10199 33282
rect 7557 33224 7562 33280
rect 7618 33224 10138 33280
rect 10194 33224 10199 33280
rect 7557 33222 10199 33224
rect 7557 33219 7623 33222
rect 10133 33219 10199 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 7465 32874 7531 32877
rect 11329 32874 11395 32877
rect 7465 32872 11395 32874
rect 7465 32816 7470 32872
rect 7526 32816 11334 32872
rect 11390 32816 11395 32872
rect 7465 32814 11395 32816
rect 7465 32811 7531 32814
rect 11329 32811 11395 32814
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 5717 32602 5783 32605
rect 5717 32600 8770 32602
rect 5717 32544 5722 32600
rect 5778 32544 8770 32600
rect 5717 32542 8770 32544
rect 5717 32539 5783 32542
rect 6637 32466 6703 32469
rect 8017 32466 8083 32469
rect 6637 32464 8083 32466
rect 6637 32408 6642 32464
rect 6698 32408 8022 32464
rect 8078 32408 8083 32464
rect 6637 32406 8083 32408
rect 8710 32466 8770 32542
rect 10777 32466 10843 32469
rect 8710 32464 10843 32466
rect 8710 32408 10782 32464
rect 10838 32408 10843 32464
rect 8710 32406 10843 32408
rect 6637 32403 6703 32406
rect 8017 32403 8083 32406
rect 10777 32403 10843 32406
rect 7373 32330 7439 32333
rect 12525 32330 12591 32333
rect 7373 32328 12591 32330
rect 7373 32272 7378 32328
rect 7434 32272 12530 32328
rect 12586 32272 12591 32328
rect 7373 32270 12591 32272
rect 7373 32267 7439 32270
rect 12525 32267 12591 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 933 31514 999 31517
rect 2865 31514 2931 31517
rect 933 31512 2931 31514
rect 933 31456 938 31512
rect 994 31456 2870 31512
rect 2926 31456 2931 31512
rect 933 31454 2931 31456
rect 933 31451 999 31454
rect 2865 31451 2931 31454
rect 4981 31378 5047 31381
rect 9673 31378 9739 31381
rect 4981 31376 9739 31378
rect 4981 31320 4986 31376
rect 5042 31320 9678 31376
rect 9734 31320 9739 31376
rect 4981 31318 9739 31320
rect 4981 31315 5047 31318
rect 9673 31315 9739 31318
rect 10317 31378 10383 31381
rect 10961 31378 11027 31381
rect 10317 31376 11027 31378
rect 10317 31320 10322 31376
rect 10378 31320 10966 31376
rect 11022 31320 11027 31376
rect 10317 31318 11027 31320
rect 10317 31315 10383 31318
rect 10961 31315 11027 31318
rect 8201 31242 8267 31245
rect 12525 31242 12591 31245
rect 8201 31240 12591 31242
rect 8201 31184 8206 31240
rect 8262 31184 12530 31240
rect 12586 31184 12591 31240
rect 8201 31182 12591 31184
rect 8201 31179 8267 31182
rect 12525 31179 12591 31182
rect 7373 31106 7439 31109
rect 9305 31106 9371 31109
rect 7373 31104 9371 31106
rect 7373 31048 7378 31104
rect 7434 31048 9310 31104
rect 9366 31048 9371 31104
rect 7373 31046 9371 31048
rect 7373 31043 7439 31046
rect 9305 31043 9371 31046
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 4061 30834 4127 30837
rect 10317 30834 10383 30837
rect 4061 30832 10383 30834
rect 4061 30776 4066 30832
rect 4122 30776 10322 30832
rect 10378 30776 10383 30832
rect 4061 30774 10383 30776
rect 4061 30771 4127 30774
rect 10317 30771 10383 30774
rect 5349 30698 5415 30701
rect 10041 30698 10107 30701
rect 5349 30696 10107 30698
rect 5349 30640 5354 30696
rect 5410 30640 10046 30696
rect 10102 30640 10107 30696
rect 5349 30638 10107 30640
rect 5349 30635 5415 30638
rect 10041 30635 10107 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6177 30154 6243 30157
rect 11329 30154 11395 30157
rect 6177 30152 11395 30154
rect 6177 30096 6182 30152
rect 6238 30096 11334 30152
rect 11390 30096 11395 30152
rect 6177 30094 11395 30096
rect 6177 30091 6243 30094
rect 11329 30091 11395 30094
rect 12249 30018 12315 30021
rect 15520 30018 16000 30048
rect 12249 30016 16000 30018
rect 12249 29960 12254 30016
rect 12310 29960 16000 30016
rect 12249 29958 16000 29960
rect 12249 29955 12315 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 5441 29610 5507 29613
rect 9673 29610 9739 29613
rect 5441 29608 9739 29610
rect 5441 29552 5446 29608
rect 5502 29552 9678 29608
rect 9734 29552 9739 29608
rect 5441 29550 9739 29552
rect 5441 29547 5507 29550
rect 9673 29547 9739 29550
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 5165 28522 5231 28525
rect 10041 28522 10107 28525
rect 5165 28520 10107 28522
rect 5165 28464 5170 28520
rect 5226 28464 10046 28520
rect 10102 28464 10107 28520
rect 5165 28462 10107 28464
rect 5165 28459 5231 28462
rect 10041 28459 10107 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 6821 27434 6887 27437
rect 15009 27434 15075 27437
rect 6821 27432 15075 27434
rect 6821 27376 6826 27432
rect 6882 27376 15014 27432
rect 15070 27376 15075 27432
rect 6821 27374 15075 27376
rect 6821 27371 6887 27374
rect 15009 27371 15075 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6177 25938 6243 25941
rect 11329 25938 11395 25941
rect 6177 25936 11395 25938
rect 6177 25880 6182 25936
rect 6238 25880 11334 25936
rect 11390 25880 11395 25936
rect 6177 25878 11395 25880
rect 6177 25875 6243 25878
rect 11329 25875 11395 25878
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 9949 24986 10015 24989
rect 12433 24986 12499 24989
rect 9949 24984 12499 24986
rect 9949 24928 9954 24984
rect 10010 24928 12438 24984
rect 12494 24928 12499 24984
rect 9949 24926 12499 24928
rect 9949 24923 10015 24926
rect 12433 24923 12499 24926
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 5717 24170 5783 24173
rect 10501 24170 10567 24173
rect 5717 24168 10567 24170
rect 5717 24112 5722 24168
rect 5778 24112 10506 24168
rect 10562 24112 10567 24168
rect 5717 24110 10567 24112
rect 5717 24107 5783 24110
rect 10501 24107 10567 24110
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 10961 23626 11027 23629
rect 12525 23626 12591 23629
rect 10961 23624 12591 23626
rect 10961 23568 10966 23624
rect 11022 23568 12530 23624
rect 12586 23568 12591 23624
rect 10961 23566 12591 23568
rect 10961 23563 11027 23566
rect 12525 23563 12591 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 4153 22674 4219 22677
rect 9673 22674 9739 22677
rect 4153 22672 9739 22674
rect 4153 22616 4158 22672
rect 4214 22616 9678 22672
rect 9734 22616 9739 22672
rect 4153 22614 9739 22616
rect 4153 22611 4219 22614
rect 9673 22611 9739 22614
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 4705 22130 4771 22133
rect 6085 22130 6151 22133
rect 4705 22128 6151 22130
rect 4705 22072 4710 22128
rect 4766 22072 6090 22128
rect 6146 22072 6151 22128
rect 4705 22070 6151 22072
rect 4705 22067 4771 22070
rect 6085 22067 6151 22070
rect 10869 22130 10935 22133
rect 12709 22130 12775 22133
rect 10869 22128 12775 22130
rect 10869 22072 10874 22128
rect 10930 22072 12714 22128
rect 12770 22072 12775 22128
rect 10869 22070 12775 22072
rect 10869 22067 10935 22070
rect 12709 22067 12775 22070
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3417 21042 3483 21045
rect 7741 21042 7807 21045
rect 3417 21040 7807 21042
rect 3417 20984 3422 21040
rect 3478 20984 7746 21040
rect 7802 20984 7807 21040
rect 3417 20982 7807 20984
rect 3417 20979 3483 20982
rect 7741 20979 7807 20982
rect 7833 20906 7899 20909
rect 10317 20906 10383 20909
rect 7833 20904 10383 20906
rect 7833 20848 7838 20904
rect 7894 20848 10322 20904
rect 10378 20848 10383 20904
rect 7833 20846 10383 20848
rect 7833 20843 7899 20846
rect 10317 20843 10383 20846
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 8109 20226 8175 20229
rect 9857 20226 9923 20229
rect 8109 20224 9923 20226
rect 8109 20168 8114 20224
rect 8170 20168 9862 20224
rect 9918 20168 9923 20224
rect 8109 20166 9923 20168
rect 8109 20163 8175 20166
rect 9857 20163 9923 20166
rect 6277 20160 6597 20161
rect 0 20090 480 20120
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 2957 20090 3023 20093
rect 3509 20090 3575 20093
rect 0 20088 3575 20090
rect 0 20032 2962 20088
rect 3018 20032 3514 20088
rect 3570 20032 3575 20088
rect 0 20030 3575 20032
rect 0 20000 480 20030
rect 2957 20027 3023 20030
rect 3509 20027 3575 20030
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 3877 19410 3943 19413
rect 8109 19410 8175 19413
rect 3877 19408 8175 19410
rect 3877 19352 3882 19408
rect 3938 19352 8114 19408
rect 8170 19352 8175 19408
rect 3877 19350 8175 19352
rect 3877 19347 3943 19350
rect 8109 19347 8175 19350
rect 9949 19410 10015 19413
rect 12065 19410 12131 19413
rect 9949 19408 12131 19410
rect 9949 19352 9954 19408
rect 10010 19352 12070 19408
rect 12126 19352 12131 19408
rect 9949 19350 12131 19352
rect 9949 19347 10015 19350
rect 12065 19347 12131 19350
rect 3049 19274 3115 19277
rect 5625 19274 5691 19277
rect 3049 19272 5691 19274
rect 3049 19216 3054 19272
rect 3110 19216 5630 19272
rect 5686 19216 5691 19272
rect 3049 19214 5691 19216
rect 3049 19211 3115 19214
rect 5625 19211 5691 19214
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3233 18866 3299 18869
rect 6729 18866 6795 18869
rect 3233 18864 6795 18866
rect 3233 18808 3238 18864
rect 3294 18808 6734 18864
rect 6790 18808 6795 18864
rect 3233 18806 6795 18808
rect 3233 18803 3299 18806
rect 6729 18803 6795 18806
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 3417 18050 3483 18053
rect 6085 18050 6151 18053
rect 3417 18048 6151 18050
rect 3417 17992 3422 18048
rect 3478 17992 6090 18048
rect 6146 17992 6151 18048
rect 3417 17990 6151 17992
rect 3417 17987 3483 17990
rect 6085 17987 6151 17990
rect 6729 18050 6795 18053
rect 8477 18050 8543 18053
rect 6729 18048 8543 18050
rect 6729 17992 6734 18048
rect 6790 17992 8482 18048
rect 8538 17992 8543 18048
rect 6729 17990 8543 17992
rect 6729 17987 6795 17990
rect 8477 17987 8543 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 5073 17778 5139 17781
rect 7281 17778 7347 17781
rect 5073 17776 7347 17778
rect 5073 17720 5078 17776
rect 5134 17720 7286 17776
rect 7342 17720 7347 17776
rect 5073 17718 7347 17720
rect 5073 17715 5139 17718
rect 7281 17715 7347 17718
rect 7925 17778 7991 17781
rect 13997 17778 14063 17781
rect 7925 17776 14063 17778
rect 7925 17720 7930 17776
rect 7986 17720 14002 17776
rect 14058 17720 14063 17776
rect 7925 17718 14063 17720
rect 7925 17715 7991 17718
rect 13997 17715 14063 17718
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3509 17234 3575 17237
rect 8845 17234 8911 17237
rect 3509 17232 8911 17234
rect 3509 17176 3514 17232
rect 3570 17176 8850 17232
rect 8906 17176 8911 17232
rect 3509 17174 8911 17176
rect 3509 17171 3575 17174
rect 8845 17171 8911 17174
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3233 16554 3299 16557
rect 7373 16554 7439 16557
rect 3233 16552 7439 16554
rect 3233 16496 3238 16552
rect 3294 16496 7378 16552
rect 7434 16496 7439 16552
rect 3233 16494 7439 16496
rect 3233 16491 3299 16494
rect 7373 16491 7439 16494
rect 9305 16554 9371 16557
rect 11237 16554 11303 16557
rect 9305 16552 11303 16554
rect 9305 16496 9310 16552
rect 9366 16496 11242 16552
rect 11298 16496 11303 16552
rect 9305 16494 11303 16496
rect 9305 16491 9371 16494
rect 11237 16491 11303 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 5533 11250 5599 11253
rect 8017 11250 8083 11253
rect 12157 11250 12223 11253
rect 5533 11248 12223 11250
rect 5533 11192 5538 11248
rect 5594 11192 8022 11248
rect 8078 11192 12162 11248
rect 12218 11192 12223 11248
rect 5533 11190 12223 11192
rect 5533 11187 5599 11190
rect 8017 11187 8083 11190
rect 12157 11187 12223 11190
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 4337 10570 4403 10573
rect 7097 10570 7163 10573
rect 10685 10570 10751 10573
rect 4337 10568 6746 10570
rect 4337 10512 4342 10568
rect 4398 10512 6746 10568
rect 4337 10510 6746 10512
rect 4337 10507 4403 10510
rect 6686 10437 6746 10510
rect 7097 10568 10751 10570
rect 7097 10512 7102 10568
rect 7158 10512 10690 10568
rect 10746 10512 10751 10568
rect 7097 10510 10751 10512
rect 7097 10507 7163 10510
rect 10685 10507 10751 10510
rect 6686 10434 6795 10437
rect 7281 10434 7347 10437
rect 9765 10434 9831 10437
rect 6686 10432 9831 10434
rect 6686 10376 6734 10432
rect 6790 10376 7286 10432
rect 7342 10376 9770 10432
rect 9826 10376 9831 10432
rect 6686 10374 9831 10376
rect 6729 10371 6795 10374
rect 7281 10371 7347 10374
rect 9765 10371 9831 10374
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 1669 10298 1735 10301
rect 5625 10298 5691 10301
rect 1669 10296 5691 10298
rect 1669 10240 1674 10296
rect 1730 10240 5630 10296
rect 5686 10240 5691 10296
rect 1669 10238 5691 10240
rect 1669 10235 1735 10238
rect 5625 10235 5691 10238
rect 1393 10026 1459 10029
rect 5993 10026 6059 10029
rect 7465 10026 7531 10029
rect 1393 10024 7531 10026
rect 1393 9968 1398 10024
rect 1454 9968 5998 10024
rect 6054 9968 7470 10024
rect 7526 9968 7531 10024
rect 1393 9966 7531 9968
rect 1393 9963 1459 9966
rect 5993 9963 6059 9966
rect 7465 9963 7531 9966
rect 7833 10026 7899 10029
rect 10041 10026 10107 10029
rect 10225 10026 10291 10029
rect 15520 10026 16000 10056
rect 7833 10024 10107 10026
rect 7833 9968 7838 10024
rect 7894 9968 10046 10024
rect 10102 9968 10107 10024
rect 7833 9966 10107 9968
rect 7833 9963 7899 9966
rect 10041 9963 10107 9966
rect 10182 10024 16000 10026
rect 10182 9968 10230 10024
rect 10286 9968 16000 10024
rect 10182 9966 16000 9968
rect 10182 9963 10291 9966
rect 9489 9890 9555 9893
rect 10182 9890 10242 9963
rect 15520 9936 16000 9966
rect 9489 9888 10242 9890
rect 9489 9832 9494 9888
rect 9550 9832 10242 9888
rect 9489 9830 10242 9832
rect 9489 9827 9555 9830
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 5901 7850 5967 7853
rect 12525 7850 12591 7853
rect 5901 7848 12591 7850
rect 5901 7792 5906 7848
rect 5962 7792 12530 7848
rect 12586 7792 12591 7848
rect 5901 7790 12591 7792
rect 5901 7787 5967 7790
rect 12525 7787 12591 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 0 6762 480 6792
rect 4153 6762 4219 6765
rect 0 6760 4219 6762
rect 0 6704 4158 6760
rect 4214 6704 4219 6760
rect 0 6702 4219 6704
rect 0 6672 480 6702
rect 4153 6699 4219 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3325 5674 3391 5677
rect 7649 5674 7715 5677
rect 3325 5672 7715 5674
rect 3325 5616 3330 5672
rect 3386 5616 7654 5672
rect 7710 5616 7715 5672
rect 3325 5614 7715 5616
rect 3325 5611 3391 5614
rect 7649 5611 7715 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 10593 5130 10659 5133
rect 13813 5130 13879 5133
rect 10593 5128 13879 5130
rect 10593 5072 10598 5128
rect 10654 5072 13818 5128
rect 13874 5072 13879 5128
rect 10593 5070 13879 5072
rect 10593 5067 10659 5070
rect 13813 5067 13879 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 5993 4722 6059 4725
rect 8201 4722 8267 4725
rect 5993 4720 8267 4722
rect 5993 4664 5998 4720
rect 6054 4664 8206 4720
rect 8262 4664 8267 4720
rect 5993 4662 8267 4664
rect 5993 4659 6059 4662
rect 8201 4659 8267 4662
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 2405 4178 2471 4181
rect 4153 4178 4219 4181
rect 2405 4176 4219 4178
rect 2405 4120 2410 4176
rect 2466 4120 4158 4176
rect 4214 4120 4219 4176
rect 2405 4118 4219 4120
rect 2405 4115 2471 4118
rect 4153 4115 4219 4118
rect 7373 4042 7439 4045
rect 8845 4042 8911 4045
rect 7373 4040 8911 4042
rect 7373 3984 7378 4040
rect 7434 3984 8850 4040
rect 8906 3984 8911 4040
rect 7373 3982 8911 3984
rect 7373 3979 7439 3982
rect 8845 3979 8911 3982
rect 10225 4042 10291 4045
rect 14641 4042 14707 4045
rect 10225 4040 14707 4042
rect 10225 3984 10230 4040
rect 10286 3984 14646 4040
rect 14702 3984 14707 4040
rect 10225 3982 14707 3984
rect 10225 3979 10291 3982
rect 14641 3979 14707 3982
rect 12985 3906 13051 3909
rect 15377 3906 15443 3909
rect 12985 3904 15443 3906
rect 12985 3848 12990 3904
rect 13046 3848 15382 3904
rect 15438 3848 15443 3904
rect 12985 3846 15443 3848
rect 12985 3843 13051 3846
rect 15377 3843 15443 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 7741 3634 7807 3637
rect 12801 3634 12867 3637
rect 7741 3632 12867 3634
rect 7741 3576 7746 3632
rect 7802 3576 12806 3632
rect 12862 3576 12867 3632
rect 7741 3574 12867 3576
rect 7741 3571 7807 3574
rect 12801 3571 12867 3574
rect 2589 3498 2655 3501
rect 4245 3498 4311 3501
rect 2589 3496 4311 3498
rect 2589 3440 2594 3496
rect 2650 3440 4250 3496
rect 4306 3440 4311 3496
rect 2589 3438 4311 3440
rect 2589 3435 2655 3438
rect 4245 3435 4311 3438
rect 7925 3498 7991 3501
rect 10593 3498 10659 3501
rect 7925 3496 10659 3498
rect 7925 3440 7930 3496
rect 7986 3440 10598 3496
rect 10654 3440 10659 3496
rect 7925 3438 10659 3440
rect 7925 3435 7991 3438
rect 10593 3435 10659 3438
rect 11973 3498 12039 3501
rect 14181 3498 14247 3501
rect 11973 3496 14247 3498
rect 11973 3440 11978 3496
rect 12034 3440 14186 3496
rect 14242 3440 14247 3496
rect 11973 3438 14247 3440
rect 11973 3435 12039 3438
rect 14181 3435 14247 3438
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 1485 3090 1551 3093
rect 4245 3090 4311 3093
rect 1485 3088 4311 3090
rect 1485 3032 1490 3088
rect 1546 3032 4250 3088
rect 4306 3032 4311 3088
rect 1485 3030 4311 3032
rect 1485 3027 1551 3030
rect 4245 3027 4311 3030
rect 4613 3090 4679 3093
rect 10593 3090 10659 3093
rect 4613 3088 10659 3090
rect 4613 3032 4618 3088
rect 4674 3032 10598 3088
rect 10654 3032 10659 3088
rect 4613 3030 10659 3032
rect 4613 3027 4679 3030
rect 10593 3027 10659 3030
rect 933 2954 999 2957
rect 2865 2954 2931 2957
rect 933 2952 2931 2954
rect 933 2896 938 2952
rect 994 2896 2870 2952
rect 2926 2896 2931 2952
rect 933 2894 2931 2896
rect 933 2891 999 2894
rect 2865 2891 2931 2894
rect 4337 2954 4403 2957
rect 7465 2954 7531 2957
rect 4337 2952 7531 2954
rect 4337 2896 4342 2952
rect 4398 2896 7470 2952
rect 7526 2896 7531 2952
rect 4337 2894 7531 2896
rect 4337 2891 4403 2894
rect 7465 2891 7531 2894
rect 7649 2954 7715 2957
rect 13629 2954 13695 2957
rect 7649 2952 13695 2954
rect 7649 2896 7654 2952
rect 7710 2896 13634 2952
rect 13690 2896 13695 2952
rect 7649 2894 13695 2896
rect 7649 2891 7715 2894
rect 13629 2891 13695 2894
rect 565 2818 631 2821
rect 3049 2818 3115 2821
rect 565 2816 3115 2818
rect 565 2760 570 2816
rect 626 2760 3054 2816
rect 3110 2760 3115 2816
rect 565 2758 3115 2760
rect 565 2755 631 2758
rect 3049 2755 3115 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 4705 2546 4771 2549
rect 7189 2546 7255 2549
rect 4705 2544 7255 2546
rect 4705 2488 4710 2544
rect 4766 2488 7194 2544
rect 7250 2488 7255 2544
rect 4705 2486 7255 2488
rect 4705 2483 4771 2486
rect 7189 2483 7255 2486
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 197 1458 263 1461
rect 1577 1458 1643 1461
rect 197 1456 1643 1458
rect 197 1400 202 1456
rect 258 1400 1582 1456
rect 1638 1400 1643 1456
rect 197 1398 1643 1400
rect 197 1395 263 1398
rect 1577 1395 1643 1398
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_fill_2  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _40_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 774 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _14_
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_48
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_40
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_52
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_60
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _24_
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_87
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _29_
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_48
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_78
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_96
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _02_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_3_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_12  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_140
timestamp 1586364061
transform 1 0 13984 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_63
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_109
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_21
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_24
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_49
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_48
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_69
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_73
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_50
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_54
timestamp 1586364061
transform 1 0 6072 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_100
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_120
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_75
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_79
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9752 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_113
timestamp 1586364061
transform 1 0 11500 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_125
timestamp 1586364061
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_38
timestamp 1586364061
transform 1 0 4600 0 -1 21216
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_61
timestamp 1586364061
transform 1 0 6716 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_33
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_45
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_38
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_62
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_74
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_86
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_21
timestamp 1586364061
transform 1 0 3036 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_24
timestamp 1586364061
transform 1 0 3312 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_19
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3128 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_31
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_43
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_41_55
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12052 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_121
timestamp 1586364061
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_21
timestamp 1586364061
transform 1 0 3036 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_24
timestamp 1586364061
transform 1 0 3312 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_30
timestamp 1586364061
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_buf_1  mux_left_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12052 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_122
timestamp 1586364061
transform 1 0 12328 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4876 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5244 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_43
timestamp 1586364061
transform 1 0 5060 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_47
timestamp 1586364061
transform 1 0 5428 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_8  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4876 0 -1 26656
box -38 -48 866 592
use scs8hd_fill_1  FILLER_44_40
timestamp 1586364061
transform 1 0 4784 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_50
timestamp 1586364061
transform 1 0 5704 0 -1 26656
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6808 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_64
timestamp 1586364061
transform 1 0 6992 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_buf_1  mux_right_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_6
timestamp 1586364061
transform 1 0 1656 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_10
timestamp 1586364061
transform 1 0 2024 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_22
timestamp 1586364061
transform 1 0 3128 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_34
timestamp 1586364061
transform 1 0 4232 0 1 26656
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_46
timestamp 1586364061
transform 1 0 5336 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_50
timestamp 1586364061
transform 1 0 5704 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_53
timestamp 1586364061
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_71
timestamp 1586364061
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_75
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_87
timestamp 1586364061
transform 1 0 9108 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_99
timestamp 1586364061
transform 1 0 10212 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_111
timestamp 1586364061
transform 1 0 11316 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_45_119
timestamp 1586364061
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6532 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_conb_1  _03_
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_65
timestamp 1586364061
transform 1 0 7084 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_77
timestamp 1586364061
transform 1 0 8188 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_89
timestamp 1586364061
transform 1 0 9292 0 1 27744
box -38 -48 774 592
use scs8hd_fill_1  FILLER_47_97
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 130 592
use scs8hd_buf_2  _26_
timestamp 1586364061
transform 1 0 10304 0 1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 10856 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_104
timestamp 1586364061
transform 1 0 10672 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_108
timestamp 1586364061
transform 1 0 11040 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_120
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_48_99
timestamp 1586364061
transform 1 0 10212 0 -1 28832
box -38 -48 130 592
use scs8hd_buf_2  _06_
timestamp 1586364061
transform 1 0 10304 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_104
timestamp 1586364061
transform 1 0 10672 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_116
timestamp 1586364061
transform 1 0 11776 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_128
timestamp 1586364061
transform 1 0 12880 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_48_140
timestamp 1586364061
transform 1 0 13984 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_106
timestamp 1586364061
transform 1 0 10856 0 1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_49_111
timestamp 1586364061
transform 1 0 11316 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  FILLER_49_119
timestamp 1586364061
transform 1 0 12052 0 1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_buf_2  _25_
timestamp 1586364061
transform 1 0 11132 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_4  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_113
timestamp 1586364061
transform 1 0 11500 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_125
timestamp 1586364061
transform 1 0 12604 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_137
timestamp 1586364061
transform 1 0 13708 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 4048 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_31
timestamp 1586364061
transform 1 0 3956 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_34
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_46
timestamp 1586364061
transform 1 0 5336 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_51_58
timestamp 1586364061
transform 1 0 6440 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_buf_2  _27_
timestamp 1586364061
transform 1 0 9844 0 1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_51_92
timestamp 1586364061
transform 1 0 9568 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_99
timestamp 1586364061
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use scs8hd_buf_2  _05_
timestamp 1586364061
transform 1 0 11132 0 1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 11684 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_103
timestamp 1586364061
transform 1 0 10580 0 1 29920
box -38 -48 590 592
use scs8hd_fill_2  FILLER_51_113
timestamp 1586364061
transform 1 0 11500 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_117
timestamp 1586364061
transform 1 0 11868 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_121
timestamp 1586364061
transform 1 0 12236 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_53_8
timestamp 1586364061
transform 1 0 1840 0 1 31008
box -38 -48 590 592
use scs8hd_decap_3  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 1656 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_53_14
timestamp 1586364061
transform 1 0 2392 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 222 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 2668 0 1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_25
timestamp 1586364061
transform 1 0 3404 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_21
timestamp 1586364061
transform 1 0 3036 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 3220 0 1 31008
box -38 -48 222 592
use scs8hd_buf_2  _15_
timestamp 1586364061
transform 1 0 3772 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_37
timestamp 1586364061
transform 1 0 4508 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_33
timestamp 1586364061
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_36
timestamp 1586364061
transform 1 0 4416 0 -1 31008
box -38 -48 1142 592
use scs8hd_buf_2  _09_
timestamp 1586364061
transform 1 0 4876 0 1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 6440 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_48
timestamp 1586364061
transform 1 0 5520 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_45
timestamp 1586364061
transform 1 0 5244 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_53_49
timestamp 1586364061
transform 1 0 5612 0 1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_53_57
timestamp 1586364061
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_66
timestamp 1586364061
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_60
timestamp 1586364061
transform 1 0 6624 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_buf_2  _12_
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_53_70
timestamp 1586364061
transform 1 0 7544 0 1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_75
timestamp 1586364061
transform 1 0 8004 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_72
timestamp 1586364061
transform 1 0 7728 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_60
timestamp 1586364061
transform 1 0 6624 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_53_87
timestamp 1586364061
transform 1 0 9108 0 1 31008
box -38 -48 406 592
use scs8hd_decap_8  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_53_99
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_buf_2  _08_
timestamp 1586364061
transform 1 0 9476 0 1 31008
box -38 -48 406 592
use scs8hd_buf_2  _07_
timestamp 1586364061
transform 1 0 9844 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_99
timestamp 1586364061
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_111
timestamp 1586364061
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_103
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_53_115
timestamp 1586364061
transform 1 0 11684 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_119
timestamp 1586364061
transform 1 0 12052 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_127
timestamp 1586364061
transform 1 0 12788 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use scs8hd_decap_8  FILLER_53_136
timestamp 1586364061
transform 1 0 13616 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  FILLER_53_131
timestamp 1586364061
transform 1 0 13156 0 1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_52_135
timestamp 1586364061
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 13432 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 12972 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_123
timestamp 1586364061
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_143
timestamp 1586364061
transform 1 0 14260 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_144
timestamp 1586364061
transform 1 0 14352 0 1 31008
box -38 -48 222 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 2760 0 -1 32096
box -38 -48 406 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 1656 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_8  FILLER_54_10
timestamp 1586364061
transform 1 0 2024 0 -1 32096
box -38 -48 774 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_22
timestamp 1586364061
transform 1 0 3128 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_30
timestamp 1586364061
transform 1 0 3864 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_36
timestamp 1586364061
transform 1 0 4416 0 -1 32096
box -38 -48 774 592
use scs8hd_buf_2  _10_
timestamp 1586364061
transform 1 0 5336 0 -1 32096
box -38 -48 406 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 6440 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_50
timestamp 1586364061
transform 1 0 5704 0 -1 32096
box -38 -48 774 592
use scs8hd_buf_2  _04_
timestamp 1586364061
transform 1 0 7820 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_8  FILLER_54_62
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_54_70
timestamp 1586364061
transform 1 0 7544 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_77
timestamp 1586364061
transform 1 0 8188 0 -1 32096
box -38 -48 1142 592
use scs8hd_buf_2  _11_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_89
timestamp 1586364061
transform 1 0 9292 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_97
timestamp 1586364061
transform 1 0 10028 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_109
timestamp 1586364061
transform 1 0 11132 0 -1 32096
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 13432 0 -1 32096
box -38 -48 406 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 12328 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_121
timestamp 1586364061
transform 1 0 12236 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_126
timestamp 1586364061
transform 1 0 12696 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_8  FILLER_54_138
timestamp 1586364061
transform 1 0 13800 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 590 592
use scs8hd_buf_2  _13_
timestamp 1586364061
transform 1 0 4140 0 1 32096
box -38 -48 406 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 3036 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_25
timestamp 1586364061
transform 1 0 3404 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_29
timestamp 1586364061
transform 1 0 3772 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_37
timestamp 1586364061
transform 1 0 4508 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_41
timestamp 1586364061
transform 1 0 4876 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 774 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 7360 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_66
timestamp 1586364061
transform 1 0 7176 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_70
timestamp 1586364061
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use scs8hd_buf_2  _28_
timestamp 1586364061
transform 1 0 10028 0 1 32096
box -38 -48 406 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 8924 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 9476 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_82
timestamp 1586364061
transform 1 0 8648 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_89
timestamp 1586364061
transform 1 0 9292 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_93
timestamp 1586364061
transform 1 0 9660 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 10580 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_101
timestamp 1586364061
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_105
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 406 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_121
timestamp 1586364061
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_127
timestamp 1586364061
transform 1 0 12788 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_131
timestamp 1586364061
transform 1 0 13156 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 6672 480 6792 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 20000 480 20120 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 33328 480 33448 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 prog_clk
port 83 nsew default input
rlabel metal3 s 15520 29928 16000 30048 6 right_grid_pin_52_
port 84 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 85 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 86 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
