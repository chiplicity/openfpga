magic
tech EFS8A
magscale 1 2
timestamp 1602269619
<< locali >>
rect 2639 11169 2766 11203
rect 5583 11169 5618 11203
rect 6595 11169 6630 11203
rect 8251 11169 8286 11203
rect 7935 6953 7941 6987
rect 7935 6885 7969 6953
rect 13679 6817 13714 6851
rect 2697 6239 2731 6409
rect 6377 6239 6411 6409
rect 4111 4641 4238 4675
rect 4905 4471 4939 4573
rect 8309 4539 8343 4709
rect 4445 4131 4479 4165
rect 4353 4097 4479 4131
rect 8125 3383 8159 3621
rect 15243 3553 15370 3587
rect 9873 2975 9907 3077
rect 14105 2907 14139 3145
rect 3709 2295 3743 2465
rect 6561 2295 6595 2533
<< viali >>
rect 6193 18377 6227 18411
rect 7389 18377 7423 18411
rect 13001 18377 13035 18411
rect 5641 18173 5675 18207
rect 7205 18173 7239 18207
rect 12817 18173 12851 18207
rect 13369 18173 13403 18207
rect 5825 18037 5859 18071
rect 7849 18037 7883 18071
rect 4813 17833 4847 17867
rect 4629 17697 4663 17731
rect 19257 17289 19291 17323
rect 19073 17085 19107 17119
rect 19625 17085 19659 17119
rect 4629 16949 4663 16983
rect 19073 14433 19107 14467
rect 19257 14229 19291 14263
rect 19073 14025 19107 14059
rect 1593 11781 1627 11815
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 8100 11645 8134 11679
rect 8171 11509 8205 11543
rect 8585 11509 8619 11543
rect 7113 11305 7147 11339
rect 12633 11305 12667 11339
rect 2605 11169 2639 11203
rect 5549 11169 5583 11203
rect 6561 11169 6595 11203
rect 8217 11169 8251 11203
rect 12449 11169 12483 11203
rect 2835 10965 2869 10999
rect 3801 10965 3835 10999
rect 5687 10965 5721 10999
rect 6699 10965 6733 10999
rect 8355 10965 8389 10999
rect 1593 10761 1627 10795
rect 3341 10761 3375 10795
rect 6285 10761 6319 10795
rect 6653 10761 6687 10795
rect 12633 10761 12667 10795
rect 3801 10625 3835 10659
rect 4721 10625 4755 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 1409 10557 1443 10591
rect 1961 10557 1995 10591
rect 2548 10557 2582 10591
rect 2973 10557 3007 10591
rect 5784 10557 5818 10591
rect 8436 10557 8470 10591
rect 8861 10557 8895 10591
rect 3893 10489 3927 10523
rect 4445 10489 4479 10523
rect 5871 10489 5905 10523
rect 7021 10489 7055 10523
rect 8539 10489 8573 10523
rect 2651 10421 2685 10455
rect 5641 10421 5675 10455
rect 8309 10421 8343 10455
rect 10333 10421 10367 10455
rect 7297 10217 7331 10251
rect 10793 10217 10827 10251
rect 15485 10217 15519 10251
rect 3893 10149 3927 10183
rect 4261 10149 4295 10183
rect 4813 10149 4847 10183
rect 5089 10149 5123 10183
rect 6009 10149 6043 10183
rect 6101 10149 6135 10183
rect 7021 10149 7055 10183
rect 7573 10149 7607 10183
rect 7665 10149 7699 10183
rect 12403 10149 12437 10183
rect 2513 10081 2547 10115
rect 10241 10081 10275 10115
rect 11320 10081 11354 10115
rect 12316 10081 12350 10115
rect 15301 10081 15335 10115
rect 2605 10013 2639 10047
rect 2973 10013 3007 10047
rect 4169 10013 4203 10047
rect 6653 10013 6687 10047
rect 7941 10013 7975 10047
rect 9689 10013 9723 10047
rect 1777 9877 1811 9911
rect 3249 9877 3283 9911
rect 11391 9877 11425 9911
rect 2697 9673 2731 9707
rect 5917 9673 5951 9707
rect 6285 9673 6319 9707
rect 8217 9673 8251 9707
rect 10241 9673 10275 9707
rect 4169 9605 4203 9639
rect 6929 9537 6963 9571
rect 7205 9537 7239 9571
rect 9321 9537 9355 9571
rect 10885 9537 10919 9571
rect 11161 9537 11195 9571
rect 12633 9537 12667 9571
rect 1777 9469 1811 9503
rect 3249 9469 3283 9503
rect 4537 9469 4571 9503
rect 4997 9469 5031 9503
rect 3611 9401 3645 9435
rect 5318 9401 5352 9435
rect 6653 9401 6687 9435
rect 7021 9401 7055 9435
rect 9413 9401 9447 9435
rect 9965 9401 9999 9435
rect 10701 9401 10735 9435
rect 10977 9401 11011 9435
rect 1961 9333 1995 9367
rect 3065 9333 3099 9367
rect 4813 9333 4847 9367
rect 7849 9333 7883 9367
rect 9137 9333 9171 9367
rect 11805 9333 11839 9367
rect 15393 9333 15427 9367
rect 1685 9129 1719 9163
rect 3157 9129 3191 9163
rect 4537 9129 4571 9163
rect 6009 9129 6043 9163
rect 6469 9129 6503 9163
rect 9321 9129 9355 9163
rect 2599 9061 2633 9095
rect 6653 9061 6687 9095
rect 6745 9061 6779 9095
rect 10517 9061 10551 9095
rect 10609 9061 10643 9095
rect 11989 9061 12023 9095
rect 4445 8993 4479 9027
rect 4721 8993 4755 9027
rect 5089 8993 5123 9027
rect 5457 8993 5491 9027
rect 8652 8993 8686 9027
rect 11161 8993 11195 9027
rect 12357 8993 12391 9027
rect 2237 8925 2271 8959
rect 3525 8857 3559 8891
rect 7205 8857 7239 8891
rect 8723 8857 8757 8891
rect 2145 8789 2179 8823
rect 3893 8789 3927 8823
rect 7573 8789 7607 8823
rect 9873 8789 9907 8823
rect 8033 8585 8067 8619
rect 9505 8585 9539 8619
rect 10241 8585 10275 8619
rect 11345 8585 11379 8619
rect 12081 8585 12115 8619
rect 9873 8517 9907 8551
rect 10977 8517 11011 8551
rect 2329 8449 2363 8483
rect 8585 8449 8619 8483
rect 10425 8449 10459 8483
rect 2789 8381 2823 8415
rect 3341 8381 3375 8415
rect 3801 8381 3835 8415
rect 4169 8381 4203 8415
rect 4997 8381 5031 8415
rect 5733 8381 5767 8415
rect 6101 8381 6135 8415
rect 6837 8381 6871 8415
rect 12484 8381 12518 8415
rect 12587 8381 12621 8415
rect 5089 8313 5123 8347
rect 7158 8313 7192 8347
rect 8906 8313 8940 8347
rect 10517 8313 10551 8347
rect 12909 8313 12943 8347
rect 1593 8245 1627 8279
rect 2697 8245 2731 8279
rect 2881 8245 2915 8279
rect 4537 8245 4571 8279
rect 6561 8245 6595 8279
rect 7757 8245 7791 8279
rect 8493 8245 8527 8279
rect 10609 8041 10643 8075
rect 11253 8041 11287 8075
rect 2145 7973 2179 8007
rect 6285 7973 6319 8007
rect 7297 7973 7331 8007
rect 10010 7973 10044 8007
rect 10977 7973 11011 8007
rect 13001 7973 13035 8007
rect 1501 7905 1535 7939
rect 2421 7905 2455 7939
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 5825 7905 5859 7939
rect 6009 7905 6043 7939
rect 8585 7905 8619 7939
rect 11713 7905 11747 7939
rect 11897 7905 11931 7939
rect 3157 7837 3191 7871
rect 6561 7837 6595 7871
rect 7205 7837 7239 7871
rect 8125 7837 8159 7871
rect 9689 7837 9723 7871
rect 11989 7837 12023 7871
rect 7757 7769 7791 7803
rect 2881 7701 2915 7735
rect 3617 7701 3651 7735
rect 4261 7701 4295 7735
rect 4629 7701 4663 7735
rect 6929 7701 6963 7735
rect 8953 7701 8987 7735
rect 9321 7701 9355 7735
rect 2513 7497 2547 7531
rect 4997 7497 5031 7531
rect 7757 7497 7791 7531
rect 9137 7497 9171 7531
rect 10241 7497 10275 7531
rect 12633 7497 12667 7531
rect 6285 7429 6319 7463
rect 12173 7429 12207 7463
rect 5917 7361 5951 7395
rect 10885 7361 10919 7395
rect 11253 7361 11287 7395
rect 1409 7293 1443 7327
rect 2789 7293 2823 7327
rect 3341 7293 3375 7327
rect 3617 7293 3651 7327
rect 3985 7293 4019 7327
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 8033 7293 8067 7327
rect 12449 7293 12483 7327
rect 7158 7225 7192 7259
rect 9321 7225 9355 7259
rect 9413 7225 9447 7259
rect 9965 7225 9999 7259
rect 10701 7225 10735 7259
rect 10977 7225 11011 7259
rect 1593 7157 1627 7191
rect 2237 7157 2271 7191
rect 2973 7157 3007 7191
rect 4629 7157 4663 7191
rect 6653 7157 6687 7191
rect 8769 7157 8803 7191
rect 11897 7157 11931 7191
rect 13093 7157 13127 7191
rect 1685 6953 1719 6987
rect 2053 6953 2087 6987
rect 3433 6953 3467 6987
rect 7389 6953 7423 6987
rect 7941 6953 7975 6987
rect 13783 6953 13817 6987
rect 6745 6885 6779 6919
rect 10701 6885 10735 6919
rect 11253 6885 11287 6919
rect 2973 6817 3007 6851
rect 5273 6817 5307 6851
rect 6009 6817 6043 6851
rect 6101 6817 6135 6851
rect 6469 6817 6503 6851
rect 7021 6817 7055 6851
rect 12081 6817 12115 6851
rect 12357 6817 12391 6851
rect 13645 6817 13679 6851
rect 3065 6749 3099 6783
rect 4261 6749 4295 6783
rect 7573 6749 7607 6783
rect 8769 6749 8803 6783
rect 10609 6749 10643 6783
rect 11897 6749 11931 6783
rect 9873 6681 9907 6715
rect 3709 6613 3743 6647
rect 4905 6613 4939 6647
rect 8493 6613 8527 6647
rect 9137 6613 9171 6647
rect 10241 6613 10275 6647
rect 11621 6613 11655 6647
rect 1685 6409 1719 6443
rect 2053 6409 2087 6443
rect 2697 6409 2731 6443
rect 2789 6409 2823 6443
rect 5273 6409 5307 6443
rect 6377 6409 6411 6443
rect 9045 6409 9079 6443
rect 12173 6409 12207 6443
rect 1777 6273 1811 6307
rect 5871 6273 5905 6307
rect 6561 6341 6595 6375
rect 12449 6273 12483 6307
rect 1556 6205 1590 6239
rect 2697 6205 2731 6239
rect 2973 6205 3007 6239
rect 3433 6205 3467 6239
rect 3801 6205 3835 6239
rect 4353 6205 4387 6239
rect 5784 6205 5818 6239
rect 6377 6205 6411 6239
rect 6837 6205 6871 6239
rect 7389 6205 7423 6239
rect 8125 6205 8159 6239
rect 9873 6205 9907 6239
rect 10793 6205 10827 6239
rect 11161 6205 11195 6239
rect 12541 6205 12575 6239
rect 1409 6137 1443 6171
rect 4445 6137 4479 6171
rect 8466 6137 8500 6171
rect 9321 6137 9355 6171
rect 9689 6137 9723 6171
rect 10194 6137 10228 6171
rect 2421 6069 2455 6103
rect 4905 6069 4939 6103
rect 6193 6069 6227 6103
rect 7021 6069 7055 6103
rect 7941 6069 7975 6103
rect 11437 6069 11471 6103
rect 13737 6069 13771 6103
rect 3801 5865 3835 5899
rect 8585 5865 8619 5899
rect 12541 5865 12575 5899
rect 13047 5865 13081 5899
rect 3525 5797 3559 5831
rect 4813 5797 4847 5831
rect 6745 5797 6779 5831
rect 7665 5797 7699 5831
rect 7757 5797 7791 5831
rect 8953 5797 8987 5831
rect 9873 5797 9907 5831
rect 9965 5797 9999 5831
rect 10517 5797 10551 5831
rect 11529 5797 11563 5831
rect 1777 5729 1811 5763
rect 2329 5729 2363 5763
rect 2513 5729 2547 5763
rect 3065 5729 3099 5763
rect 5273 5729 5307 5763
rect 5733 5729 5767 5763
rect 6285 5729 6319 5763
rect 6469 5729 6503 5763
rect 7389 5729 7423 5763
rect 12944 5729 12978 5763
rect 4261 5661 4295 5695
rect 7941 5661 7975 5695
rect 10885 5661 10919 5695
rect 11437 5661 11471 5695
rect 11713 5661 11747 5695
rect 13921 5661 13955 5695
rect 3065 5593 3099 5627
rect 5089 5525 5123 5559
rect 7113 5525 7147 5559
rect 9321 5525 9355 5559
rect 11161 5525 11195 5559
rect 2421 5321 2455 5355
rect 4261 5321 4295 5355
rect 8033 5321 8067 5355
rect 8769 5321 8803 5355
rect 10241 5321 10275 5355
rect 14151 5321 14185 5355
rect 5825 5253 5859 5287
rect 13829 5253 13863 5287
rect 2053 5185 2087 5219
rect 6837 5185 6871 5219
rect 10517 5185 10551 5219
rect 10885 5185 10919 5219
rect 13461 5185 13495 5219
rect 1501 5117 1535 5151
rect 1685 5117 1719 5151
rect 2973 5117 3007 5151
rect 4445 5117 4479 5151
rect 4905 5117 4939 5151
rect 5273 5117 5307 5151
rect 5825 5117 5859 5151
rect 8953 5117 8987 5151
rect 12541 5117 12575 5151
rect 14080 5117 14114 5151
rect 14473 5117 14507 5151
rect 3617 5049 3651 5083
rect 7158 5049 7192 5083
rect 9274 5049 9308 5083
rect 10977 5049 11011 5083
rect 11529 5049 11563 5083
rect 12449 5049 12483 5083
rect 2697 4981 2731 5015
rect 3985 4981 4019 5015
rect 6193 4981 6227 5015
rect 6561 4981 6595 5015
rect 7757 4981 7791 5015
rect 8401 4981 8435 5015
rect 9873 4981 9907 5015
rect 11805 4981 11839 5015
rect 12173 4981 12207 5015
rect 1685 4777 1719 4811
rect 1961 4777 1995 4811
rect 3709 4777 3743 4811
rect 4629 4777 4663 4811
rect 7297 4777 7331 4811
rect 10885 4777 10919 4811
rect 13277 4777 13311 4811
rect 2329 4709 2363 4743
rect 6653 4709 6687 4743
rect 7573 4709 7607 4743
rect 7665 4709 7699 4743
rect 8217 4709 8251 4743
rect 8309 4709 8343 4743
rect 10010 4709 10044 4743
rect 11805 4709 11839 4743
rect 4077 4641 4111 4675
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 5641 4641 5675 4675
rect 6009 4641 6043 4675
rect 6377 4641 6411 4675
rect 2476 4573 2510 4607
rect 2697 4573 2731 4607
rect 4905 4573 4939 4607
rect 2605 4505 2639 4539
rect 2973 4505 3007 4539
rect 10609 4641 10643 4675
rect 13461 4641 13495 4675
rect 13645 4641 13679 4675
rect 8861 4573 8895 4607
rect 9689 4573 9723 4607
rect 11713 4573 11747 4607
rect 11989 4573 12023 4607
rect 8309 4505 8343 4539
rect 9229 4505 9263 4539
rect 4307 4437 4341 4471
rect 4905 4437 4939 4471
rect 6929 4437 6963 4471
rect 8585 4437 8619 4471
rect 11253 4437 11287 4471
rect 12633 4437 12667 4471
rect 13001 4437 13035 4471
rect 2191 4233 2225 4267
rect 2329 4233 2363 4267
rect 3065 4233 3099 4267
rect 3433 4233 3467 4267
rect 6193 4233 6227 4267
rect 13461 4233 13495 4267
rect 13829 4233 13863 4267
rect 4445 4165 4479 4199
rect 11161 4165 11195 4199
rect 2421 4097 2455 4131
rect 2789 4097 2823 4131
rect 5273 4097 5307 4131
rect 6837 4097 6871 4131
rect 8677 4097 8711 4131
rect 8953 4097 8987 4131
rect 10609 4097 10643 4131
rect 11989 4097 12023 4131
rect 3801 4029 3835 4063
rect 4169 4029 4203 4063
rect 12541 4029 12575 4063
rect 14048 4029 14082 4063
rect 14473 4029 14507 4063
rect 2053 3961 2087 3995
rect 4721 3961 4755 3995
rect 5365 3961 5399 3995
rect 5917 3961 5951 3995
rect 7158 3961 7192 3995
rect 8769 3961 8803 3995
rect 10425 3961 10459 3995
rect 10701 3961 10735 3995
rect 11713 3961 11747 3995
rect 12449 3961 12483 3995
rect 1869 3893 1903 3927
rect 4997 3893 5031 3927
rect 6561 3893 6595 3927
rect 7757 3893 7791 3927
rect 8033 3893 8067 3927
rect 8401 3893 8435 3927
rect 9689 3893 9723 3927
rect 14151 3893 14185 3927
rect 1547 3689 1581 3723
rect 3525 3689 3559 3723
rect 6837 3689 6871 3723
rect 11345 3689 11379 3723
rect 12541 3689 12575 3723
rect 14013 3689 14047 3723
rect 2421 3621 2455 3655
rect 6469 3621 6503 3655
rect 7481 3621 7515 3655
rect 8125 3621 8159 3655
rect 9413 3621 9447 3655
rect 10057 3621 10091 3655
rect 11621 3621 11655 3655
rect 13001 3621 13035 3655
rect 1476 3553 1510 3587
rect 2568 3553 2602 3587
rect 3893 3553 3927 3587
rect 4997 3553 5031 3587
rect 5273 3553 5307 3587
rect 5733 3553 5767 3587
rect 5917 3553 5951 3587
rect 2789 3485 2823 3519
rect 6193 3485 6227 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 4445 3417 4479 3451
rect 8309 3553 8343 3587
rect 8677 3553 8711 3587
rect 13553 3553 13587 3587
rect 15209 3553 15243 3587
rect 9965 3485 9999 3519
rect 11529 3485 11563 3519
rect 9045 3417 9079 3451
rect 10517 3417 10551 3451
rect 12081 3417 12115 3451
rect 15439 3417 15473 3451
rect 2145 3349 2179 3383
rect 2697 3349 2731 3383
rect 3065 3349 3099 3383
rect 8125 3349 8159 3383
rect 10885 3349 10919 3383
rect 12817 3349 12851 3383
rect 1685 3145 1719 3179
rect 4353 3145 4387 3179
rect 6561 3145 6595 3179
rect 11069 3145 11103 3179
rect 11529 3145 11563 3179
rect 13553 3145 13587 3179
rect 14105 3145 14139 3179
rect 3893 3077 3927 3111
rect 5825 3077 5859 3111
rect 9873 3077 9907 3111
rect 6929 3009 6963 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 9689 3009 9723 3043
rect 12541 3009 12575 3043
rect 12909 3009 12943 3043
rect 2053 2941 2087 2975
rect 2421 2941 2455 2975
rect 2697 2941 2731 2975
rect 3157 2941 3191 2975
rect 3341 2941 3375 2975
rect 4721 2941 4755 2975
rect 5089 2941 5123 2975
rect 5273 2941 5307 2975
rect 5641 2941 5675 2975
rect 8401 2941 8435 2975
rect 9321 2941 9355 2975
rect 9873 2941 9907 2975
rect 10149 2941 10183 2975
rect 11805 2941 11839 2975
rect 14749 3077 14783 3111
rect 14565 2941 14599 2975
rect 15117 2941 15151 2975
rect 15704 2941 15738 2975
rect 16129 2941 16163 2975
rect 3617 2873 3651 2907
rect 6193 2873 6227 2907
rect 7021 2873 7055 2907
rect 8309 2873 8343 2907
rect 8722 2873 8756 2907
rect 9965 2873 9999 2907
rect 10470 2873 10504 2907
rect 12633 2873 12667 2907
rect 14105 2873 14139 2907
rect 14289 2873 14323 2907
rect 15807 2873 15841 2907
rect 12265 2805 12299 2839
rect 13921 2805 13955 2839
rect 15485 2805 15519 2839
rect 1685 2601 1719 2635
rect 2145 2601 2179 2635
rect 3157 2601 3191 2635
rect 4353 2601 4387 2635
rect 5917 2601 5951 2635
rect 8815 2601 8849 2635
rect 10885 2601 10919 2635
rect 13921 2601 13955 2635
rect 15623 2601 15657 2635
rect 17141 2601 17175 2635
rect 2558 2533 2592 2567
rect 6285 2533 6319 2567
rect 6561 2533 6595 2567
rect 7250 2533 7284 2567
rect 8125 2533 8159 2567
rect 8493 2533 8527 2567
rect 9965 2533 9999 2567
rect 13553 2533 13587 2567
rect 3709 2465 3743 2499
rect 4537 2465 4571 2499
rect 4997 2465 5031 2499
rect 5365 2465 5399 2499
rect 5733 2465 5767 2499
rect 2237 2397 2271 2431
rect 3433 2397 3467 2431
rect 6929 2465 6963 2499
rect 7849 2465 7883 2499
rect 8744 2465 8778 2499
rect 10517 2465 10551 2499
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12265 2465 12299 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13725 2465 13759 2499
rect 15552 2465 15586 2499
rect 16037 2465 16071 2499
rect 16497 2465 16531 2499
rect 9873 2397 9907 2431
rect 11161 2397 11195 2431
rect 9505 2329 9539 2363
rect 11529 2329 11563 2363
rect 16681 2329 16715 2363
rect 3709 2261 3743 2295
rect 3801 2261 3835 2295
rect 6561 2261 6595 2295
rect 6653 2261 6687 2295
rect 9229 2261 9263 2295
rect 12817 2261 12851 2295
rect 14381 2261 14415 2295
<< metal1 >>
rect 14 21496 20 21548
rect 72 21536 78 21548
rect 842 21536 848 21548
rect 72 21508 848 21536
rect 72 21496 78 21508
rect 842 21496 848 21508
rect 900 21496 906 21548
rect 1670 21496 1676 21548
rect 1728 21536 1734 21548
rect 2498 21536 2504 21548
rect 1728 21508 2504 21536
rect 1728 21496 1734 21508
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 9214 21536 9220 21548
rect 8720 21508 9220 21536
rect 8720 21496 8726 21508
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 10962 21536 10968 21548
rect 9732 21508 10968 21536
rect 9732 21496 9738 21508
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 15194 21496 15200 21548
rect 15252 21536 15258 21548
rect 16022 21536 16028 21548
rect 15252 21508 16028 21536
rect 15252 21496 15258 21508
rect 16022 21496 16028 21508
rect 16080 21496 16086 21548
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17678 21536 17684 21548
rect 16632 21508 17684 21536
rect 16632 21496 16638 21508
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 19702 21496 19708 21548
rect 19760 21536 19766 21548
rect 21082 21536 21088 21548
rect 19760 21508 21088 21536
rect 19760 21496 19766 21508
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 1104 19610 20884 19632
rect 1104 19558 4648 19610
rect 4700 19558 4712 19610
rect 4764 19558 4776 19610
rect 4828 19558 4840 19610
rect 4892 19558 11982 19610
rect 12034 19558 12046 19610
rect 12098 19558 12110 19610
rect 12162 19558 12174 19610
rect 12226 19558 19315 19610
rect 19367 19558 19379 19610
rect 19431 19558 19443 19610
rect 19495 19558 19507 19610
rect 19559 19558 20884 19610
rect 1104 19536 20884 19558
rect 1104 19066 20884 19088
rect 1104 19014 8315 19066
rect 8367 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 15648 19066
rect 15700 19014 15712 19066
rect 15764 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 20884 19066
rect 1104 18992 20884 19014
rect 1104 18522 20884 18544
rect 1104 18470 4648 18522
rect 4700 18470 4712 18522
rect 4764 18470 4776 18522
rect 4828 18470 4840 18522
rect 4892 18470 11982 18522
rect 12034 18470 12046 18522
rect 12098 18470 12110 18522
rect 12162 18470 12174 18522
rect 12226 18470 19315 18522
rect 19367 18470 19379 18522
rect 19431 18470 19443 18522
rect 19495 18470 19507 18522
rect 19559 18470 20884 18522
rect 1104 18448 20884 18470
rect 6178 18408 6184 18420
rect 6139 18380 6184 18408
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 7374 18408 7380 18420
rect 7335 18380 7380 18408
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 12989 18411 13047 18417
rect 12989 18377 13001 18411
rect 13035 18408 13047 18411
rect 14458 18408 14464 18420
rect 13035 18380 14464 18408
rect 13035 18377 13047 18380
rect 12989 18371 13047 18377
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 5629 18207 5687 18213
rect 5629 18173 5641 18207
rect 5675 18204 5687 18207
rect 6178 18204 6184 18216
rect 5675 18176 6184 18204
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 7193 18207 7251 18213
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 7239 18176 7880 18204
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 7852 18077 7880 18176
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 11848 18176 12817 18204
rect 11848 18164 11854 18176
rect 12805 18173 12817 18176
rect 12851 18204 12863 18207
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 12851 18176 13369 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 13357 18173 13369 18176
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 5813 18071 5871 18077
rect 5813 18068 5825 18071
rect 5132 18040 5825 18068
rect 5132 18028 5138 18040
rect 5813 18037 5825 18040
rect 5859 18037 5871 18071
rect 5813 18031 5871 18037
rect 7837 18071 7895 18077
rect 7837 18037 7849 18071
rect 7883 18068 7895 18071
rect 8018 18068 8024 18080
rect 7883 18040 8024 18068
rect 7883 18037 7895 18040
rect 7837 18031 7895 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 1104 17978 20884 18000
rect 1104 17926 8315 17978
rect 8367 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 15648 17978
rect 15700 17926 15712 17978
rect 15764 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 20884 17978
rect 1104 17904 20884 17926
rect 4798 17864 4804 17876
rect 4759 17836 4804 17864
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 4212 17700 4629 17728
rect 4212 17688 4218 17700
rect 4617 17697 4629 17700
rect 4663 17697 4675 17731
rect 4617 17691 4675 17697
rect 1104 17434 20884 17456
rect 1104 17382 4648 17434
rect 4700 17382 4712 17434
rect 4764 17382 4776 17434
rect 4828 17382 4840 17434
rect 4892 17382 11982 17434
rect 12034 17382 12046 17434
rect 12098 17382 12110 17434
rect 12162 17382 12174 17434
rect 12226 17382 19315 17434
rect 19367 17382 19379 17434
rect 19431 17382 19443 17434
rect 19495 17382 19507 17434
rect 19559 17382 20884 17434
rect 1104 17360 20884 17382
rect 19245 17323 19303 17329
rect 19245 17289 19257 17323
rect 19291 17320 19303 17323
rect 19886 17320 19892 17332
rect 19291 17292 19892 17320
rect 19291 17289 19303 17292
rect 19245 17283 19303 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 12400 17088 19073 17116
rect 12400 17076 12406 17088
rect 19061 17085 19073 17088
rect 19107 17116 19119 17119
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 19107 17088 19625 17116
rect 19107 17085 19119 17088
rect 19061 17079 19119 17085
rect 19613 17085 19625 17088
rect 19659 17085 19671 17119
rect 19613 17079 19671 17085
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4617 16983 4675 16989
rect 4617 16980 4629 16983
rect 4212 16952 4629 16980
rect 4212 16940 4218 16952
rect 4617 16949 4629 16952
rect 4663 16949 4675 16983
rect 4617 16943 4675 16949
rect 1104 16890 20884 16912
rect 1104 16838 8315 16890
rect 8367 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 15648 16890
rect 15700 16838 15712 16890
rect 15764 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 20884 16890
rect 1104 16816 20884 16838
rect 1104 16346 20884 16368
rect 1104 16294 4648 16346
rect 4700 16294 4712 16346
rect 4764 16294 4776 16346
rect 4828 16294 4840 16346
rect 4892 16294 11982 16346
rect 12034 16294 12046 16346
rect 12098 16294 12110 16346
rect 12162 16294 12174 16346
rect 12226 16294 19315 16346
rect 19367 16294 19379 16346
rect 19431 16294 19443 16346
rect 19495 16294 19507 16346
rect 19559 16294 20884 16346
rect 1104 16272 20884 16294
rect 1104 15802 20884 15824
rect 1104 15750 8315 15802
rect 8367 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 15648 15802
rect 15700 15750 15712 15802
rect 15764 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 20884 15802
rect 1104 15728 20884 15750
rect 1104 15258 20884 15280
rect 1104 15206 4648 15258
rect 4700 15206 4712 15258
rect 4764 15206 4776 15258
rect 4828 15206 4840 15258
rect 4892 15206 11982 15258
rect 12034 15206 12046 15258
rect 12098 15206 12110 15258
rect 12162 15206 12174 15258
rect 12226 15206 19315 15258
rect 19367 15206 19379 15258
rect 19431 15206 19443 15258
rect 19495 15206 19507 15258
rect 19559 15206 20884 15258
rect 1104 15184 20884 15206
rect 1104 14714 20884 14736
rect 1104 14662 8315 14714
rect 8367 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 15648 14714
rect 15700 14662 15712 14714
rect 15764 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 20884 14714
rect 1104 14640 20884 14662
rect 19058 14464 19064 14476
rect 19019 14436 19064 14464
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 19150 14220 19156 14272
rect 19208 14260 19214 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 19208 14232 19257 14260
rect 19208 14220 19214 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 1104 14170 20884 14192
rect 1104 14118 4648 14170
rect 4700 14118 4712 14170
rect 4764 14118 4776 14170
rect 4828 14118 4840 14170
rect 4892 14118 11982 14170
rect 12034 14118 12046 14170
rect 12098 14118 12110 14170
rect 12162 14118 12174 14170
rect 12226 14118 19315 14170
rect 19367 14118 19379 14170
rect 19431 14118 19443 14170
rect 19495 14118 19507 14170
rect 19559 14118 20884 14170
rect 1104 14096 20884 14118
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 1104 13626 20884 13648
rect 1104 13574 8315 13626
rect 8367 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 15648 13626
rect 15700 13574 15712 13626
rect 15764 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 20884 13626
rect 1104 13552 20884 13574
rect 1104 13082 20884 13104
rect 1104 13030 4648 13082
rect 4700 13030 4712 13082
rect 4764 13030 4776 13082
rect 4828 13030 4840 13082
rect 4892 13030 11982 13082
rect 12034 13030 12046 13082
rect 12098 13030 12110 13082
rect 12162 13030 12174 13082
rect 12226 13030 19315 13082
rect 19367 13030 19379 13082
rect 19431 13030 19443 13082
rect 19495 13030 19507 13082
rect 19559 13030 20884 13082
rect 1104 13008 20884 13030
rect 1104 12538 20884 12560
rect 1104 12486 8315 12538
rect 8367 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 15648 12538
rect 15700 12486 15712 12538
rect 15764 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 20884 12538
rect 1104 12464 20884 12486
rect 1104 11994 20884 12016
rect 1104 11942 4648 11994
rect 4700 11942 4712 11994
rect 4764 11942 4776 11994
rect 4828 11942 4840 11994
rect 4892 11942 11982 11994
rect 12034 11942 12046 11994
rect 12098 11942 12110 11994
rect 12162 11942 12174 11994
rect 12226 11942 19315 11994
rect 19367 11942 19379 11994
rect 19431 11942 19443 11994
rect 19495 11942 19507 11994
rect 19559 11942 20884 11994
rect 1104 11920 20884 11942
rect 1578 11812 1584 11824
rect 1539 11784 1584 11812
rect 1578 11772 1584 11784
rect 1636 11772 1642 11824
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1360 11648 1409 11676
rect 1360 11636 1366 11648
rect 1397 11645 1409 11648
rect 1443 11676 1455 11679
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1443 11648 1961 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1949 11645 1961 11648
rect 1995 11676 2007 11679
rect 2590 11676 2596 11688
rect 1995 11648 2596 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 8088 11679 8146 11685
rect 8088 11645 8100 11679
rect 8134 11676 8146 11679
rect 8134 11648 8616 11676
rect 8134 11645 8146 11648
rect 8088 11639 8146 11645
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 8588 11549 8616 11648
rect 8159 11543 8217 11549
rect 8159 11540 8171 11543
rect 7156 11512 8171 11540
rect 7156 11500 7162 11512
rect 8159 11509 8171 11512
rect 8205 11509 8217 11543
rect 8159 11503 8217 11509
rect 8573 11543 8631 11549
rect 8573 11509 8585 11543
rect 8619 11540 8631 11543
rect 9030 11540 9036 11552
rect 8619 11512 9036 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9030 11500 9036 11512
rect 9088 11540 9094 11552
rect 9674 11540 9680 11552
rect 9088 11512 9680 11540
rect 9088 11500 9094 11512
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 1104 11450 20884 11472
rect 1104 11398 8315 11450
rect 8367 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 15648 11450
rect 15700 11398 15712 11450
rect 15764 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 20884 11450
rect 1104 11376 20884 11398
rect 7098 11336 7104 11348
rect 7059 11308 7104 11336
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 2590 11200 2596 11212
rect 2551 11172 2596 11200
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 5537 11203 5595 11209
rect 5537 11200 5549 11203
rect 4304 11172 5549 11200
rect 4304 11160 4310 11172
rect 5537 11169 5549 11172
rect 5583 11200 5595 11203
rect 5626 11200 5632 11212
rect 5583 11172 5632 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6638 11200 6644 11212
rect 6595 11172 6644 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 8202 11200 8208 11212
rect 7616 11172 8208 11200
rect 7616 11160 7622 11172
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 12434 11200 12440 11212
rect 12395 11172 12440 11200
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 7374 11064 7380 11076
rect 6328 11036 7380 11064
rect 6328 11024 6334 11036
rect 7374 11024 7380 11036
rect 7432 11064 7438 11076
rect 8662 11064 8668 11076
rect 7432 11036 8668 11064
rect 7432 11024 7438 11036
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 2823 10999 2881 11005
rect 2823 10965 2835 10999
rect 2869 10996 2881 10999
rect 3602 10996 3608 11008
rect 2869 10968 3608 10996
rect 2869 10965 2881 10968
rect 2823 10959 2881 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 3786 10996 3792 11008
rect 3747 10968 3792 10996
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 5675 10999 5733 11005
rect 5675 10965 5687 10999
rect 5721 10996 5733 10999
rect 5994 10996 6000 11008
rect 5721 10968 6000 10996
rect 5721 10965 5733 10968
rect 5675 10959 5733 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6546 10956 6552 11008
rect 6604 10996 6610 11008
rect 6687 10999 6745 11005
rect 6687 10996 6699 10999
rect 6604 10968 6699 10996
rect 6604 10956 6610 10968
rect 6687 10965 6699 10968
rect 6733 10965 6745 10999
rect 6687 10959 6745 10965
rect 8343 10999 8401 11005
rect 8343 10965 8355 10999
rect 8389 10996 8401 10999
rect 9306 10996 9312 11008
rect 8389 10968 9312 10996
rect 8389 10965 8401 10968
rect 8343 10959 8401 10965
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 1104 10906 20884 10928
rect 1104 10854 4648 10906
rect 4700 10854 4712 10906
rect 4764 10854 4776 10906
rect 4828 10854 4840 10906
rect 4892 10854 11982 10906
rect 12034 10854 12046 10906
rect 12098 10854 12110 10906
rect 12162 10854 12174 10906
rect 12226 10854 19315 10906
rect 19367 10854 19379 10906
rect 19431 10854 19443 10906
rect 19495 10854 19507 10906
rect 19559 10854 20884 10906
rect 1104 10832 20884 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1452 10764 1593 10792
rect 1452 10752 1458 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 2648 10764 3341 10792
rect 2648 10752 2654 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 3329 10755 3387 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12492 10764 12633 10792
rect 12492 10752 12498 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 4430 10684 4436 10736
rect 4488 10724 4494 10736
rect 4488 10696 7236 10724
rect 4488 10684 4494 10696
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3660 10628 3801 10656
rect 3660 10616 3666 10628
rect 3789 10625 3801 10628
rect 3835 10656 3847 10659
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 3835 10628 4721 10656
rect 3835 10625 3847 10628
rect 3789 10619 3847 10625
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7098 10656 7104 10668
rect 6963 10628 7104 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7208 10665 7236 10696
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7558 10656 7564 10668
rect 7239 10628 7564 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10588 1458 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1452 10560 1961 10588
rect 1452 10548 1458 10560
rect 1949 10557 1961 10560
rect 1995 10588 2007 10591
rect 2536 10591 2594 10597
rect 2536 10588 2548 10591
rect 1995 10560 2548 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2536 10557 2548 10560
rect 2582 10588 2594 10591
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2582 10560 2973 10588
rect 2582 10557 2594 10560
rect 2536 10551 2594 10557
rect 2961 10557 2973 10560
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 5772 10591 5830 10597
rect 5772 10557 5784 10591
rect 5818 10588 5830 10591
rect 6270 10588 6276 10600
rect 5818 10560 6276 10588
rect 5818 10557 5830 10560
rect 5772 10551 5830 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8424 10591 8482 10597
rect 8424 10588 8436 10591
rect 7984 10560 8436 10588
rect 7984 10548 7990 10560
rect 8424 10557 8436 10560
rect 8470 10588 8482 10591
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8470 10560 8861 10588
rect 8470 10557 8482 10560
rect 8424 10551 8482 10557
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 3786 10480 3792 10532
rect 3844 10520 3850 10532
rect 3881 10523 3939 10529
rect 3881 10520 3893 10523
rect 3844 10492 3893 10520
rect 3844 10480 3850 10492
rect 3881 10489 3893 10492
rect 3927 10489 3939 10523
rect 4430 10520 4436 10532
rect 4391 10492 4436 10520
rect 3881 10483 3939 10489
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 5859 10523 5917 10529
rect 5859 10489 5871 10523
rect 5905 10520 5917 10523
rect 6914 10520 6920 10532
rect 5905 10492 6920 10520
rect 5905 10489 5917 10492
rect 5859 10483 5917 10489
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 8527 10523 8585 10529
rect 7064 10492 7109 10520
rect 7064 10480 7070 10492
rect 8527 10489 8539 10523
rect 8573 10520 8585 10523
rect 12434 10520 12440 10532
rect 8573 10492 12440 10520
rect 8573 10489 8585 10492
rect 8527 10483 8585 10489
rect 12434 10480 12440 10492
rect 12492 10480 12498 10532
rect 2639 10455 2697 10461
rect 2639 10421 2651 10455
rect 2685 10452 2697 10455
rect 4982 10452 4988 10464
rect 2685 10424 4988 10452
rect 2685 10421 2697 10424
rect 2639 10415 2697 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 5626 10452 5632 10464
rect 5587 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8297 10455 8355 10461
rect 8297 10452 8309 10455
rect 8260 10424 8309 10452
rect 8260 10412 8266 10424
rect 8297 10421 8309 10424
rect 8343 10452 8355 10455
rect 8846 10452 8852 10464
rect 8343 10424 8852 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 10318 10452 10324 10464
rect 10279 10424 10324 10452
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 1104 10362 20884 10384
rect 1104 10310 8315 10362
rect 8367 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 15648 10362
rect 15700 10310 15712 10362
rect 15764 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 20884 10362
rect 1104 10288 20884 10310
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10376 10220 10793 10248
rect 10376 10208 10382 10220
rect 10781 10217 10793 10220
rect 10827 10248 10839 10251
rect 10870 10248 10876 10260
rect 10827 10220 10876 10248
rect 10827 10217 10839 10220
rect 10781 10211 10839 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15252 10220 15485 10248
rect 15252 10208 15258 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 3881 10183 3939 10189
rect 3881 10149 3893 10183
rect 3927 10180 3939 10183
rect 4246 10180 4252 10192
rect 3927 10152 4252 10180
rect 3927 10149 3939 10152
rect 3881 10143 3939 10149
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 4801 10183 4859 10189
rect 4801 10180 4813 10183
rect 4488 10152 4813 10180
rect 4488 10140 4494 10152
rect 4801 10149 4813 10152
rect 4847 10149 4859 10183
rect 4801 10143 4859 10149
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 5077 10183 5135 10189
rect 5077 10180 5089 10183
rect 5040 10152 5089 10180
rect 5040 10140 5046 10152
rect 5077 10149 5089 10152
rect 5123 10149 5135 10183
rect 5994 10180 6000 10192
rect 5955 10152 6000 10180
rect 5077 10143 5135 10149
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 6089 10183 6147 10189
rect 6089 10149 6101 10183
rect 6135 10180 6147 10183
rect 6270 10180 6276 10192
rect 6135 10152 6276 10180
rect 6135 10149 6147 10152
rect 6089 10143 6147 10149
rect 6270 10140 6276 10152
rect 6328 10180 6334 10192
rect 7006 10180 7012 10192
rect 6328 10152 7012 10180
rect 6328 10140 6334 10152
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 7558 10180 7564 10192
rect 7519 10152 7564 10180
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 7653 10183 7711 10189
rect 7653 10149 7665 10183
rect 7699 10180 7711 10183
rect 7742 10180 7748 10192
rect 7699 10152 7748 10180
rect 7699 10149 7711 10152
rect 7653 10143 7711 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 12391 10183 12449 10189
rect 12391 10149 12403 10183
rect 12437 10180 12449 10183
rect 17218 10180 17224 10192
rect 12437 10152 17224 10180
rect 12437 10149 12449 10152
rect 12391 10143 12449 10149
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3878 10044 3884 10056
rect 3007 10016 3884 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 5000 10044 5028 10140
rect 10226 10112 10232 10124
rect 10187 10084 10232 10112
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11308 10115 11366 10121
rect 11308 10081 11320 10115
rect 11354 10112 11366 10115
rect 11514 10112 11520 10124
rect 11354 10084 11520 10112
rect 11354 10081 11366 10084
rect 11308 10075 11366 10081
rect 11514 10072 11520 10084
rect 11572 10112 11578 10124
rect 12158 10112 12164 10124
rect 11572 10084 12164 10112
rect 11572 10072 11578 10084
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12304 10115 12362 10121
rect 12304 10081 12316 10115
rect 12350 10112 12362 10115
rect 12526 10112 12532 10124
rect 12350 10084 12532 10112
rect 12350 10081 12362 10084
rect 12304 10075 12362 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 15378 10112 15384 10124
rect 15335 10084 15384 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 4203 10016 5028 10044
rect 6641 10047 6699 10053
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 7190 10044 7196 10056
rect 6687 10016 7196 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 3016 9880 3249 9908
rect 3016 9868 3022 9880
rect 3237 9877 3249 9880
rect 3283 9877 3295 9911
rect 3237 9871 3295 9877
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 11379 9911 11437 9917
rect 11379 9908 11391 9911
rect 11296 9880 11391 9908
rect 11296 9868 11302 9880
rect 11379 9877 11391 9880
rect 11425 9877 11437 9911
rect 11379 9871 11437 9877
rect 1104 9818 20884 9840
rect 1104 9766 4648 9818
rect 4700 9766 4712 9818
rect 4764 9766 4776 9818
rect 4828 9766 4840 9818
rect 4892 9766 11982 9818
rect 12034 9766 12046 9818
rect 12098 9766 12110 9818
rect 12162 9766 12174 9818
rect 12226 9766 19315 9818
rect 19367 9766 19379 9818
rect 19431 9766 19443 9818
rect 19495 9766 19507 9818
rect 19559 9766 20884 9818
rect 1104 9744 20884 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 2556 9676 2697 9704
rect 2556 9664 2562 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 2685 9667 2743 9673
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6270 9704 6276 9716
rect 5951 9676 6276 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7616 9676 8217 9704
rect 7616 9664 7622 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 8205 9667 8263 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 4157 9639 4215 9645
rect 4157 9636 4169 9639
rect 3844 9608 4169 9636
rect 3844 9596 3850 9608
rect 4157 9605 4169 9608
rect 4203 9636 4215 9639
rect 6730 9636 6736 9648
rect 4203 9608 6736 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 12434 9636 12440 9648
rect 8076 9608 12440 9636
rect 8076 9596 8082 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 6914 9568 6920 9580
rect 6875 9540 6920 9568
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7190 9568 7196 9580
rect 7151 9540 7196 9568
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 10870 9568 10876 9580
rect 10831 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 11146 9568 11152 9580
rect 11107 9540 11152 9568
rect 11146 9528 11152 9540
rect 11204 9568 11210 9580
rect 12526 9568 12532 9580
rect 11204 9540 12532 9568
rect 11204 9528 11210 9540
rect 12526 9528 12532 9540
rect 12584 9568 12590 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12584 9540 12633 9568
rect 12584 9528 12590 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1728 9472 1777 9500
rect 1728 9460 1734 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 3016 9472 3249 9500
rect 3016 9460 3022 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 4522 9500 4528 9512
rect 4435 9472 4528 9500
rect 3237 9463 3295 9469
rect 4522 9460 4528 9472
rect 4580 9500 4586 9512
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4580 9472 4997 9500
rect 4580 9460 4586 9472
rect 4985 9469 4997 9472
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 3599 9435 3657 9441
rect 3599 9401 3611 9435
rect 3645 9401 3657 9435
rect 3599 9395 3657 9401
rect 5306 9435 5364 9441
rect 5306 9401 5318 9435
rect 5352 9401 5364 9435
rect 5306 9395 5364 9401
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3053 9367 3111 9373
rect 3053 9364 3065 9367
rect 2740 9336 3065 9364
rect 2740 9324 2746 9336
rect 3053 9333 3065 9336
rect 3099 9364 3111 9367
rect 3614 9364 3642 9395
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 3099 9336 4813 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 4801 9333 4813 9336
rect 4847 9364 4859 9367
rect 5321 9364 5349 9395
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 5592 9404 6653 9432
rect 5592 9392 5598 9404
rect 6641 9401 6653 9404
rect 6687 9432 6699 9435
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6687 9404 7021 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9674 9432 9680 9444
rect 9447 9404 9680 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 4847 9336 5349 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7800 9336 7849 9364
rect 7800 9324 7806 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 9125 9367 9183 9373
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 9416 9364 9444 9395
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9950 9432 9956 9444
rect 9911 9404 9956 9432
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 10962 9432 10968 9444
rect 10735 9404 10968 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 9171 9336 9444 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11572 9336 11805 9364
rect 11572 9324 11578 9336
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 15378 9364 15384 9376
rect 15339 9336 15384 9364
rect 11793 9327 11851 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 1104 9274 20884 9296
rect 1104 9222 8315 9274
rect 8367 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 15648 9274
rect 15700 9222 15712 9274
rect 15764 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 20884 9274
rect 1104 9200 20884 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 4246 9160 4252 9172
rect 3191 9132 4252 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 2587 9095 2645 9101
rect 2587 9061 2599 9095
rect 2633 9092 2645 9095
rect 2682 9092 2688 9104
rect 2633 9064 2688 9092
rect 2633 9061 2645 9064
rect 2587 9055 2645 9061
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 4126 9092 4154 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 5994 9160 6000 9172
rect 5955 9132 6000 9160
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6457 9163 6515 9169
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 6546 9160 6552 9172
rect 6503 9132 6552 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6546 9120 6552 9132
rect 6604 9160 6610 9172
rect 9306 9160 9312 9172
rect 6604 9132 6684 9160
rect 9267 9132 9312 9160
rect 6604 9120 6610 9132
rect 5534 9092 5540 9104
rect 4126 9064 5540 9092
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 6656 9101 6684 9132
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 10612 9132 12388 9160
rect 10612 9104 10640 9132
rect 6641 9095 6699 9101
rect 6641 9061 6653 9095
rect 6687 9061 6699 9095
rect 6641 9055 6699 9061
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 8018 9092 8024 9104
rect 6788 9064 8024 9092
rect 6788 9052 6794 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 9950 9052 9956 9104
rect 10008 9092 10014 9104
rect 10502 9092 10508 9104
rect 10008 9064 10508 9092
rect 10008 9052 10014 9064
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 10652 9064 10745 9092
rect 10652 9052 10658 9064
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 11977 9095 12035 9101
rect 11977 9092 11989 9095
rect 11020 9064 11989 9092
rect 11020 9052 11026 9064
rect 11977 9061 11989 9064
rect 12023 9061 12035 9095
rect 11977 9055 12035 9061
rect 12360 9036 12388 9132
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4433 8987 4491 8993
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 1820 8928 2237 8956
rect 1820 8916 1826 8928
rect 2225 8925 2237 8928
rect 2271 8956 2283 8959
rect 2866 8956 2872 8968
rect 2271 8928 2872 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8888 3571 8891
rect 3786 8888 3792 8900
rect 3559 8860 3792 8888
rect 3559 8857 3571 8860
rect 3513 8851 3571 8857
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4448 8888 4476 8987
rect 4614 8984 4620 9036
rect 4672 9024 4678 9036
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 4672 8996 4721 9024
rect 4672 8984 4678 8996
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 5040 8996 5089 9024
rect 5040 8984 5046 8996
rect 5077 8993 5089 8996
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 8640 9027 8698 9033
rect 8640 8993 8652 9027
rect 8686 9024 8698 9027
rect 9030 9024 9036 9036
rect 8686 8996 9036 9024
rect 8686 8993 8698 8996
rect 8640 8987 8698 8993
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 5460 8956 5488 8987
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 12342 9024 12348 9036
rect 11204 8996 11249 9024
rect 12303 8996 12348 9024
rect 11204 8984 11210 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 4580 8928 5488 8956
rect 4580 8916 4586 8928
rect 5166 8888 5172 8900
rect 4448 8860 5172 8888
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 7190 8888 7196 8900
rect 7151 8860 7196 8888
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 8711 8891 8769 8897
rect 8711 8857 8723 8891
rect 8757 8888 8769 8891
rect 9674 8888 9680 8900
rect 8757 8860 9680 8888
rect 8757 8857 8769 8860
rect 8711 8851 8769 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 2130 8820 2136 8832
rect 2091 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 7558 8820 7564 8832
rect 7519 8792 7564 8820
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9364 8792 9873 8820
rect 9364 8780 9370 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 9861 8783 9919 8789
rect 1104 8730 20884 8752
rect 1104 8678 4648 8730
rect 4700 8678 4712 8730
rect 4764 8678 4776 8730
rect 4828 8678 4840 8730
rect 4892 8678 11982 8730
rect 12034 8678 12046 8730
rect 12098 8678 12110 8730
rect 12162 8678 12174 8730
rect 12226 8678 19315 8730
rect 19367 8678 19379 8730
rect 19431 8678 19443 8730
rect 19495 8678 19507 8730
rect 19559 8678 20884 8730
rect 1104 8656 20884 8678
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 10226 8616 10232 8628
rect 9539 8588 10232 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10594 8616 10600 8628
rect 10428 8588 10600 8616
rect 9861 8551 9919 8557
rect 9861 8517 9873 8551
rect 9907 8548 9919 8551
rect 10428 8548 10456 8588
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 11296 8588 11345 8616
rect 11296 8576 11302 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 11333 8579 11391 8585
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12342 8616 12348 8628
rect 12115 8588 12348 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 9907 8520 10456 8548
rect 9907 8517 9919 8520
rect 9861 8511 9919 8517
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 10560 8520 10977 8548
rect 10560 8508 10566 8520
rect 10965 8517 10977 8520
rect 11011 8548 11023 8551
rect 11146 8548 11152 8560
rect 11011 8520 11152 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2682 8480 2688 8492
rect 2363 8452 2688 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2682 8440 2688 8452
rect 2740 8480 2746 8492
rect 8573 8483 8631 8489
rect 2740 8452 3648 8480
rect 2740 8440 2746 8452
rect 2777 8415 2835 8421
rect 2777 8412 2789 8415
rect 2700 8384 2789 8412
rect 2700 8288 2728 8384
rect 2777 8381 2789 8384
rect 2823 8381 2835 8415
rect 3326 8412 3332 8424
rect 3287 8384 3332 8412
rect 2777 8375 2835 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3620 8344 3648 8452
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8938 8480 8944 8492
rect 8619 8452 8944 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 11256 8480 11284 8576
rect 10459 8452 11284 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 3786 8412 3792 8424
rect 3747 8384 3792 8412
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3936 8384 4169 8412
rect 3936 8372 3942 8384
rect 4157 8381 4169 8384
rect 4203 8412 4215 8415
rect 4522 8412 4528 8424
rect 4203 8384 4528 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5166 8412 5172 8424
rect 5031 8384 5172 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5718 8412 5724 8424
rect 5631 8384 5724 8412
rect 5718 8372 5724 8384
rect 5776 8412 5782 8424
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 5776 8384 6101 8412
rect 5776 8372 5782 8384
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6328 8384 6837 8412
rect 6328 8372 6334 8384
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 7558 8412 7564 8424
rect 6871 8384 7564 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12472 8415 12530 8421
rect 12472 8412 12484 8415
rect 11296 8384 12484 8412
rect 11296 8372 11302 8384
rect 12472 8381 12484 8384
rect 12518 8381 12530 8415
rect 12472 8375 12530 8381
rect 12575 8415 12633 8421
rect 12575 8381 12587 8415
rect 12621 8412 12633 8415
rect 12710 8412 12716 8424
rect 12621 8384 12716 8412
rect 12621 8381 12633 8384
rect 12575 8375 12633 8381
rect 5074 8344 5080 8356
rect 3620 8316 4936 8344
rect 5035 8316 5080 8344
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 2682 8276 2688 8288
rect 2643 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 2866 8276 2872 8288
rect 2827 8248 2872 8276
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 3660 8248 4537 8276
rect 3660 8236 3666 8248
rect 4525 8245 4537 8248
rect 4571 8276 4583 8279
rect 4798 8276 4804 8288
rect 4571 8248 4804 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 4908 8276 4936 8316
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 7146 8347 7204 8353
rect 7146 8313 7158 8347
rect 7192 8313 7204 8347
rect 7146 8307 7204 8313
rect 6546 8276 6552 8288
rect 4908 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8276 6610 8288
rect 7161 8276 7189 8307
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 8894 8347 8952 8353
rect 8894 8344 8906 8347
rect 8812 8316 8906 8344
rect 8812 8304 8818 8316
rect 8894 8313 8906 8316
rect 8940 8313 8952 8347
rect 8894 8307 8952 8313
rect 10505 8347 10563 8353
rect 10505 8313 10517 8347
rect 10551 8313 10563 8347
rect 12487 8344 12515 8375
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12487 8316 12909 8344
rect 10505 8307 10563 8313
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 6604 8248 7189 8276
rect 6604 8236 6610 8248
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 7340 8248 7757 8276
rect 7340 8236 7346 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8276 8539 8279
rect 9030 8276 9036 8288
rect 8527 8248 9036 8276
rect 8527 8245 8539 8248
rect 8481 8239 8539 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 10520 8276 10548 8307
rect 10284 8248 10548 8276
rect 10284 8236 10290 8248
rect 1104 8186 20884 8208
rect 1104 8134 8315 8186
rect 8367 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 15648 8186
rect 15700 8134 15712 8186
rect 15764 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 20884 8186
rect 1104 8112 20884 8134
rect 3694 8032 3700 8084
rect 3752 8072 3758 8084
rect 5074 8072 5080 8084
rect 3752 8044 5080 8072
rect 3752 8032 3758 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 10594 8072 10600 8084
rect 10555 8044 10600 8072
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 11204 8044 11253 8072
rect 11204 8032 11210 8044
rect 11241 8041 11253 8044
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 2130 8004 2136 8016
rect 2091 7976 2136 8004
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 4430 8004 4436 8016
rect 4304 7976 4436 8004
rect 4304 7964 4310 7976
rect 4430 7964 4436 7976
rect 4488 8004 4494 8016
rect 6270 8004 6276 8016
rect 4488 7976 5304 8004
rect 6231 7976 6276 8004
rect 4488 7964 4494 7976
rect 1026 7896 1032 7948
rect 1084 7936 1090 7948
rect 1489 7939 1547 7945
rect 1489 7936 1501 7939
rect 1084 7908 1501 7936
rect 1084 7896 1090 7908
rect 1489 7905 1501 7908
rect 1535 7936 1547 7939
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 1535 7908 2421 7936
rect 1535 7905 1547 7908
rect 1489 7899 1547 7905
rect 2409 7905 2421 7908
rect 2455 7905 2467 7939
rect 4982 7936 4988 7948
rect 4943 7908 4988 7936
rect 2409 7899 2467 7905
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 5276 7945 5304 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 7282 8004 7288 8016
rect 7243 7976 7288 8004
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 9998 8007 10056 8013
rect 9998 7973 10010 8007
rect 10044 7973 10056 8007
rect 9998 7967 10056 7973
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7905 5319 7939
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5261 7899 5319 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2832 7840 3157 7868
rect 2832 7828 2838 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 6012 7868 6040 7899
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 7892 7908 8585 7936
rect 7892 7896 7898 7908
rect 8573 7905 8585 7908
rect 8619 7936 8631 7939
rect 8754 7936 8760 7948
rect 8619 7908 8760 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8754 7896 8760 7908
rect 8812 7936 8818 7948
rect 10013 7936 10041 7967
rect 10870 7964 10876 8016
rect 10928 8004 10934 8016
rect 10965 8007 11023 8013
rect 10965 8004 10977 8007
rect 10928 7976 10977 8004
rect 10928 7964 10934 7976
rect 10965 7973 10977 7976
rect 11011 8004 11023 8007
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 11011 7976 13001 8004
rect 11011 7973 11023 7976
rect 10965 7967 11023 7973
rect 12989 7973 13001 7976
rect 13035 7973 13047 8007
rect 12989 7967 13047 7973
rect 10226 7936 10232 7948
rect 8812 7908 10232 7936
rect 8812 7896 8818 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11698 7936 11704 7948
rect 11659 7908 11704 7936
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 11931 7908 12112 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 6454 7868 6460 7880
rect 3145 7831 3203 7837
rect 4632 7840 6460 7868
rect 2866 7732 2872 7744
rect 2827 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3694 7732 3700 7744
rect 3651 7704 3700 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4522 7692 4528 7744
rect 4580 7732 4586 7744
rect 4632 7741 4660 7840
rect 6454 7828 6460 7840
rect 6512 7868 6518 7880
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6512 7840 6561 7868
rect 6512 7828 6518 7840
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 6549 7831 6607 7837
rect 7190 7828 7196 7840
rect 7248 7868 7254 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7248 7840 8125 7868
rect 7248 7828 7254 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9180 7840 9689 7868
rect 9180 7828 9186 7840
rect 9677 7837 9689 7840
rect 9723 7868 9735 7871
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 9723 7840 11989 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 7926 7800 7932 7812
rect 7791 7772 7932 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 11882 7800 11888 7812
rect 8496 7772 11888 7800
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 4580 7704 4629 7732
rect 4580 7692 4586 7704
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 4617 7695 4675 7701
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6696 7704 6929 7732
rect 6696 7692 6702 7704
rect 6917 7701 6929 7704
rect 6963 7732 6975 7735
rect 8496 7732 8524 7772
rect 11882 7760 11888 7772
rect 11940 7800 11946 7812
rect 12084 7800 12112 7908
rect 11940 7772 12112 7800
rect 11940 7760 11946 7772
rect 8938 7732 8944 7744
rect 6963 7704 8524 7732
rect 8899 7704 8944 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 9272 7704 9321 7732
rect 9272 7692 9278 7704
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 1104 7642 20884 7664
rect 1104 7590 4648 7642
rect 4700 7590 4712 7642
rect 4764 7590 4776 7642
rect 4828 7590 4840 7642
rect 4892 7590 11982 7642
rect 12034 7590 12046 7642
rect 12098 7590 12110 7642
rect 12162 7590 12174 7642
rect 12226 7590 19315 7642
rect 19367 7590 19379 7642
rect 19431 7590 19443 7642
rect 19495 7590 19507 7642
rect 19559 7590 20884 7642
rect 1104 7568 20884 7590
rect 14 7488 20 7540
rect 72 7528 78 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 72 7500 2513 7528
rect 72 7488 78 7500
rect 2501 7497 2513 7500
rect 2547 7528 2559 7531
rect 3602 7528 3608 7540
rect 2547 7500 3608 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 3602 7488 3608 7500
rect 3660 7528 3666 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 3660 7500 4997 7528
rect 3660 7488 3666 7500
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 7742 7528 7748 7540
rect 7703 7500 7748 7528
rect 4985 7491 5043 7497
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 4522 7460 4528 7472
rect 2096 7432 4528 7460
rect 2096 7420 2102 7432
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 2866 7392 2872 7404
rect 2280 7364 2872 7392
rect 2280 7352 2286 7364
rect 2866 7352 2872 7364
rect 2924 7392 2930 7404
rect 2924 7364 3372 7392
rect 2924 7352 2930 7364
rect 3344 7336 3372 7364
rect 106 7284 112 7336
rect 164 7324 170 7336
rect 1397 7327 1455 7333
rect 1397 7324 1409 7327
rect 164 7296 1409 7324
rect 164 7284 170 7296
rect 1397 7293 1409 7296
rect 1443 7324 1455 7327
rect 1578 7324 1584 7336
rect 1443 7296 1584 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3326 7324 3332 7336
rect 3239 7296 3332 7324
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 3988 7333 4016 7432
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 5000 7324 5028 7491
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 9122 7528 9128 7540
rect 9083 7500 9128 7528
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10226 7528 10232 7540
rect 10187 7500 10232 7528
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 6270 7460 6276 7472
rect 5868 7432 6276 7460
rect 5868 7420 5874 7432
rect 6270 7420 6276 7432
rect 6328 7460 6334 7472
rect 11698 7460 11704 7472
rect 6328 7432 11704 7460
rect 6328 7420 6334 7432
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11940 7432 12173 7460
rect 11940 7420 11946 7432
rect 12161 7429 12173 7432
rect 12207 7429 12219 7463
rect 12161 7423 12219 7429
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 8938 7392 8944 7404
rect 5951 7364 8944 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 5000 7296 5181 7324
rect 3973 7287 4031 7293
rect 5169 7293 5181 7296
rect 5215 7324 5227 7327
rect 5258 7324 5264 7336
rect 5215 7296 5264 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6638 7324 6644 7336
rect 5675 7296 6644 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 2866 7216 2872 7268
rect 2924 7256 2930 7268
rect 5644 7256 5672 7287
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7324 6886 7336
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 6880 7296 8033 7324
rect 6880 7284 6886 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12483 7296 13124 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 2924 7228 5672 7256
rect 7146 7259 7204 7265
rect 2924 7216 2930 7228
rect 7146 7225 7158 7259
rect 7192 7225 7204 7259
rect 9306 7256 9312 7268
rect 9267 7228 9312 7256
rect 7146 7219 7204 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2222 7188 2228 7200
rect 2183 7160 2228 7188
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 4246 7188 4252 7200
rect 3384 7160 4252 7188
rect 3384 7148 3390 7160
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4304 7160 4629 7188
rect 4304 7148 4310 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6604 7160 6653 7188
rect 6604 7148 6610 7160
rect 6641 7157 6653 7160
rect 6687 7188 6699 7191
rect 7161 7188 7189 7219
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 9953 7259 10011 7265
rect 9456 7228 9501 7256
rect 9456 7216 9462 7228
rect 9953 7225 9965 7259
rect 9999 7256 10011 7259
rect 10594 7256 10600 7268
rect 9999 7228 10600 7256
rect 9999 7225 10011 7228
rect 9953 7219 10011 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 10689 7259 10747 7265
rect 10689 7225 10701 7259
rect 10735 7256 10747 7259
rect 10962 7256 10968 7268
rect 10735 7228 10968 7256
rect 10735 7225 10747 7228
rect 10689 7219 10747 7225
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 7834 7188 7840 7200
rect 6687 7160 7840 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 8757 7191 8815 7197
rect 8757 7157 8769 7191
rect 8803 7188 8815 7191
rect 9416 7188 9444 7216
rect 13096 7200 13124 7296
rect 8803 7160 9444 7188
rect 8803 7157 8815 7160
rect 8757 7151 8815 7157
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11756 7160 11897 7188
rect 11756 7148 11762 7160
rect 11885 7157 11897 7160
rect 11931 7188 11943 7191
rect 12618 7188 12624 7200
rect 11931 7160 12624 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 13078 7188 13084 7200
rect 13039 7160 13084 7188
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 1104 7098 20884 7120
rect 1104 7046 8315 7098
rect 8367 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 15648 7098
rect 15700 7046 15712 7098
rect 15764 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 20884 7098
rect 1104 7024 20884 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 2041 6987 2099 6993
rect 2041 6953 2053 6987
rect 2087 6984 2099 6987
rect 2498 6984 2504 6996
rect 2087 6956 2504 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 5718 6984 5724 6996
rect 3467 6956 5724 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 1762 6876 1768 6928
rect 1820 6916 1826 6928
rect 3436 6916 3464 6947
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7340 6956 7389 6984
rect 7340 6944 7346 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7892 6956 7941 6984
rect 7892 6944 7898 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 13771 6987 13829 6993
rect 13771 6984 13783 6987
rect 9364 6956 13783 6984
rect 9364 6944 9370 6956
rect 13771 6953 13783 6956
rect 13817 6953 13829 6987
rect 13771 6947 13829 6953
rect 1820 6888 3464 6916
rect 1820 6876 1826 6888
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 6733 6919 6791 6925
rect 5408 6888 6132 6916
rect 5408 6876 5414 6888
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2958 6848 2964 6860
rect 2740 6820 2964 6848
rect 2740 6808 2746 6820
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 6104 6857 6132 6888
rect 6733 6885 6745 6919
rect 6779 6916 6791 6919
rect 6822 6916 6828 6928
rect 6779 6888 6828 6916
rect 6779 6885 6791 6888
rect 6733 6879 6791 6885
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 10686 6916 10692 6928
rect 10647 6888 10692 6916
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 11238 6916 11244 6928
rect 11199 6888 11244 6916
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 5224 6820 5273 6848
rect 5224 6808 5230 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 5261 6811 5319 6817
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6817 6055 6851
rect 5997 6811 6055 6817
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6817 6147 6851
rect 6454 6848 6460 6860
rect 6415 6820 6460 6848
rect 6089 6811 6147 6817
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2832 6752 3065 6780
rect 2832 6740 2838 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 4246 6780 4252 6792
rect 4207 6752 4252 6780
rect 3053 6743 3111 6749
rect 3068 6712 3096 6743
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 6012 6780 6040 6811
rect 6454 6808 6460 6820
rect 6512 6848 6518 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6512 6820 7021 6848
rect 6512 6808 6518 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 11388 6820 12081 6848
rect 11388 6808 11394 6820
rect 12069 6817 12081 6820
rect 12115 6817 12127 6851
rect 12342 6848 12348 6860
rect 12303 6820 12348 6848
rect 12069 6811 12127 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 13722 6848 13728 6860
rect 13679 6820 13728 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 6178 6780 6184 6792
rect 6012 6752 6184 6780
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 6788 6752 7573 6780
rect 6788 6740 6794 6752
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 7607 6752 8769 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 10594 6780 10600 6792
rect 10555 6752 10600 6780
rect 8757 6743 8815 6749
rect 10594 6740 10600 6752
rect 10652 6780 10658 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 10652 6752 11897 6780
rect 10652 6740 10658 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 3068 6684 4936 6712
rect 3694 6644 3700 6656
rect 3655 6616 3700 6644
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 4908 6653 4936 6684
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 9861 6715 9919 6721
rect 9861 6712 9873 6715
rect 8168 6684 9873 6712
rect 8168 6672 8174 6684
rect 9861 6681 9873 6684
rect 9907 6681 9919 6715
rect 9861 6675 9919 6681
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 4982 6644 4988 6656
rect 4939 6616 4988 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 8662 6644 8668 6656
rect 8527 6616 8668 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 10042 6604 10048 6656
rect 10100 6644 10106 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 10100 6616 10241 6644
rect 10100 6604 10106 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11698 6644 11704 6656
rect 11655 6616 11704 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 1104 6554 20884 6576
rect 1104 6502 4648 6554
rect 4700 6502 4712 6554
rect 4764 6502 4776 6554
rect 4828 6502 4840 6554
rect 4892 6502 11982 6554
rect 12034 6502 12046 6554
rect 12098 6502 12110 6554
rect 12162 6502 12174 6554
rect 12226 6502 19315 6554
rect 19367 6502 19379 6554
rect 19431 6502 19443 6554
rect 19495 6502 19507 6554
rect 19559 6502 20884 6554
rect 1104 6480 20884 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1762 6440 1768 6452
rect 1719 6412 1768 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2556 6412 2697 6440
rect 2556 6400 2562 6412
rect 2685 6409 2697 6412
rect 2731 6440 2743 6443
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2731 6412 2789 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 5258 6440 5264 6452
rect 5219 6412 5264 6440
rect 2777 6403 2835 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 9033 6443 9091 6449
rect 6411 6412 8499 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 2516 6372 2544 6400
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 1780 6344 2544 6372
rect 4126 6344 6561 6372
rect 1780 6316 1808 6344
rect 1762 6304 1768 6316
rect 1675 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 3694 6304 3700 6316
rect 2372 6276 3700 6304
rect 2372 6264 2378 6276
rect 1544 6239 1602 6245
rect 1544 6205 1556 6239
rect 1590 6236 1602 6239
rect 1670 6236 1676 6248
rect 1590 6208 1676 6236
rect 1590 6205 1602 6208
rect 1544 6199 1602 6205
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 3436 6245 3464 6276
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 4126 6304 4154 6344
rect 6549 6341 6561 6344
rect 6595 6372 6607 6375
rect 8018 6372 8024 6384
rect 6595 6344 8024 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 8471 6372 8499 6412
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9398 6440 9404 6452
rect 9079 6412 9404 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9398 6400 9404 6412
rect 9456 6440 9462 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 9456 6412 12173 6440
rect 9456 6400 9462 6412
rect 12161 6409 12173 6412
rect 12207 6440 12219 6443
rect 12342 6440 12348 6452
rect 12207 6412 12348 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 9214 6372 9220 6384
rect 8471 6344 9220 6372
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 3804 6276 4154 6304
rect 5859 6307 5917 6313
rect 3804 6245 3832 6276
rect 5859 6273 5871 6307
rect 5905 6304 5917 6307
rect 9766 6304 9772 6316
rect 5905 6276 9772 6304
rect 5905 6273 5917 6276
rect 5859 6267 5917 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11020 6276 12449 6304
rect 11020 6264 11026 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 2731 6208 2973 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4798 6236 4804 6248
rect 4387 6208 4804 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 1394 6168 1400 6180
rect 1307 6140 1400 6168
rect 1394 6128 1400 6140
rect 1452 6168 1458 6180
rect 2130 6168 2136 6180
rect 1452 6140 2136 6168
rect 1452 6128 1458 6140
rect 2130 6128 2136 6140
rect 2188 6128 2194 6180
rect 2498 6128 2504 6180
rect 2556 6168 2562 6180
rect 3804 6168 3832 6199
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5772 6239 5830 6245
rect 5772 6205 5784 6239
rect 5818 6236 5830 6239
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 5818 6208 6377 6236
rect 5818 6205 5830 6208
rect 5772 6199 5830 6205
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 6365 6199 6423 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 7374 6236 7380 6248
rect 6871 6208 7380 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8110 6236 8116 6248
rect 8071 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 8255 6208 9873 6236
rect 2556 6140 3832 6168
rect 4433 6171 4491 6177
rect 2556 6128 2562 6140
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 8255 6168 8283 6208
rect 9861 6205 9873 6208
rect 9907 6236 9919 6239
rect 10042 6236 10048 6248
rect 9907 6208 10048 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10744 6208 10793 6236
rect 10744 6196 10750 6208
rect 10781 6205 10793 6208
rect 10827 6236 10839 6239
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 10827 6208 11161 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 11149 6205 11161 6208
rect 11195 6236 11207 6239
rect 12526 6236 12532 6248
rect 11195 6208 12532 6236
rect 11195 6205 11207 6208
rect 11149 6199 11207 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 4479 6140 8283 6168
rect 8454 6171 8512 6177
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 8454 6137 8466 6171
rect 8500 6168 8512 6171
rect 8754 6168 8760 6180
rect 8500 6140 8760 6168
rect 8500 6137 8512 6140
rect 8454 6131 8512 6137
rect 8754 6128 8760 6140
rect 8812 6168 8818 6180
rect 9309 6171 9367 6177
rect 9309 6168 9321 6171
rect 8812 6140 9321 6168
rect 8812 6128 8818 6140
rect 9309 6137 9321 6140
rect 9355 6168 9367 6171
rect 9677 6171 9735 6177
rect 9677 6168 9689 6171
rect 9355 6140 9689 6168
rect 9355 6137 9367 6140
rect 9309 6131 9367 6137
rect 9677 6137 9689 6140
rect 9723 6168 9735 6171
rect 10182 6171 10240 6177
rect 10182 6168 10194 6171
rect 9723 6140 10194 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10182 6137 10194 6140
rect 10228 6137 10240 6171
rect 10182 6131 10240 6137
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 2958 6100 2964 6112
rect 2455 6072 2964 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 2958 6060 2964 6072
rect 3016 6100 3022 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 3016 6072 4905 6100
rect 3016 6060 3022 6072
rect 4893 6069 4905 6072
rect 4939 6100 4951 6103
rect 5166 6100 5172 6112
rect 4939 6072 5172 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 6178 6100 6184 6112
rect 6139 6072 6184 6100
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7006 6100 7012 6112
rect 6967 6072 7012 6100
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7892 6072 7941 6100
rect 7892 6060 7898 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 11422 6100 11428 6112
rect 11383 6072 11428 6100
rect 7929 6063 7987 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 13722 6100 13728 6112
rect 13683 6072 13728 6100
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 1104 6010 20884 6032
rect 1104 5958 8315 6010
rect 8367 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 15648 6010
rect 15700 5958 15712 6010
rect 15764 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 20884 6010
rect 1104 5936 20884 5958
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 2648 5868 3801 5896
rect 2648 5856 2654 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 4246 5856 4252 5908
rect 4304 5896 4310 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 4304 5868 8585 5896
rect 4304 5856 4310 5868
rect 3513 5831 3571 5837
rect 3513 5797 3525 5831
rect 3559 5828 3571 5831
rect 4798 5828 4804 5840
rect 3559 5800 4804 5828
rect 3559 5797 3571 5800
rect 3513 5791 3571 5797
rect 3804 5772 3832 5800
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 6178 5828 6184 5840
rect 5132 5800 6184 5828
rect 5132 5788 5138 5800
rect 1762 5760 1768 5772
rect 1723 5732 1768 5760
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2314 5760 2320 5772
rect 2275 5732 2320 5760
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 2648 5732 3065 5760
rect 2648 5720 2654 5732
rect 3053 5729 3065 5732
rect 3099 5760 3111 5763
rect 3602 5760 3608 5772
rect 3099 5732 3608 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3602 5720 3608 5732
rect 3660 5720 3666 5772
rect 3786 5720 3792 5772
rect 3844 5720 3850 5772
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 5736 5769 5764 5800
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 6730 5828 6736 5840
rect 6691 5800 6736 5828
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 7668 5837 7696 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 10226 5896 10232 5908
rect 8573 5859 8631 5865
rect 9968 5868 10232 5896
rect 7653 5831 7711 5837
rect 7653 5797 7665 5831
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 7745 5831 7803 5837
rect 7745 5797 7757 5831
rect 7791 5828 7803 5831
rect 8662 5828 8668 5840
rect 7791 5800 8668 5828
rect 7791 5797 7803 5800
rect 7745 5791 7803 5797
rect 8662 5788 8668 5800
rect 8720 5828 8726 5840
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8720 5800 8953 5828
rect 8720 5788 8726 5800
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9968 5837 9996 5868
rect 10226 5856 10232 5868
rect 10284 5896 10290 5908
rect 11330 5896 11336 5908
rect 10284 5868 11336 5896
rect 10284 5856 10290 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12526 5896 12532 5908
rect 12487 5868 12532 5896
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13035 5899 13093 5905
rect 13035 5896 13047 5899
rect 12952 5868 13047 5896
rect 12952 5856 12958 5868
rect 13035 5865 13047 5868
rect 13081 5865 13093 5899
rect 13035 5859 13093 5865
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 9732 5800 9873 5828
rect 9732 5788 9738 5800
rect 9861 5797 9873 5800
rect 9907 5797 9919 5831
rect 9861 5791 9919 5797
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5797 10011 5831
rect 9953 5791 10011 5797
rect 10505 5831 10563 5837
rect 10505 5797 10517 5831
rect 10551 5828 10563 5831
rect 10594 5828 10600 5840
rect 10551 5800 10600 5828
rect 10551 5797 10563 5800
rect 10505 5791 10563 5797
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 11517 5831 11575 5837
rect 11517 5797 11529 5831
rect 11563 5828 11575 5831
rect 11606 5828 11612 5840
rect 11563 5800 11612 5828
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 5224 5732 5273 5760
rect 5224 5720 5230 5732
rect 5261 5729 5273 5732
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5729 5779 5763
rect 6270 5760 6276 5772
rect 6231 5732 6276 5760
rect 5721 5723 5779 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6454 5720 6460 5732
rect 6512 5760 6518 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 6512 5732 7389 5760
rect 6512 5720 6518 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12894 5760 12900 5772
rect 12952 5769 12958 5772
rect 12952 5763 12990 5769
rect 12492 5732 12900 5760
rect 12492 5720 12498 5732
rect 12894 5720 12900 5732
rect 12978 5729 12990 5763
rect 12952 5723 12990 5729
rect 12952 5720 12958 5723
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 7190 5692 7196 5704
rect 4295 5664 7196 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 10962 5692 10968 5704
rect 10919 5664 10968 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11422 5692 11428 5704
rect 11383 5664 11428 5692
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13786 5664 13921 5692
rect 3053 5627 3111 5633
rect 3053 5593 3065 5627
rect 3099 5624 3111 5627
rect 8110 5624 8116 5636
rect 3099 5596 8116 5624
rect 3099 5593 3111 5596
rect 3053 5587 3111 5593
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 5074 5556 5080 5568
rect 5035 5528 5080 5556
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 7098 5556 7104 5568
rect 7059 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 9306 5556 9312 5568
rect 9267 5528 9312 5556
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 10376 5528 11161 5556
rect 10376 5516 10382 5528
rect 11149 5525 11161 5528
rect 11195 5525 11207 5559
rect 11149 5519 11207 5525
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 13786 5556 13814 5664
rect 13909 5661 13921 5664
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 11848 5528 13814 5556
rect 11848 5516 11854 5528
rect 1104 5466 20884 5488
rect 1104 5414 4648 5466
rect 4700 5414 4712 5466
rect 4764 5414 4776 5466
rect 4828 5414 4840 5466
rect 4892 5414 11982 5466
rect 12034 5414 12046 5466
rect 12098 5414 12110 5466
rect 12162 5414 12174 5466
rect 12226 5414 19315 5466
rect 19367 5414 19379 5466
rect 19431 5414 19443 5466
rect 19495 5414 19507 5466
rect 19559 5414 20884 5466
rect 1104 5392 20884 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2590 5352 2596 5364
rect 2455 5324 2596 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 3660 5324 4261 5352
rect 3660 5312 3666 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 8018 5352 8024 5364
rect 7979 5324 8024 5352
rect 4249 5315 4307 5321
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2498 5216 2504 5228
rect 2087 5188 2504 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 4264 5216 4292 5315
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8754 5352 8760 5364
rect 8715 5324 8760 5352
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10226 5352 10232 5364
rect 10187 5324 10232 5352
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 14139 5355 14197 5361
rect 14139 5352 14151 5355
rect 11480 5324 14151 5352
rect 11480 5312 11486 5324
rect 14139 5321 14151 5324
rect 14185 5321 14197 5355
rect 14139 5315 14197 5321
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 6730 5284 6736 5296
rect 5859 5256 6736 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 6730 5244 6736 5256
rect 6788 5284 6794 5296
rect 9306 5284 9312 5296
rect 6788 5256 9312 5284
rect 6788 5244 6794 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 9732 5256 13829 5284
rect 9732 5244 9738 5256
rect 13817 5253 13829 5256
rect 13863 5253 13875 5287
rect 13817 5247 13875 5253
rect 4338 5216 4344 5228
rect 4251 5188 4344 5216
rect 4338 5176 4344 5188
rect 4396 5216 4402 5228
rect 4396 5188 5304 5216
rect 4396 5176 4402 5188
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1489 5151 1547 5157
rect 1489 5148 1501 5151
rect 1452 5120 1501 5148
rect 1452 5108 1458 5120
rect 1489 5117 1501 5120
rect 1535 5117 1547 5151
rect 1670 5148 1676 5160
rect 1631 5120 1676 5148
rect 1489 5111 1547 5117
rect 1670 5108 1676 5120
rect 1728 5108 1734 5160
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2700 5120 2973 5148
rect 2130 4972 2136 5024
rect 2188 5012 2194 5024
rect 2700 5021 2728 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5117 4491 5151
rect 4890 5148 4896 5160
rect 4851 5120 4896 5148
rect 4433 5111 4491 5117
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5080 3663 5083
rect 4246 5080 4252 5092
rect 3651 5052 4252 5080
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 2188 4984 2697 5012
rect 2188 4972 2194 4984
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 2685 4975 2743 4981
rect 3973 5015 4031 5021
rect 3973 4981 3985 5015
rect 4019 5012 4031 5015
rect 4448 5012 4476 5111
rect 4890 5108 4896 5120
rect 4948 5148 4954 5160
rect 5074 5148 5080 5160
rect 4948 5120 5080 5148
rect 4948 5108 4954 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5276 5157 5304 5188
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6696 5188 6837 5216
rect 6696 5176 6702 5188
rect 6825 5185 6837 5188
rect 6871 5216 6883 5219
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 6871 5188 10517 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11146 5216 11152 5228
rect 10919 5188 11152 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11146 5176 11152 5188
rect 11204 5216 11210 5228
rect 11698 5216 11704 5228
rect 11204 5188 11704 5216
rect 11204 5176 11210 5188
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13354 5216 13360 5228
rect 12952 5188 13360 5216
rect 12952 5176 12958 5188
rect 13354 5176 13360 5188
rect 13412 5216 13418 5228
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 13412 5188 13461 5216
rect 13412 5176 13418 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 13538 5176 13544 5228
rect 13596 5216 13602 5228
rect 13596 5188 13814 5216
rect 13596 5176 13602 5188
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5442 5148 5448 5160
rect 5307 5120 5448 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6362 5148 6368 5160
rect 5859 5120 6368 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8260 5120 8953 5148
rect 8260 5108 8266 5120
rect 8941 5117 8953 5120
rect 8987 5148 8999 5151
rect 9122 5148 9128 5160
rect 8987 5120 9128 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 12529 5151 12587 5157
rect 12529 5117 12541 5151
rect 12575 5117 12587 5151
rect 13786 5148 13814 5188
rect 14068 5151 14126 5157
rect 14068 5148 14080 5151
rect 13786 5120 14080 5148
rect 12529 5111 12587 5117
rect 14068 5117 14080 5120
rect 14114 5148 14126 5151
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14114 5120 14473 5148
rect 14114 5117 14126 5120
rect 14068 5111 14126 5117
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 7146 5083 7204 5089
rect 7146 5049 7158 5083
rect 7192 5080 7204 5083
rect 7834 5080 7840 5092
rect 7192 5052 7840 5080
rect 7192 5049 7204 5052
rect 7146 5043 7204 5049
rect 5166 5012 5172 5024
rect 4019 4984 5172 5012
rect 4019 4981 4031 4984
rect 3973 4975 4031 4981
rect 5166 4972 5172 4984
rect 5224 5012 5230 5024
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 5224 4984 6193 5012
rect 5224 4972 5230 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6181 4975 6239 4981
rect 6546 4972 6552 4984
rect 6604 5012 6610 5024
rect 7161 5012 7189 5043
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 8754 5040 8760 5092
rect 8812 5080 8818 5092
rect 9262 5083 9320 5089
rect 9262 5080 9274 5083
rect 8812 5052 9274 5080
rect 8812 5040 8818 5052
rect 9262 5049 9274 5052
rect 9308 5080 9320 5083
rect 9674 5080 9680 5092
rect 9308 5052 9680 5080
rect 9308 5049 9320 5052
rect 9262 5043 9320 5049
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 10962 5080 10968 5092
rect 9876 5052 10968 5080
rect 7742 5012 7748 5024
rect 6604 4984 7189 5012
rect 7703 4984 7748 5012
rect 6604 4972 6610 4984
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 9876 5021 9904 5052
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 11974 5080 11980 5092
rect 11563 5052 11980 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 12434 5080 12440 5092
rect 12395 5052 12440 5080
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8168 4984 8401 5012
rect 8168 4972 8174 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8389 4975 8447 4981
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 4981 9919 5015
rect 9861 4975 9919 4981
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 11606 5012 11612 5024
rect 10652 4984 11612 5012
rect 10652 4972 10658 4984
rect 11606 4972 11612 4984
rect 11664 5012 11670 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11664 4984 11805 5012
rect 11664 4972 11670 4984
rect 11793 4981 11805 4984
rect 11839 5012 11851 5015
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11839 4984 12173 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12161 4981 12173 4984
rect 12207 5012 12219 5015
rect 12544 5012 12572 5111
rect 12207 4984 12572 5012
rect 12207 4981 12219 4984
rect 12161 4975 12219 4981
rect 1104 4922 20884 4944
rect 1104 4870 8315 4922
rect 8367 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 15648 4922
rect 15700 4870 15712 4922
rect 15764 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 20884 4922
rect 1104 4848 20884 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1820 4780 1961 4808
rect 1820 4768 1826 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 1949 4771 2007 4777
rect 3697 4811 3755 4817
rect 3697 4777 3709 4811
rect 3743 4808 3755 4811
rect 3786 4808 3792 4820
rect 3743 4780 3792 4808
rect 3743 4777 3755 4780
rect 3697 4771 3755 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4304 4780 4629 4808
rect 4304 4768 4310 4780
rect 4617 4777 4629 4780
rect 4663 4808 4675 4811
rect 4890 4808 4896 4820
rect 4663 4780 4896 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7156 4780 7297 4808
rect 7156 4768 7162 4780
rect 7285 4777 7297 4780
rect 7331 4808 7343 4811
rect 7834 4808 7840 4820
rect 7331 4780 7840 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 8128 4780 10885 4808
rect 1394 4700 1400 4752
rect 1452 4740 1458 4752
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 1452 4712 2329 4740
rect 1452 4700 1458 4712
rect 2317 4709 2329 4712
rect 2363 4740 2375 4743
rect 2406 4740 2412 4752
rect 2363 4712 2412 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 3804 4740 3832 4768
rect 4908 4740 4936 4768
rect 6638 4740 6644 4752
rect 3804 4712 4568 4740
rect 4908 4712 5672 4740
rect 6599 4712 6644 4740
rect 4062 4672 4068 4684
rect 2479 4644 3924 4672
rect 4023 4644 4068 4672
rect 1946 4564 1952 4616
rect 2004 4604 2010 4616
rect 2479 4613 2507 4644
rect 2464 4607 2522 4613
rect 2464 4604 2476 4607
rect 2004 4576 2476 4604
rect 2004 4564 2010 4576
rect 2464 4573 2476 4576
rect 2510 4573 2522 4607
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2464 4567 2522 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 3896 4604 3924 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4540 4672 4568 4712
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4540 4644 4997 4672
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 4985 4635 5043 4641
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 3896 4576 4905 4604
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 5000 4604 5028 4635
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5644 4681 5672 4712
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 7558 4740 7564 4752
rect 7248 4712 7564 4740
rect 7248 4700 7254 4712
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 7653 4743 7711 4749
rect 7653 4709 7665 4743
rect 7699 4740 7711 4743
rect 7742 4740 7748 4752
rect 7699 4712 7748 4740
rect 7699 4709 7711 4712
rect 7653 4703 7711 4709
rect 7742 4700 7748 4712
rect 7800 4740 7806 4752
rect 8128 4740 8156 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 11388 4780 13277 4808
rect 11388 4768 11394 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 7800 4712 8156 4740
rect 8205 4743 8263 4749
rect 7800 4700 7806 4712
rect 8205 4709 8217 4743
rect 8251 4740 8263 4743
rect 8297 4743 8355 4749
rect 8297 4740 8309 4743
rect 8251 4712 8309 4740
rect 8251 4709 8263 4712
rect 8205 4703 8263 4709
rect 8297 4709 8309 4712
rect 8343 4740 8355 4743
rect 9214 4740 9220 4752
rect 8343 4712 9220 4740
rect 8343 4709 8355 4712
rect 8297 4703 8355 4709
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 9998 4743 10056 4749
rect 9998 4740 10010 4743
rect 9732 4712 10010 4740
rect 9732 4700 9738 4712
rect 9998 4709 10010 4712
rect 10044 4709 10056 4743
rect 11790 4740 11796 4752
rect 11751 4712 11796 4740
rect 9998 4703 10056 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 5902 4672 5908 4684
rect 5675 4644 5908 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 5997 4635 6055 4641
rect 5718 4604 5724 4616
rect 5000 4576 5724 4604
rect 4893 4567 4951 4573
rect 5718 4564 5724 4576
rect 5776 4604 5782 4616
rect 6012 4604 6040 4635
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 5776 4576 6040 4604
rect 5776 4564 5782 4576
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 7616 4576 8861 4604
rect 7616 4564 7622 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 11330 4604 11336 4616
rect 9723 4576 11336 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11698 4604 11704 4616
rect 11659 4576 11704 4604
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 1854 4496 1860 4548
rect 1912 4536 1918 4548
rect 2314 4536 2320 4548
rect 1912 4508 2320 4536
rect 1912 4496 1918 4508
rect 2314 4496 2320 4508
rect 2372 4536 2378 4548
rect 2593 4539 2651 4545
rect 2593 4536 2605 4539
rect 2372 4508 2605 4536
rect 2372 4496 2378 4508
rect 2593 4505 2605 4508
rect 2639 4505 2651 4539
rect 2593 4499 2651 4505
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 4430 4536 4436 4548
rect 3007 4508 4436 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 4430 4496 4436 4508
rect 4488 4536 4494 4548
rect 4488 4508 7052 4536
rect 4488 4496 4494 4508
rect 4295 4471 4353 4477
rect 4295 4437 4307 4471
rect 4341 4468 4353 4471
rect 4522 4468 4528 4480
rect 4341 4440 4528 4468
rect 4341 4437 4353 4440
rect 4295 4431 4353 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 6822 4468 6828 4480
rect 4939 4440 6828 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 6822 4428 6828 4440
rect 6880 4468 6886 4480
rect 6917 4471 6975 4477
rect 6917 4468 6929 4471
rect 6880 4440 6929 4468
rect 6880 4428 6886 4440
rect 6917 4437 6929 4440
rect 6963 4437 6975 4471
rect 7024 4468 7052 4508
rect 8018 4496 8024 4548
rect 8076 4536 8082 4548
rect 8297 4539 8355 4545
rect 8297 4536 8309 4539
rect 8076 4508 8309 4536
rect 8076 4496 8082 4508
rect 8297 4505 8309 4508
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9217 4539 9275 4545
rect 9217 4536 9229 4539
rect 8812 4508 9229 4536
rect 8812 4496 8818 4508
rect 9217 4505 9229 4508
rect 9263 4505 9275 4539
rect 11992 4536 12020 4564
rect 13814 4536 13820 4548
rect 11992 4508 13820 4536
rect 9217 4499 9275 4505
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 8570 4468 8576 4480
rect 7024 4440 8576 4468
rect 6917 4431 6975 4437
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 11238 4468 11244 4480
rect 11199 4440 11244 4468
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 11480 4440 12633 4468
rect 11480 4428 11486 4440
rect 12621 4437 12633 4440
rect 12667 4437 12679 4471
rect 12986 4468 12992 4480
rect 12947 4440 12992 4468
rect 12621 4431 12679 4437
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 1104 4378 20884 4400
rect 1104 4326 4648 4378
rect 4700 4326 4712 4378
rect 4764 4326 4776 4378
rect 4828 4326 4840 4378
rect 4892 4326 11982 4378
rect 12034 4326 12046 4378
rect 12098 4326 12110 4378
rect 12162 4326 12174 4378
rect 12226 4326 19315 4378
rect 19367 4326 19379 4378
rect 19431 4326 19443 4378
rect 19495 4326 19507 4378
rect 19559 4326 20884 4378
rect 1104 4304 20884 4326
rect 1946 4224 1952 4276
rect 2004 4264 2010 4276
rect 2179 4267 2237 4273
rect 2179 4264 2191 4267
rect 2004 4236 2191 4264
rect 2004 4224 2010 4236
rect 2179 4233 2191 4236
rect 2225 4233 2237 4267
rect 2314 4264 2320 4276
rect 2275 4236 2320 4264
rect 2179 4227 2237 4233
rect 2314 4224 2320 4236
rect 2372 4264 2378 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 2372 4236 3065 4264
rect 2372 4224 2378 4236
rect 3053 4233 3065 4236
rect 3099 4264 3111 4267
rect 3421 4267 3479 4273
rect 3421 4264 3433 4267
rect 3099 4236 3433 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3421 4233 3433 4236
rect 3467 4233 3479 4267
rect 3421 4227 3479 4233
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 5960 4236 6193 4264
rect 5960 4224 5966 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 6181 4227 6239 4233
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 12526 4264 12532 4276
rect 11020 4236 12532 4264
rect 11020 4224 11026 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 13446 4264 13452 4276
rect 13228 4236 13452 4264
rect 13228 4224 13234 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 13817 4267 13875 4273
rect 13817 4264 13829 4267
rect 13688 4236 13829 4264
rect 13688 4224 13694 4236
rect 13817 4233 13829 4236
rect 13863 4233 13875 4267
rect 13817 4227 13875 4233
rect 4433 4199 4491 4205
rect 4433 4165 4445 4199
rect 4479 4196 4491 4199
rect 8202 4196 8208 4208
rect 4479 4168 8208 4196
rect 4479 4165 4491 4168
rect 4433 4159 4491 4165
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 11146 4196 11152 4208
rect 11107 4168 11152 4196
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 12986 4196 12992 4208
rect 11348 4168 12992 4196
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1912 4100 2421 4128
rect 1912 4088 1918 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 2866 4128 2872 4140
rect 2823 4100 2872 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 3016 4100 5273 4128
rect 3016 4088 3022 4100
rect 5261 4097 5273 4100
rect 5307 4128 5319 4131
rect 5307 4100 5948 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 3786 4060 3792 4072
rect 3747 4032 3792 4060
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4430 4060 4436 4072
rect 4203 4032 4436 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 5920 4060 5948 4100
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6788 4100 6837 4128
rect 6788 4088 6794 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 8938 4128 8944 4140
rect 8720 4100 8765 4128
rect 8899 4100 8944 4128
rect 8720 4088 8726 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 11348 4128 11376 4168
rect 12986 4156 12992 4168
rect 13044 4156 13050 4208
rect 10643 4100 11376 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11940 4100 11989 4128
rect 11940 4088 11946 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12526 4060 12532 4072
rect 5920 4032 8524 4060
rect 12487 4032 12532 4060
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 2406 3992 2412 4004
rect 2087 3964 2412 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 2406 3952 2412 3964
rect 2464 3952 2470 4004
rect 4706 3992 4712 4004
rect 4126 3964 4712 3992
rect 4126 3936 4154 3964
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5902 3992 5908 4004
rect 5408 3964 5453 3992
rect 5863 3964 5908 3992
rect 5408 3952 5414 3964
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7146 3995 7204 4001
rect 7146 3992 7158 3995
rect 6564 3964 7158 3992
rect 6564 3936 6592 3964
rect 7146 3961 7158 3964
rect 7192 3961 7204 3995
rect 7146 3955 7204 3961
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 3970 3924 3976 3936
rect 2004 3896 3976 3924
rect 2004 3884 2010 3896
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4062 3884 4068 3936
rect 4120 3896 4154 3936
rect 4120 3884 4126 3896
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 4985 3927 5043 3933
rect 4985 3924 4997 3927
rect 4580 3896 4997 3924
rect 4580 3884 4586 3896
rect 4985 3893 4997 3896
rect 5031 3924 5043 3927
rect 5166 3924 5172 3936
rect 5031 3896 5172 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 7834 3884 7840 3936
rect 7892 3924 7898 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 7892 3896 8033 3924
rect 7892 3884 7898 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8168 3896 8401 3924
rect 8168 3884 8174 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8496 3924 8524 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14036 4063 14094 4069
rect 14036 4060 14048 4063
rect 13872 4032 14048 4060
rect 13872 4020 13878 4032
rect 14036 4029 14048 4032
rect 14082 4060 14094 4063
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 14082 4032 14473 4060
rect 14082 4029 14094 4032
rect 14036 4023 14094 4029
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 8754 3992 8760 4004
rect 8715 3964 8760 3992
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 10318 3992 10324 4004
rect 8864 3964 10324 3992
rect 8864 3924 8892 3964
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10459 3964 10701 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 10689 3961 10701 3964
rect 10735 3961 10747 3995
rect 10689 3955 10747 3961
rect 11701 3995 11759 4001
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 11790 3992 11796 4004
rect 11747 3964 11796 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 9674 3924 9680 3936
rect 8496 3896 8892 3924
rect 9635 3896 9680 3924
rect 8389 3887 8447 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10704 3924 10732 3955
rect 11790 3952 11796 3964
rect 11848 3992 11854 4004
rect 12437 3995 12495 4001
rect 12437 3992 12449 3995
rect 11848 3964 12449 3992
rect 11848 3952 11854 3964
rect 12437 3961 12449 3964
rect 12483 3961 12495 3995
rect 12437 3955 12495 3961
rect 12342 3924 12348 3936
rect 10704 3896 12348 3924
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 14139 3927 14197 3933
rect 14139 3893 14151 3927
rect 14185 3924 14197 3927
rect 20990 3924 20996 3936
rect 14185 3896 20996 3924
rect 14185 3893 14197 3896
rect 14139 3887 14197 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 1104 3834 20884 3856
rect 1104 3782 8315 3834
rect 8367 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 15648 3834
rect 15700 3782 15712 3834
rect 15764 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 20884 3834
rect 1104 3760 20884 3782
rect 1535 3723 1593 3729
rect 1535 3689 1547 3723
rect 1581 3720 1593 3723
rect 2958 3720 2964 3732
rect 1581 3692 2964 3720
rect 1581 3689 1593 3692
rect 1535 3683 1593 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3200 3692 3525 3720
rect 3200 3680 3206 3692
rect 3513 3689 3525 3692
rect 3559 3720 3571 3723
rect 3786 3720 3792 3732
rect 3559 3692 3792 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4154 3720 4160 3732
rect 4028 3692 4160 3720
rect 4028 3680 4034 3692
rect 4154 3680 4160 3692
rect 4212 3720 4218 3732
rect 5534 3720 5540 3732
rect 4212 3692 5540 3720
rect 4212 3680 4218 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7742 3720 7748 3732
rect 7484 3692 7748 3720
rect 2314 3612 2320 3664
rect 2372 3652 2378 3664
rect 2409 3655 2467 3661
rect 2409 3652 2421 3655
rect 2372 3624 2421 3652
rect 2372 3612 2378 3624
rect 2409 3621 2421 3624
rect 2455 3621 2467 3655
rect 2409 3615 2467 3621
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 7484 3661 7512 3692
rect 7742 3680 7748 3692
rect 7800 3720 7806 3732
rect 10962 3720 10968 3732
rect 7800 3692 10968 3720
rect 7800 3680 7806 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11330 3720 11336 3732
rect 11291 3692 11336 3720
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 12526 3720 12532 3732
rect 12487 3692 12532 3720
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 14001 3723 14059 3729
rect 14001 3720 14013 3723
rect 12768 3692 14013 3720
rect 12768 3680 12774 3692
rect 14001 3689 14013 3692
rect 14047 3689 14059 3723
rect 14001 3683 14059 3689
rect 6457 3655 6515 3661
rect 6457 3652 6469 3655
rect 2832 3624 6469 3652
rect 2832 3612 2838 3624
rect 6457 3621 6469 3624
rect 6503 3621 6515 3655
rect 6457 3615 6515 3621
rect 7469 3655 7527 3661
rect 7469 3621 7481 3655
rect 7515 3621 7527 3655
rect 7469 3615 7527 3621
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3652 8171 3655
rect 8754 3652 8760 3664
rect 8159 3624 8760 3652
rect 8159 3621 8171 3624
rect 8113 3615 8171 3621
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 9401 3655 9459 3661
rect 9401 3652 9413 3655
rect 8812 3624 9413 3652
rect 8812 3612 8818 3624
rect 9401 3621 9413 3624
rect 9447 3621 9459 3655
rect 10042 3652 10048 3664
rect 10003 3624 10048 3652
rect 9401 3615 9459 3621
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 11606 3652 11612 3664
rect 11567 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12676 3624 13001 3652
rect 12676 3612 12682 3624
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 1464 3587 1522 3593
rect 1464 3553 1476 3587
rect 1510 3584 1522 3587
rect 1946 3584 1952 3596
rect 1510 3556 1952 3584
rect 1510 3553 1522 3556
rect 1464 3547 1522 3553
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2556 3587 2614 3593
rect 2556 3553 2568 3587
rect 2602 3584 2614 3587
rect 2792 3584 2820 3612
rect 2602 3556 2820 3584
rect 3881 3587 3939 3593
rect 2602 3553 2614 3556
rect 2556 3547 2614 3553
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 4982 3584 4988 3596
rect 3927 3556 4988 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3553 5319 3587
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5261 3547 5319 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2777 3519 2835 3525
rect 2777 3516 2789 3519
rect 1728 3488 2789 3516
rect 1728 3476 1734 3488
rect 2777 3485 2789 3488
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4433 3451 4491 3457
rect 4433 3448 4445 3451
rect 3936 3420 4445 3448
rect 3936 3408 3942 3420
rect 4433 3417 4445 3420
rect 4479 3448 4491 3451
rect 5074 3448 5080 3460
rect 4479 3420 5080 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 5074 3408 5080 3420
rect 5132 3448 5138 3460
rect 5276 3448 5304 3547
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5810 3544 5816 3596
rect 5868 3584 5874 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5868 3556 5917 3584
rect 5868 3544 5874 3556
rect 5905 3553 5917 3556
rect 5951 3584 5963 3587
rect 6362 3584 6368 3596
rect 5951 3556 6368 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 8260 3556 8309 3584
rect 8260 3544 8266 3556
rect 8297 3553 8309 3556
rect 8343 3584 8355 3587
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 8343 3556 8677 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 13538 3584 13544 3596
rect 13228 3556 13544 3584
rect 13228 3544 13234 3556
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 15194 3584 15200 3596
rect 15155 3556 15200 3584
rect 15194 3544 15200 3556
rect 15252 3544 15258 3596
rect 6178 3516 6184 3528
rect 6139 3488 6184 3516
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7650 3516 7656 3528
rect 7611 3488 7656 3516
rect 7377 3479 7435 3485
rect 5132 3420 5304 3448
rect 5132 3408 5138 3420
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 7392 3448 7420 3479
rect 7650 3476 7656 3488
rect 7708 3516 7714 3528
rect 8018 3516 8024 3528
rect 7708 3488 8024 3516
rect 7708 3476 7714 3488
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 9953 3519 10011 3525
rect 8128 3488 9812 3516
rect 8128 3448 8156 3488
rect 5960 3420 8156 3448
rect 5960 3408 5966 3420
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 9033 3451 9091 3457
rect 9033 3448 9045 3451
rect 8260 3420 9045 3448
rect 8260 3408 8266 3420
rect 9033 3417 9045 3420
rect 9079 3417 9091 3451
rect 9784 3448 9812 3488
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 11517 3519 11575 3525
rect 9999 3488 11376 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10502 3448 10508 3460
rect 9784 3420 10508 3448
rect 9033 3411 9091 3417
rect 10502 3408 10508 3420
rect 10560 3448 10566 3460
rect 11238 3448 11244 3460
rect 10560 3420 11244 3448
rect 10560 3408 10566 3420
rect 11238 3408 11244 3420
rect 11296 3408 11302 3460
rect 2130 3380 2136 3392
rect 2091 3352 2136 3380
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 3326 3380 3332 3392
rect 3099 3352 3332 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 5350 3380 5356 3392
rect 4212 3352 5356 3380
rect 4212 3340 4218 3352
rect 5350 3340 5356 3352
rect 5408 3380 5414 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 5408 3352 8125 3380
rect 5408 3340 5414 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8113 3343 8171 3349
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10836 3352 10885 3380
rect 10836 3340 10842 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 11348 3380 11376 3488
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 13998 3516 14004 3528
rect 11563 3488 14004 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 12069 3451 12127 3457
rect 12069 3448 12081 3451
rect 11848 3420 12081 3448
rect 11848 3408 11854 3420
rect 12069 3417 12081 3420
rect 12115 3448 12127 3451
rect 12618 3448 12624 3460
rect 12115 3420 12624 3448
rect 12115 3417 12127 3420
rect 12069 3411 12127 3417
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 13630 3448 13636 3460
rect 12728 3420 13636 3448
rect 12728 3380 12756 3420
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 15427 3451 15485 3457
rect 15427 3448 15439 3451
rect 13786 3420 15439 3448
rect 11348 3352 12756 3380
rect 10873 3343 10931 3349
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 12860 3352 12905 3380
rect 12860 3340 12866 3352
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 13786 3380 13814 3420
rect 15427 3417 15439 3420
rect 15473 3417 15485 3451
rect 15427 3411 15485 3417
rect 13412 3352 13814 3380
rect 13412 3340 13418 3352
rect 1104 3290 20884 3312
rect 1104 3238 4648 3290
rect 4700 3238 4712 3290
rect 4764 3238 4776 3290
rect 4828 3238 4840 3290
rect 4892 3238 11982 3290
rect 12034 3238 12046 3290
rect 12098 3238 12110 3290
rect 12162 3238 12174 3290
rect 12226 3238 19315 3290
rect 19367 3238 19379 3290
rect 19431 3238 19443 3290
rect 19495 3238 19507 3290
rect 19559 3238 20884 3290
rect 1104 3216 20884 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 4338 3176 4344 3188
rect 4299 3148 4344 3176
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5776 3148 6561 3176
rect 5776 3136 5782 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 8938 3176 8944 3188
rect 6972 3148 8944 3176
rect 6972 3136 6978 3148
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 10686 3176 10692 3188
rect 9180 3148 10692 3176
rect 9180 3136 9186 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 11057 3179 11115 3185
rect 11057 3176 11069 3179
rect 10928 3148 11069 3176
rect 10928 3136 10934 3148
rect 11057 3145 11069 3148
rect 11103 3176 11115 3179
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11103 3148 11529 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 11517 3145 11529 3148
rect 11563 3176 11575 3179
rect 11606 3176 11612 3188
rect 11563 3148 11612 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 13538 3176 13544 3188
rect 13499 3148 13544 3176
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13688 3148 14105 3176
rect 13688 3136 13694 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 14093 3139 14151 3145
rect 2130 3068 2136 3120
rect 2188 3108 2194 3120
rect 3878 3108 3884 3120
rect 2188 3080 3884 3108
rect 2188 3068 2194 3080
rect 2700 2981 2728 3080
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 4356 3040 4384 3136
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 9861 3111 9919 3117
rect 9861 3108 9873 3111
rect 5859 3080 9873 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 9861 3077 9873 3080
rect 9907 3077 9919 3111
rect 9861 3071 9919 3077
rect 9950 3068 9956 3120
rect 10008 3108 10014 3120
rect 12802 3108 12808 3120
rect 10008 3080 12808 3108
rect 10008 3068 10014 3080
rect 6914 3040 6920 3052
rect 4356 3012 5304 3040
rect 6875 3012 6920 3040
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2409 2975 2467 2981
rect 2409 2972 2421 2975
rect 2087 2944 2421 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2409 2941 2421 2944
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2941 2743 2975
rect 3142 2972 3148 2984
rect 3103 2944 3148 2972
rect 2685 2935 2743 2941
rect 2424 2836 2452 2935
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3326 2972 3332 2984
rect 3287 2944 3332 2972
rect 3326 2932 3332 2944
rect 3384 2972 3390 2984
rect 4709 2975 4767 2981
rect 3384 2944 4154 2972
rect 3384 2932 3390 2944
rect 3602 2904 3608 2916
rect 3563 2876 3608 2904
rect 3602 2864 3608 2876
rect 3660 2864 3666 2916
rect 3510 2836 3516 2848
rect 2424 2808 3516 2836
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4126 2836 4154 2944
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 4709 2935 4767 2941
rect 4724 2904 4752 2935
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5276 2981 5304 3012
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7650 3040 7656 3052
rect 7607 3012 7656 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7834 3040 7840 3052
rect 7795 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9324 3012 9689 3040
rect 5261 2975 5319 2981
rect 5261 2941 5273 2975
rect 5307 2972 5319 2975
rect 5350 2972 5356 2984
rect 5307 2944 5356 2972
rect 5307 2941 5319 2944
rect 5261 2935 5319 2941
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 9324 2981 9352 3012
rect 9677 3009 9689 3012
rect 9723 3040 9735 3043
rect 10042 3040 10048 3052
rect 9723 3012 10048 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 10042 3000 10048 3012
rect 10100 3040 10106 3052
rect 12544 3049 12572 3080
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 14737 3111 14795 3117
rect 14737 3077 14749 3111
rect 14783 3108 14795 3111
rect 15930 3108 15936 3120
rect 14783 3080 15936 3108
rect 14783 3077 14795 3080
rect 14737 3071 14795 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 12529 3043 12587 3049
rect 10100 3012 12296 3040
rect 10100 3000 10106 3012
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8260 2944 8401 2972
rect 8260 2932 8266 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2941 9367 2975
rect 9309 2935 9367 2941
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2972 9919 2975
rect 10137 2975 10195 2981
rect 10137 2972 10149 2975
rect 9907 2944 10149 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10137 2941 10149 2944
rect 10183 2972 10195 2975
rect 10778 2972 10784 2984
rect 10183 2944 10784 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11020 2944 11805 2972
rect 11020 2932 11026 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 4982 2904 4988 2916
rect 4724 2876 4988 2904
rect 4982 2864 4988 2876
rect 5040 2904 5046 2916
rect 6181 2907 6239 2913
rect 6181 2904 6193 2907
rect 5040 2876 6193 2904
rect 5040 2864 5046 2876
rect 6181 2873 6193 2876
rect 6227 2873 6239 2907
rect 6181 2867 6239 2873
rect 7009 2907 7067 2913
rect 7009 2873 7021 2907
rect 7055 2904 7067 2907
rect 7098 2904 7104 2916
rect 7055 2876 7104 2904
rect 7055 2873 7067 2876
rect 7009 2867 7067 2873
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7926 2864 7932 2916
rect 7984 2904 7990 2916
rect 8297 2907 8355 2913
rect 8297 2904 8309 2907
rect 7984 2876 8309 2904
rect 7984 2864 7990 2876
rect 8297 2873 8309 2876
rect 8343 2904 8355 2907
rect 8710 2907 8768 2913
rect 8710 2904 8722 2907
rect 8343 2876 8722 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 8710 2873 8722 2876
rect 8756 2904 8768 2907
rect 9674 2904 9680 2916
rect 8756 2876 9680 2904
rect 8756 2873 8768 2876
rect 8710 2867 8768 2873
rect 9674 2864 9680 2876
rect 9732 2904 9738 2916
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 9732 2876 9965 2904
rect 9732 2864 9738 2876
rect 9953 2873 9965 2876
rect 9999 2904 10011 2907
rect 10458 2907 10516 2913
rect 10458 2904 10470 2907
rect 9999 2876 10470 2904
rect 9999 2873 10011 2876
rect 9953 2867 10011 2873
rect 10458 2873 10470 2876
rect 10504 2873 10516 2907
rect 10458 2867 10516 2873
rect 5626 2836 5632 2848
rect 4126 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2836 5690 2848
rect 8110 2836 8116 2848
rect 5684 2808 8116 2836
rect 5684 2796 5690 2808
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 11238 2836 11244 2848
rect 8904 2808 11244 2836
rect 8904 2796 8910 2808
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 12268 2845 12296 3012
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12676 3012 12909 3040
rect 12676 3000 12682 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13044 3012 13814 3040
rect 13044 3000 13050 3012
rect 13786 2972 13814 3012
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 13786 2944 14565 2972
rect 14553 2941 14565 2944
rect 14599 2972 14611 2975
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14599 2944 15117 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15692 2975 15750 2981
rect 15692 2972 15704 2975
rect 15528 2944 15704 2972
rect 15528 2932 15534 2944
rect 15692 2941 15704 2944
rect 15738 2972 15750 2975
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15738 2944 16129 2972
rect 15738 2941 15750 2944
rect 15692 2935 15750 2941
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 16117 2935 16175 2941
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 14277 2907 14335 2913
rect 14277 2904 14289 2907
rect 14139 2876 14289 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 14277 2873 14289 2876
rect 14323 2904 14335 2907
rect 15795 2907 15853 2913
rect 15795 2904 15807 2907
rect 14323 2876 15807 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 15795 2873 15807 2876
rect 15841 2873 15853 2907
rect 15795 2867 15853 2873
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12636 2836 12664 2867
rect 12299 2808 12664 2836
rect 13909 2839 13967 2845
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 13998 2836 14004 2848
rect 13955 2808 14004 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 13998 2796 14004 2808
rect 14056 2796 14062 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 15194 2836 15200 2848
rect 14608 2808 15200 2836
rect 14608 2796 14614 2808
rect 15194 2796 15200 2808
rect 15252 2836 15258 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15252 2808 15485 2836
rect 15252 2796 15258 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 1104 2746 20884 2768
rect 1104 2694 8315 2746
rect 8367 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 15648 2746
rect 15700 2694 15712 2746
rect 15764 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 20884 2746
rect 1104 2672 20884 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1946 2632 1952 2644
rect 1719 2604 1952 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2314 2632 2320 2644
rect 2179 2604 2320 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2314 2592 2320 2604
rect 2372 2632 2378 2644
rect 3145 2635 3203 2641
rect 2372 2604 3096 2632
rect 2372 2592 2378 2604
rect 2222 2524 2228 2576
rect 2280 2564 2286 2576
rect 2546 2567 2604 2573
rect 2546 2564 2558 2567
rect 2280 2536 2558 2564
rect 2280 2524 2286 2536
rect 2546 2533 2558 2536
rect 2592 2533 2604 2567
rect 3068 2564 3096 2604
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 4154 2632 4160 2644
rect 3191 2604 4160 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 5905 2635 5963 2641
rect 5092 2604 5304 2632
rect 5092 2576 5120 2604
rect 4246 2564 4252 2576
rect 3068 2536 4252 2564
rect 2546 2527 2604 2533
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2561 2428 2589 2527
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 5074 2564 5080 2576
rect 5000 2536 5080 2564
rect 3697 2499 3755 2505
rect 3697 2465 3709 2499
rect 3743 2496 3755 2499
rect 4522 2496 4528 2508
rect 3743 2468 4528 2496
rect 3743 2465 3755 2468
rect 3697 2459 3755 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 5000 2505 5028 2536
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5276 2564 5304 2604
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 8202 2632 8208 2644
rect 5951 2604 8208 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8803 2635 8861 2641
rect 8803 2601 8815 2635
rect 8849 2632 8861 2635
rect 9858 2632 9864 2644
rect 8849 2604 9864 2632
rect 8849 2601 8861 2604
rect 8803 2595 8861 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10870 2632 10876 2644
rect 9968 2604 10876 2632
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 5276 2536 6285 2564
rect 6273 2533 6285 2536
rect 6319 2533 6331 2567
rect 6546 2564 6552 2576
rect 6459 2536 6552 2564
rect 6273 2527 6331 2533
rect 6546 2524 6552 2536
rect 6604 2564 6610 2576
rect 7238 2567 7296 2573
rect 7238 2564 7250 2567
rect 6604 2536 7250 2564
rect 6604 2524 6610 2536
rect 7238 2533 7250 2536
rect 7284 2564 7296 2567
rect 7926 2564 7932 2576
rect 7284 2536 7932 2564
rect 7284 2533 7296 2536
rect 7238 2527 7296 2533
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 8110 2564 8116 2576
rect 8071 2536 8116 2564
rect 8110 2524 8116 2536
rect 8168 2564 8174 2576
rect 9968 2573 9996 2604
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11330 2592 11336 2644
rect 11388 2632 11394 2644
rect 13909 2635 13967 2641
rect 13909 2632 13921 2635
rect 11388 2604 13921 2632
rect 11388 2592 11394 2604
rect 13909 2601 13921 2604
rect 13955 2601 13967 2635
rect 13909 2595 13967 2601
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 15611 2635 15669 2641
rect 15611 2632 15623 2635
rect 14056 2604 15623 2632
rect 14056 2592 14062 2604
rect 15611 2601 15623 2604
rect 15657 2601 15669 2635
rect 17126 2632 17132 2644
rect 17087 2604 17132 2632
rect 15611 2595 15669 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 8168 2536 8493 2564
rect 8168 2524 8174 2536
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 8481 2527 8539 2533
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10042 2524 10048 2576
rect 10100 2564 10106 2576
rect 13354 2564 13360 2576
rect 10100 2536 13360 2564
rect 10100 2524 10106 2536
rect 13354 2524 13360 2536
rect 13412 2564 13418 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 13412 2536 13553 2564
rect 13412 2524 13418 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2465 5043 2499
rect 5350 2496 5356 2508
rect 5311 2468 5356 2496
rect 4985 2459 5043 2465
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5684 2468 5733 2496
rect 5684 2456 5690 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 6914 2496 6920 2508
rect 6236 2468 6920 2496
rect 6236 2456 6242 2468
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7156 2468 7849 2496
rect 7156 2456 7162 2468
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 8732 2499 8790 2505
rect 8732 2465 8744 2499
rect 8778 2496 8790 2499
rect 9214 2496 9220 2508
rect 8778 2468 9220 2496
rect 8778 2465 8790 2468
rect 8732 2459 8790 2465
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 2561 2400 3433 2428
rect 2225 2391 2283 2397
rect 3421 2397 3433 2400
rect 3467 2428 3479 2431
rect 5442 2428 5448 2440
rect 3467 2400 5448 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 2240 2360 2268 2391
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 7852 2428 7880 2459
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 10560 2468 10605 2496
rect 10560 2456 10566 2468
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 10744 2468 11345 2496
rect 10744 2456 10750 2468
rect 11333 2465 11345 2468
rect 11379 2496 11391 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11379 2468 11897 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 11885 2459 11943 2465
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12667 2468 13185 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13713 2499 13771 2505
rect 13713 2465 13725 2499
rect 13759 2465 13771 2499
rect 13713 2459 13771 2465
rect 15540 2499 15598 2505
rect 15540 2465 15552 2499
rect 15586 2496 15598 2499
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15586 2468 16037 2496
rect 15586 2465 15598 2468
rect 15540 2459 15598 2465
rect 16025 2465 16037 2468
rect 16071 2496 16083 2499
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 16071 2468 16497 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16485 2465 16497 2468
rect 16531 2496 16543 2499
rect 17144 2496 17172 2592
rect 16531 2468 17172 2496
rect 16531 2465 16543 2468
rect 16485 2459 16543 2465
rect 9861 2431 9919 2437
rect 5828 2400 6868 2428
rect 7852 2400 9628 2428
rect 3602 2360 3608 2372
rect 2240 2332 3608 2360
rect 3602 2320 3608 2332
rect 3660 2360 3666 2372
rect 5828 2360 5856 2400
rect 3660 2332 5856 2360
rect 6840 2360 6868 2400
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 6840 2332 9505 2360
rect 3660 2320 3666 2332
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 9600 2360 9628 2400
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10042 2428 10048 2440
rect 9907 2400 10048 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10152 2400 11161 2428
rect 10152 2360 10180 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 12636 2428 12664 2459
rect 11296 2400 12664 2428
rect 11296 2388 11302 2400
rect 11517 2363 11575 2369
rect 11517 2360 11529 2363
rect 9600 2332 10180 2360
rect 10520 2332 11529 2360
rect 9493 2323 9551 2329
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3697 2295 3755 2301
rect 3697 2292 3709 2295
rect 3568 2264 3709 2292
rect 3568 2252 3574 2264
rect 3697 2261 3709 2264
rect 3743 2292 3755 2295
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3743 2264 3801 2292
rect 3743 2261 3755 2264
rect 3697 2255 3755 2261
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 5442 2252 5448 2304
rect 5500 2292 5506 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 5500 2264 6561 2292
rect 5500 2252 5506 2264
rect 6549 2261 6561 2264
rect 6595 2292 6607 2295
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6595 2264 6653 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 6641 2255 6699 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9582 2252 9588 2304
rect 9640 2292 9646 2304
rect 10520 2292 10548 2332
rect 11517 2329 11529 2332
rect 11563 2329 11575 2363
rect 13740 2360 13768 2459
rect 16669 2363 16727 2369
rect 13740 2332 14412 2360
rect 11517 2323 11575 2329
rect 12802 2292 12808 2304
rect 9640 2264 10548 2292
rect 12763 2264 12808 2292
rect 9640 2252 9646 2264
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 14384 2301 14412 2332
rect 16669 2329 16681 2363
rect 16715 2360 16727 2363
rect 17126 2360 17132 2372
rect 16715 2332 17132 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 14550 2292 14556 2304
rect 14415 2264 14556 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14550 2252 14556 2264
rect 14608 2252 14614 2304
rect 1104 2202 20884 2224
rect 1104 2150 4648 2202
rect 4700 2150 4712 2202
rect 4764 2150 4776 2202
rect 4828 2150 4840 2202
rect 4892 2150 11982 2202
rect 12034 2150 12046 2202
rect 12098 2150 12110 2202
rect 12162 2150 12174 2202
rect 12226 2150 19315 2202
rect 19367 2150 19379 2202
rect 19431 2150 19443 2202
rect 19495 2150 19507 2202
rect 19559 2150 20884 2202
rect 1104 2128 20884 2150
rect 9214 2048 9220 2100
rect 9272 2088 9278 2100
rect 11514 2088 11520 2100
rect 9272 2060 11520 2088
rect 9272 2048 9278 2060
rect 11514 2048 11520 2060
rect 11572 2048 11578 2100
rect 12618 2048 12624 2100
rect 12676 2088 12682 2100
rect 13078 2088 13084 2100
rect 12676 2060 13084 2088
rect 12676 2048 12682 2060
rect 13078 2048 13084 2060
rect 13136 2088 13142 2100
rect 15470 2088 15476 2100
rect 13136 2060 15476 2088
rect 13136 2048 13142 2060
rect 15470 2048 15476 2060
rect 15528 2048 15534 2100
rect 8386 76 8392 128
rect 8444 116 8450 128
rect 12802 116 12808 128
rect 8444 88 12808 116
rect 8444 76 8450 88
rect 12802 76 12808 88
rect 12860 76 12866 128
<< via1 >>
rect 20 21496 72 21548
rect 848 21496 900 21548
rect 1676 21496 1728 21548
rect 2504 21496 2556 21548
rect 8668 21496 8720 21548
rect 9220 21496 9272 21548
rect 9680 21496 9732 21548
rect 10968 21496 11020 21548
rect 15200 21496 15252 21548
rect 16028 21496 16080 21548
rect 16580 21496 16632 21548
rect 17684 21496 17736 21548
rect 19708 21496 19760 21548
rect 21088 21496 21140 21548
rect 4648 19558 4700 19610
rect 4712 19558 4764 19610
rect 4776 19558 4828 19610
rect 4840 19558 4892 19610
rect 11982 19558 12034 19610
rect 12046 19558 12098 19610
rect 12110 19558 12162 19610
rect 12174 19558 12226 19610
rect 19315 19558 19367 19610
rect 19379 19558 19431 19610
rect 19443 19558 19495 19610
rect 19507 19558 19559 19610
rect 8315 19014 8367 19066
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 15648 19014 15700 19066
rect 15712 19014 15764 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 4648 18470 4700 18522
rect 4712 18470 4764 18522
rect 4776 18470 4828 18522
rect 4840 18470 4892 18522
rect 11982 18470 12034 18522
rect 12046 18470 12098 18522
rect 12110 18470 12162 18522
rect 12174 18470 12226 18522
rect 19315 18470 19367 18522
rect 19379 18470 19431 18522
rect 19443 18470 19495 18522
rect 19507 18470 19559 18522
rect 6184 18411 6236 18420
rect 6184 18377 6193 18411
rect 6193 18377 6227 18411
rect 6227 18377 6236 18411
rect 6184 18368 6236 18377
rect 7380 18411 7432 18420
rect 7380 18377 7389 18411
rect 7389 18377 7423 18411
rect 7423 18377 7432 18411
rect 7380 18368 7432 18377
rect 14464 18368 14516 18420
rect 6184 18164 6236 18216
rect 5080 18028 5132 18080
rect 11796 18164 11848 18216
rect 8024 18028 8076 18080
rect 8315 17926 8367 17978
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 15648 17926 15700 17978
rect 15712 17926 15764 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 4160 17688 4212 17740
rect 4648 17382 4700 17434
rect 4712 17382 4764 17434
rect 4776 17382 4828 17434
rect 4840 17382 4892 17434
rect 11982 17382 12034 17434
rect 12046 17382 12098 17434
rect 12110 17382 12162 17434
rect 12174 17382 12226 17434
rect 19315 17382 19367 17434
rect 19379 17382 19431 17434
rect 19443 17382 19495 17434
rect 19507 17382 19559 17434
rect 19892 17280 19944 17332
rect 12348 17076 12400 17128
rect 4160 16940 4212 16992
rect 8315 16838 8367 16890
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 15648 16838 15700 16890
rect 15712 16838 15764 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 4648 16294 4700 16346
rect 4712 16294 4764 16346
rect 4776 16294 4828 16346
rect 4840 16294 4892 16346
rect 11982 16294 12034 16346
rect 12046 16294 12098 16346
rect 12110 16294 12162 16346
rect 12174 16294 12226 16346
rect 19315 16294 19367 16346
rect 19379 16294 19431 16346
rect 19443 16294 19495 16346
rect 19507 16294 19559 16346
rect 8315 15750 8367 15802
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 15648 15750 15700 15802
rect 15712 15750 15764 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 4648 15206 4700 15258
rect 4712 15206 4764 15258
rect 4776 15206 4828 15258
rect 4840 15206 4892 15258
rect 11982 15206 12034 15258
rect 12046 15206 12098 15258
rect 12110 15206 12162 15258
rect 12174 15206 12226 15258
rect 19315 15206 19367 15258
rect 19379 15206 19431 15258
rect 19443 15206 19495 15258
rect 19507 15206 19559 15258
rect 8315 14662 8367 14714
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 15648 14662 15700 14714
rect 15712 14662 15764 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 19064 14467 19116 14476
rect 19064 14433 19073 14467
rect 19073 14433 19107 14467
rect 19107 14433 19116 14467
rect 19064 14424 19116 14433
rect 19156 14220 19208 14272
rect 4648 14118 4700 14170
rect 4712 14118 4764 14170
rect 4776 14118 4828 14170
rect 4840 14118 4892 14170
rect 11982 14118 12034 14170
rect 12046 14118 12098 14170
rect 12110 14118 12162 14170
rect 12174 14118 12226 14170
rect 19315 14118 19367 14170
rect 19379 14118 19431 14170
rect 19443 14118 19495 14170
rect 19507 14118 19559 14170
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 8315 13574 8367 13626
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 15648 13574 15700 13626
rect 15712 13574 15764 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 4648 13030 4700 13082
rect 4712 13030 4764 13082
rect 4776 13030 4828 13082
rect 4840 13030 4892 13082
rect 11982 13030 12034 13082
rect 12046 13030 12098 13082
rect 12110 13030 12162 13082
rect 12174 13030 12226 13082
rect 19315 13030 19367 13082
rect 19379 13030 19431 13082
rect 19443 13030 19495 13082
rect 19507 13030 19559 13082
rect 8315 12486 8367 12538
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 15648 12486 15700 12538
rect 15712 12486 15764 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 4648 11942 4700 11994
rect 4712 11942 4764 11994
rect 4776 11942 4828 11994
rect 4840 11942 4892 11994
rect 11982 11942 12034 11994
rect 12046 11942 12098 11994
rect 12110 11942 12162 11994
rect 12174 11942 12226 11994
rect 19315 11942 19367 11994
rect 19379 11942 19431 11994
rect 19443 11942 19495 11994
rect 19507 11942 19559 11994
rect 1584 11815 1636 11824
rect 1584 11781 1593 11815
rect 1593 11781 1627 11815
rect 1627 11781 1636 11815
rect 1584 11772 1636 11781
rect 1308 11636 1360 11688
rect 2596 11636 2648 11688
rect 7104 11500 7156 11552
rect 9036 11500 9088 11552
rect 9680 11500 9732 11552
rect 8315 11398 8367 11450
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 15648 11398 15700 11450
rect 15712 11398 15764 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 7104 11339 7156 11348
rect 7104 11305 7113 11339
rect 7113 11305 7147 11339
rect 7147 11305 7156 11339
rect 7104 11296 7156 11305
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 2596 11203 2648 11212
rect 2596 11169 2605 11203
rect 2605 11169 2639 11203
rect 2639 11169 2648 11203
rect 2596 11160 2648 11169
rect 4252 11160 4304 11212
rect 5632 11160 5684 11212
rect 6644 11160 6696 11212
rect 7564 11160 7616 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 6276 11024 6328 11076
rect 7380 11024 7432 11076
rect 8668 11024 8720 11076
rect 3608 10956 3660 11008
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 6000 10956 6052 11008
rect 6552 10956 6604 11008
rect 9312 10956 9364 11008
rect 4648 10854 4700 10906
rect 4712 10854 4764 10906
rect 4776 10854 4828 10906
rect 4840 10854 4892 10906
rect 11982 10854 12034 10906
rect 12046 10854 12098 10906
rect 12110 10854 12162 10906
rect 12174 10854 12226 10906
rect 19315 10854 19367 10906
rect 19379 10854 19431 10906
rect 19443 10854 19495 10906
rect 19507 10854 19559 10906
rect 1400 10752 1452 10804
rect 2596 10752 2648 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 12440 10752 12492 10804
rect 4436 10684 4488 10736
rect 3608 10616 3660 10668
rect 7104 10616 7156 10668
rect 7564 10616 7616 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 6276 10548 6328 10600
rect 7932 10548 7984 10600
rect 3792 10480 3844 10532
rect 4436 10523 4488 10532
rect 4436 10489 4445 10523
rect 4445 10489 4479 10523
rect 4479 10489 4488 10523
rect 4436 10480 4488 10489
rect 6920 10480 6972 10532
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 12440 10480 12492 10532
rect 4988 10412 5040 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 8208 10412 8260 10464
rect 8852 10412 8904 10464
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 8315 10310 8367 10362
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 15648 10310 15700 10362
rect 15712 10310 15764 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 6920 10208 6972 10260
rect 10324 10208 10376 10260
rect 10876 10208 10928 10260
rect 15200 10208 15252 10260
rect 4252 10183 4304 10192
rect 4252 10149 4261 10183
rect 4261 10149 4295 10183
rect 4295 10149 4304 10183
rect 4252 10140 4304 10149
rect 4436 10140 4488 10192
rect 4988 10140 5040 10192
rect 6000 10183 6052 10192
rect 6000 10149 6009 10183
rect 6009 10149 6043 10183
rect 6043 10149 6052 10183
rect 6000 10140 6052 10149
rect 6276 10140 6328 10192
rect 7012 10183 7064 10192
rect 7012 10149 7021 10183
rect 7021 10149 7055 10183
rect 7055 10149 7064 10183
rect 7012 10140 7064 10149
rect 7564 10183 7616 10192
rect 7564 10149 7573 10183
rect 7573 10149 7607 10183
rect 7607 10149 7616 10183
rect 7564 10140 7616 10149
rect 7748 10140 7800 10192
rect 17224 10140 17276 10192
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3884 10004 3936 10056
rect 10232 10115 10284 10124
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 11520 10072 11572 10124
rect 12164 10072 12216 10124
rect 12532 10072 12584 10124
rect 15384 10072 15436 10124
rect 7196 10004 7248 10056
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 2964 9868 3016 9920
rect 11244 9868 11296 9920
rect 4648 9766 4700 9818
rect 4712 9766 4764 9818
rect 4776 9766 4828 9818
rect 4840 9766 4892 9818
rect 11982 9766 12034 9818
rect 12046 9766 12098 9818
rect 12110 9766 12162 9818
rect 12174 9766 12226 9818
rect 19315 9766 19367 9818
rect 19379 9766 19431 9818
rect 19443 9766 19495 9818
rect 19507 9766 19559 9818
rect 2504 9664 2556 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 7564 9664 7616 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 3792 9596 3844 9648
rect 6736 9596 6788 9648
rect 8024 9596 8076 9648
rect 12440 9596 12492 9648
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 12532 9528 12584 9580
rect 1676 9460 1728 9512
rect 2964 9460 3016 9512
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4528 9460 4580 9469
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 2688 9324 2740 9376
rect 5540 9392 5592 9444
rect 7748 9324 7800 9376
rect 9680 9392 9732 9444
rect 9956 9435 10008 9444
rect 9956 9401 9965 9435
rect 9965 9401 9999 9435
rect 9999 9401 10008 9435
rect 9956 9392 10008 9401
rect 10968 9435 11020 9444
rect 10968 9401 10977 9435
rect 10977 9401 11011 9435
rect 11011 9401 11020 9435
rect 10968 9392 11020 9401
rect 11520 9324 11572 9376
rect 15384 9367 15436 9376
rect 15384 9333 15393 9367
rect 15393 9333 15427 9367
rect 15427 9333 15436 9367
rect 15384 9324 15436 9333
rect 8315 9222 8367 9274
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 15648 9222 15700 9274
rect 15712 9222 15764 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 2688 9052 2740 9104
rect 4252 9120 4304 9172
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 6552 9120 6604 9172
rect 9312 9163 9364 9172
rect 5540 9052 5592 9104
rect 9312 9129 9321 9163
rect 9321 9129 9355 9163
rect 9355 9129 9364 9163
rect 9312 9120 9364 9129
rect 6736 9095 6788 9104
rect 6736 9061 6745 9095
rect 6745 9061 6779 9095
rect 6779 9061 6788 9095
rect 6736 9052 6788 9061
rect 8024 9052 8076 9104
rect 9956 9052 10008 9104
rect 10508 9095 10560 9104
rect 10508 9061 10517 9095
rect 10517 9061 10551 9095
rect 10551 9061 10560 9095
rect 10508 9052 10560 9061
rect 10600 9095 10652 9104
rect 10600 9061 10609 9095
rect 10609 9061 10643 9095
rect 10643 9061 10652 9095
rect 10600 9052 10652 9061
rect 10968 9052 11020 9104
rect 1768 8916 1820 8968
rect 2872 8916 2924 8968
rect 3792 8848 3844 8900
rect 4620 8984 4672 9036
rect 4988 8984 5040 9036
rect 4528 8916 4580 8968
rect 9036 8984 9088 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 12348 9027 12400 9036
rect 11152 8984 11204 8993
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 5172 8848 5224 8900
rect 7196 8891 7248 8900
rect 7196 8857 7205 8891
rect 7205 8857 7239 8891
rect 7239 8857 7248 8891
rect 7196 8848 7248 8857
rect 9680 8848 9732 8900
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2136 8780 2188 8789
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 9312 8780 9364 8832
rect 4648 8678 4700 8730
rect 4712 8678 4764 8730
rect 4776 8678 4828 8730
rect 4840 8678 4892 8730
rect 11982 8678 12034 8730
rect 12046 8678 12098 8730
rect 12110 8678 12162 8730
rect 12174 8678 12226 8730
rect 19315 8678 19367 8730
rect 19379 8678 19431 8730
rect 19443 8678 19495 8730
rect 19507 8678 19559 8730
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 10600 8576 10652 8628
rect 11244 8576 11296 8628
rect 12348 8576 12400 8628
rect 10508 8508 10560 8560
rect 11152 8508 11204 8560
rect 2688 8440 2740 8492
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 8944 8440 8996 8492
rect 3792 8415 3844 8424
rect 3792 8381 3801 8415
rect 3801 8381 3835 8415
rect 3835 8381 3844 8415
rect 3792 8372 3844 8381
rect 3884 8372 3936 8424
rect 4528 8372 4580 8424
rect 5172 8372 5224 8424
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 6276 8372 6328 8424
rect 7564 8372 7616 8424
rect 11244 8372 11296 8424
rect 5080 8347 5132 8356
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 2688 8279 2740 8288
rect 2688 8245 2697 8279
rect 2697 8245 2731 8279
rect 2731 8245 2740 8279
rect 2688 8236 2740 8245
rect 2872 8279 2924 8288
rect 2872 8245 2881 8279
rect 2881 8245 2915 8279
rect 2915 8245 2924 8279
rect 2872 8236 2924 8245
rect 3608 8236 3660 8288
rect 4804 8236 4856 8288
rect 5080 8313 5089 8347
rect 5089 8313 5123 8347
rect 5123 8313 5132 8347
rect 5080 8304 5132 8313
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 8760 8304 8812 8356
rect 12716 8372 12768 8424
rect 6552 8236 6604 8245
rect 7288 8236 7340 8288
rect 9036 8236 9088 8288
rect 10232 8236 10284 8288
rect 8315 8134 8367 8186
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 15648 8134 15700 8186
rect 15712 8134 15764 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 3700 8032 3752 8084
rect 5080 8032 5132 8084
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 11152 8032 11204 8084
rect 2136 8007 2188 8016
rect 2136 7973 2145 8007
rect 2145 7973 2179 8007
rect 2179 7973 2188 8007
rect 2136 7964 2188 7973
rect 4252 7964 4304 8016
rect 4436 7964 4488 8016
rect 6276 8007 6328 8016
rect 1032 7896 1084 7948
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 6276 7973 6285 8007
rect 6285 7973 6319 8007
rect 6319 7973 6328 8007
rect 6276 7964 6328 7973
rect 7288 8007 7340 8016
rect 7288 7973 7297 8007
rect 7297 7973 7331 8007
rect 7331 7973 7340 8007
rect 7288 7964 7340 7973
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 2780 7828 2832 7880
rect 7840 7896 7892 7948
rect 8760 7896 8812 7948
rect 10876 7964 10928 8016
rect 10232 7896 10284 7948
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 3700 7692 3752 7744
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 4528 7692 4580 7744
rect 6460 7828 6512 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 9128 7828 9180 7880
rect 7932 7760 7984 7812
rect 6644 7692 6696 7744
rect 11888 7760 11940 7812
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9220 7692 9272 7744
rect 4648 7590 4700 7642
rect 4712 7590 4764 7642
rect 4776 7590 4828 7642
rect 4840 7590 4892 7642
rect 11982 7590 12034 7642
rect 12046 7590 12098 7642
rect 12110 7590 12162 7642
rect 12174 7590 12226 7642
rect 19315 7590 19367 7642
rect 19379 7590 19431 7642
rect 19443 7590 19495 7642
rect 19507 7590 19559 7642
rect 20 7488 72 7540
rect 3608 7488 3660 7540
rect 7748 7531 7800 7540
rect 2044 7420 2096 7472
rect 2228 7352 2280 7404
rect 2872 7352 2924 7404
rect 112 7284 164 7336
rect 1584 7284 1636 7336
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 4528 7420 4580 7472
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 10232 7531 10284 7540
rect 10232 7497 10241 7531
rect 10241 7497 10275 7531
rect 10275 7497 10284 7531
rect 10232 7488 10284 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 5816 7420 5868 7472
rect 6276 7463 6328 7472
rect 6276 7429 6285 7463
rect 6285 7429 6319 7463
rect 6319 7429 6328 7463
rect 6276 7420 6328 7429
rect 11704 7420 11756 7472
rect 11888 7420 11940 7472
rect 8944 7352 8996 7404
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 5264 7284 5316 7336
rect 2872 7216 2924 7268
rect 6644 7284 6696 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9312 7259 9364 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2228 7191 2280 7200
rect 2228 7157 2237 7191
rect 2237 7157 2271 7191
rect 2271 7157 2280 7191
rect 2228 7148 2280 7157
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3332 7148 3384 7200
rect 4252 7148 4304 7200
rect 6552 7148 6604 7200
rect 9312 7225 9321 7259
rect 9321 7225 9355 7259
rect 9355 7225 9364 7259
rect 9312 7216 9364 7225
rect 9404 7259 9456 7268
rect 9404 7225 9413 7259
rect 9413 7225 9447 7259
rect 9447 7225 9456 7259
rect 9404 7216 9456 7225
rect 10600 7216 10652 7268
rect 10968 7259 11020 7268
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 7840 7148 7892 7200
rect 11704 7148 11756 7200
rect 12624 7148 12676 7200
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 8315 7046 8367 7098
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 15648 7046 15700 7098
rect 15712 7046 15764 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2504 6944 2556 6996
rect 1768 6876 1820 6928
rect 5724 6944 5776 6996
rect 7288 6944 7340 6996
rect 7840 6944 7892 6996
rect 9312 6944 9364 6996
rect 5356 6876 5408 6928
rect 2688 6808 2740 6860
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 5172 6808 5224 6860
rect 6828 6876 6880 6928
rect 10692 6919 10744 6928
rect 10692 6885 10701 6919
rect 10701 6885 10735 6919
rect 10735 6885 10744 6919
rect 10692 6876 10744 6885
rect 11244 6919 11296 6928
rect 11244 6885 11253 6919
rect 11253 6885 11287 6919
rect 11287 6885 11296 6919
rect 11244 6876 11296 6885
rect 6460 6851 6512 6860
rect 2780 6740 2832 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 11336 6808 11388 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 13728 6808 13780 6860
rect 6184 6740 6236 6792
rect 6736 6740 6788 6792
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 3700 6647 3752 6656
rect 3700 6613 3709 6647
rect 3709 6613 3743 6647
rect 3743 6613 3752 6647
rect 3700 6604 3752 6613
rect 8116 6672 8168 6724
rect 4988 6604 5040 6656
rect 8668 6604 8720 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 10048 6604 10100 6656
rect 11704 6604 11756 6656
rect 4648 6502 4700 6554
rect 4712 6502 4764 6554
rect 4776 6502 4828 6554
rect 4840 6502 4892 6554
rect 11982 6502 12034 6554
rect 12046 6502 12098 6554
rect 12110 6502 12162 6554
rect 12174 6502 12226 6554
rect 19315 6502 19367 6554
rect 19379 6502 19431 6554
rect 19443 6502 19495 6554
rect 19507 6502 19559 6554
rect 1768 6400 1820 6452
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2504 6400 2556 6452
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 2320 6264 2372 6316
rect 1676 6196 1728 6248
rect 3700 6264 3752 6316
rect 8024 6332 8076 6384
rect 9404 6400 9456 6452
rect 12348 6400 12400 6452
rect 9220 6332 9272 6384
rect 9772 6264 9824 6316
rect 10968 6264 11020 6316
rect 1400 6171 1452 6180
rect 1400 6137 1409 6171
rect 1409 6137 1443 6171
rect 1443 6137 1452 6171
rect 1400 6128 1452 6137
rect 2136 6128 2188 6180
rect 2504 6128 2556 6180
rect 4804 6196 4856 6248
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 10048 6196 10100 6248
rect 10692 6196 10744 6248
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 8760 6128 8812 6180
rect 2964 6060 3016 6112
rect 5172 6060 5224 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 7840 6060 7892 6112
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 8315 5958 8367 6010
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 15648 5958 15700 6010
rect 15712 5958 15764 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 2596 5856 2648 5908
rect 4252 5856 4304 5908
rect 4804 5831 4856 5840
rect 4804 5797 4813 5831
rect 4813 5797 4847 5831
rect 4847 5797 4856 5831
rect 4804 5788 4856 5797
rect 5080 5788 5132 5840
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 2596 5720 2648 5772
rect 3608 5720 3660 5772
rect 3792 5720 3844 5772
rect 5172 5720 5224 5772
rect 6184 5788 6236 5840
rect 6736 5831 6788 5840
rect 6736 5797 6745 5831
rect 6745 5797 6779 5831
rect 6779 5797 6788 5831
rect 6736 5788 6788 5797
rect 8668 5788 8720 5840
rect 9680 5788 9732 5840
rect 10232 5856 10284 5908
rect 11336 5856 11388 5908
rect 12532 5899 12584 5908
rect 12532 5865 12541 5899
rect 12541 5865 12575 5899
rect 12575 5865 12584 5899
rect 12532 5856 12584 5865
rect 12900 5856 12952 5908
rect 10600 5788 10652 5840
rect 11612 5788 11664 5840
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 12440 5720 12492 5772
rect 12900 5763 12952 5772
rect 12900 5729 12944 5763
rect 12944 5729 12952 5763
rect 12900 5720 12952 5729
rect 7196 5652 7248 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 10968 5652 11020 5704
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 8116 5584 8168 5636
rect 5080 5559 5132 5568
rect 5080 5525 5089 5559
rect 5089 5525 5123 5559
rect 5123 5525 5132 5559
rect 5080 5516 5132 5525
rect 7104 5559 7156 5568
rect 7104 5525 7113 5559
rect 7113 5525 7147 5559
rect 7147 5525 7156 5559
rect 7104 5516 7156 5525
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 10324 5516 10376 5568
rect 11796 5516 11848 5568
rect 4648 5414 4700 5466
rect 4712 5414 4764 5466
rect 4776 5414 4828 5466
rect 4840 5414 4892 5466
rect 11982 5414 12034 5466
rect 12046 5414 12098 5466
rect 12110 5414 12162 5466
rect 12174 5414 12226 5466
rect 19315 5414 19367 5466
rect 19379 5414 19431 5466
rect 19443 5414 19495 5466
rect 19507 5414 19559 5466
rect 2596 5312 2648 5364
rect 3608 5312 3660 5364
rect 8024 5355 8076 5364
rect 2504 5176 2556 5228
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 11428 5312 11480 5364
rect 6736 5244 6788 5296
rect 9312 5244 9364 5296
rect 9680 5244 9732 5296
rect 4344 5176 4396 5228
rect 1400 5108 1452 5160
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 2136 4972 2188 5024
rect 4896 5151 4948 5160
rect 4252 5040 4304 5092
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 5080 5108 5132 5160
rect 6644 5176 6696 5228
rect 11152 5176 11204 5228
rect 11704 5176 11756 5228
rect 12900 5176 12952 5228
rect 13360 5176 13412 5228
rect 13544 5176 13596 5228
rect 5448 5108 5500 5160
rect 6368 5108 6420 5160
rect 8208 5108 8260 5160
rect 9128 5108 9180 5160
rect 5172 4972 5224 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 7840 5040 7892 5092
rect 8760 5040 8812 5092
rect 9680 5040 9732 5092
rect 10968 5083 11020 5092
rect 7748 5015 7800 5024
rect 6552 4972 6604 4981
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8116 4972 8168 5024
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 11980 5040 12032 5092
rect 12440 5083 12492 5092
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 10600 4972 10652 5024
rect 11612 4972 11664 5024
rect 8315 4870 8367 4922
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 15648 4870 15700 4922
rect 15712 4870 15764 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 1768 4768 1820 4820
rect 3792 4768 3844 4820
rect 4252 4768 4304 4820
rect 4896 4768 4948 4820
rect 7104 4768 7156 4820
rect 7840 4768 7892 4820
rect 1400 4700 1452 4752
rect 2412 4700 2464 4752
rect 6644 4743 6696 4752
rect 4068 4675 4120 4684
rect 1952 4564 2004 4616
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 6644 4709 6653 4743
rect 6653 4709 6687 4743
rect 6687 4709 6696 4743
rect 6644 4700 6696 4709
rect 7196 4700 7248 4752
rect 7564 4743 7616 4752
rect 7564 4709 7573 4743
rect 7573 4709 7607 4743
rect 7607 4709 7616 4743
rect 7564 4700 7616 4709
rect 7748 4700 7800 4752
rect 11336 4768 11388 4820
rect 9220 4700 9272 4752
rect 9680 4700 9732 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 5908 4632 5960 4684
rect 6368 4675 6420 4684
rect 5724 4564 5776 4616
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 7564 4564 7616 4616
rect 11336 4564 11388 4616
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 1860 4496 1912 4548
rect 2320 4496 2372 4548
rect 4436 4496 4488 4548
rect 4528 4428 4580 4480
rect 6828 4428 6880 4480
rect 8024 4496 8076 4548
rect 8760 4496 8812 4548
rect 13820 4496 13872 4548
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 11428 4428 11480 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 4648 4326 4700 4378
rect 4712 4326 4764 4378
rect 4776 4326 4828 4378
rect 4840 4326 4892 4378
rect 11982 4326 12034 4378
rect 12046 4326 12098 4378
rect 12110 4326 12162 4378
rect 12174 4326 12226 4378
rect 19315 4326 19367 4378
rect 19379 4326 19431 4378
rect 19443 4326 19495 4378
rect 19507 4326 19559 4378
rect 1952 4224 2004 4276
rect 2320 4267 2372 4276
rect 2320 4233 2329 4267
rect 2329 4233 2363 4267
rect 2363 4233 2372 4267
rect 2320 4224 2372 4233
rect 5908 4224 5960 4276
rect 10968 4224 11020 4276
rect 12532 4224 12584 4276
rect 13176 4224 13228 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 13636 4224 13688 4276
rect 8208 4156 8260 4208
rect 11152 4199 11204 4208
rect 11152 4165 11161 4199
rect 11161 4165 11195 4199
rect 11195 4165 11204 4199
rect 11152 4156 11204 4165
rect 1860 4088 1912 4140
rect 2872 4088 2924 4140
rect 2964 4088 3016 4140
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 4436 4020 4488 4072
rect 6736 4088 6788 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8944 4131 8996 4140
rect 8668 4088 8720 4097
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 12992 4156 13044 4208
rect 11888 4088 11940 4140
rect 12532 4063 12584 4072
rect 2412 3952 2464 4004
rect 4712 3995 4764 4004
rect 4712 3961 4721 3995
rect 4721 3961 4755 3995
rect 4755 3961 4764 3995
rect 4712 3952 4764 3961
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5908 3995 5960 4004
rect 5356 3952 5408 3961
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 1952 3884 2004 3936
rect 3976 3884 4028 3936
rect 4068 3884 4120 3936
rect 4528 3884 4580 3936
rect 5172 3884 5224 3936
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 7840 3884 7892 3936
rect 8116 3884 8168 3936
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 13820 4020 13872 4072
rect 8760 3995 8812 4004
rect 8760 3961 8769 3995
rect 8769 3961 8803 3995
rect 8803 3961 8812 3995
rect 8760 3952 8812 3961
rect 10324 3952 10376 4004
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 11796 3952 11848 4004
rect 12348 3884 12400 3936
rect 20996 3884 21048 3936
rect 8315 3782 8367 3834
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 15648 3782 15700 3834
rect 15712 3782 15764 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 2964 3680 3016 3732
rect 3148 3680 3200 3732
rect 3792 3680 3844 3732
rect 3976 3680 4028 3732
rect 4160 3680 4212 3732
rect 5540 3680 5592 3732
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 2320 3612 2372 3664
rect 2780 3612 2832 3664
rect 7748 3680 7800 3732
rect 10968 3680 11020 3732
rect 11336 3723 11388 3732
rect 11336 3689 11345 3723
rect 11345 3689 11379 3723
rect 11379 3689 11388 3723
rect 11336 3680 11388 3689
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 12716 3680 12768 3732
rect 8760 3612 8812 3664
rect 10048 3655 10100 3664
rect 10048 3621 10057 3655
rect 10057 3621 10091 3655
rect 10091 3621 10100 3655
rect 10048 3612 10100 3621
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 12624 3612 12676 3664
rect 1952 3544 2004 3596
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 5724 3587 5776 3596
rect 1676 3476 1728 3528
rect 3884 3408 3936 3460
rect 5080 3408 5132 3460
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 5816 3544 5868 3596
rect 6368 3544 6420 3596
rect 8208 3544 8260 3596
rect 13176 3544 13228 3596
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 15200 3587 15252 3596
rect 15200 3553 15209 3587
rect 15209 3553 15243 3587
rect 15243 3553 15252 3587
rect 15200 3544 15252 3553
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 7656 3519 7708 3528
rect 5908 3408 5960 3460
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8024 3476 8076 3528
rect 8208 3408 8260 3460
rect 10508 3451 10560 3460
rect 10508 3417 10517 3451
rect 10517 3417 10551 3451
rect 10551 3417 10560 3451
rect 10508 3408 10560 3417
rect 11244 3408 11296 3460
rect 2136 3383 2188 3392
rect 2136 3349 2145 3383
rect 2145 3349 2179 3383
rect 2179 3349 2188 3383
rect 2136 3340 2188 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 3332 3340 3384 3392
rect 4160 3340 4212 3392
rect 5356 3340 5408 3392
rect 10784 3340 10836 3392
rect 14004 3476 14056 3528
rect 11796 3408 11848 3460
rect 12624 3408 12676 3460
rect 13636 3408 13688 3460
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 13360 3340 13412 3392
rect 4648 3238 4700 3290
rect 4712 3238 4764 3290
rect 4776 3238 4828 3290
rect 4840 3238 4892 3290
rect 11982 3238 12034 3290
rect 12046 3238 12098 3290
rect 12110 3238 12162 3290
rect 12174 3238 12226 3290
rect 19315 3238 19367 3290
rect 19379 3238 19431 3290
rect 19443 3238 19495 3290
rect 19507 3238 19559 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 4344 3179 4396 3188
rect 4344 3145 4353 3179
rect 4353 3145 4387 3179
rect 4387 3145 4396 3179
rect 4344 3136 4396 3145
rect 5724 3136 5776 3188
rect 6920 3136 6972 3188
rect 8944 3136 8996 3188
rect 9128 3136 9180 3188
rect 10692 3136 10744 3188
rect 10876 3136 10928 3188
rect 11612 3136 11664 3188
rect 13544 3179 13596 3188
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 13636 3136 13688 3188
rect 2136 3068 2188 3120
rect 3884 3111 3936 3120
rect 3884 3077 3893 3111
rect 3893 3077 3927 3111
rect 3927 3077 3936 3111
rect 3884 3068 3936 3077
rect 9956 3068 10008 3120
rect 6920 3043 6972 3052
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 3608 2907 3660 2916
rect 3608 2873 3617 2907
rect 3617 2873 3651 2907
rect 3651 2873 3660 2907
rect 3608 2864 3660 2873
rect 3516 2796 3568 2848
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7656 3000 7708 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 5356 2932 5408 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 8208 2932 8260 2984
rect 10048 3000 10100 3052
rect 12808 3068 12860 3120
rect 15936 3068 15988 3120
rect 10784 2932 10836 2984
rect 10968 2932 11020 2984
rect 4988 2864 5040 2916
rect 7104 2864 7156 2916
rect 7932 2864 7984 2916
rect 9680 2864 9732 2916
rect 5632 2796 5684 2848
rect 8116 2796 8168 2848
rect 8852 2796 8904 2848
rect 11244 2796 11296 2848
rect 12624 3000 12676 3052
rect 12992 3000 13044 3052
rect 15476 2932 15528 2984
rect 14004 2796 14056 2848
rect 14556 2796 14608 2848
rect 15200 2796 15252 2848
rect 8315 2694 8367 2746
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 15648 2694 15700 2746
rect 15712 2694 15764 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 1952 2592 2004 2644
rect 2320 2592 2372 2644
rect 2228 2524 2280 2576
rect 4160 2592 4212 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4252 2524 4304 2576
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 4528 2456 4580 2465
rect 5080 2524 5132 2576
rect 8208 2592 8260 2644
rect 9864 2592 9916 2644
rect 10876 2635 10928 2644
rect 6552 2567 6604 2576
rect 6552 2533 6561 2567
rect 6561 2533 6595 2567
rect 6595 2533 6604 2567
rect 6552 2524 6604 2533
rect 7932 2524 7984 2576
rect 8116 2567 8168 2576
rect 8116 2533 8125 2567
rect 8125 2533 8159 2567
rect 8159 2533 8168 2567
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 11336 2592 11388 2644
rect 14004 2592 14056 2644
rect 17132 2635 17184 2644
rect 17132 2601 17141 2635
rect 17141 2601 17175 2635
rect 17175 2601 17184 2635
rect 17132 2592 17184 2601
rect 8116 2524 8168 2533
rect 10048 2524 10100 2576
rect 13360 2524 13412 2576
rect 5356 2499 5408 2508
rect 5356 2465 5365 2499
rect 5365 2465 5399 2499
rect 5399 2465 5408 2499
rect 5356 2456 5408 2465
rect 5632 2456 5684 2508
rect 6184 2456 6236 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7104 2456 7156 2508
rect 5448 2388 5500 2440
rect 9220 2456 9272 2508
rect 10508 2499 10560 2508
rect 10508 2465 10517 2499
rect 10517 2465 10551 2499
rect 10551 2465 10560 2499
rect 10508 2456 10560 2465
rect 10692 2456 10744 2508
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 3608 2320 3660 2372
rect 10048 2388 10100 2440
rect 11244 2388 11296 2440
rect 3516 2252 3568 2304
rect 5448 2252 5500 2304
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 9588 2252 9640 2304
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 17132 2320 17184 2372
rect 14556 2252 14608 2304
rect 4648 2150 4700 2202
rect 4712 2150 4764 2202
rect 4776 2150 4828 2202
rect 4840 2150 4892 2202
rect 11982 2150 12034 2202
rect 12046 2150 12098 2202
rect 12110 2150 12162 2202
rect 12174 2150 12226 2202
rect 19315 2150 19367 2202
rect 19379 2150 19431 2202
rect 19443 2150 19495 2202
rect 19507 2150 19559 2202
rect 9220 2048 9272 2100
rect 11520 2048 11572 2100
rect 12624 2048 12676 2100
rect 13084 2048 13136 2100
rect 15476 2048 15528 2100
rect 8392 76 8444 128
rect 12808 76 12860 128
<< metal2 >>
rect 20 21548 72 21554
rect 846 21548 902 22000
rect 846 21520 848 21548
rect 20 21490 72 21496
rect 900 21520 902 21548
rect 1676 21548 1728 21554
rect 848 21490 900 21496
rect 2502 21548 2558 22000
rect 4158 21570 4214 22000
rect 2502 21520 2504 21548
rect 1676 21490 1728 21496
rect 2556 21520 2558 21548
rect 4080 21542 4214 21570
rect 2504 21490 2556 21496
rect 32 7546 60 21490
rect 860 21459 888 21490
rect 1398 20360 1454 20369
rect 1398 20295 1454 20304
rect 1306 16008 1362 16017
rect 1306 15943 1362 15952
rect 1320 11694 1348 15943
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1412 10810 1440 20295
rect 1582 11928 1638 11937
rect 1582 11863 1638 11872
rect 1596 11830 1624 11863
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 10441 1440 10542
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1688 9518 1716 21490
rect 2516 21459 2544 21490
rect 4080 19334 4108 21542
rect 4158 21520 4214 21542
rect 5906 21570 5962 22000
rect 7562 21570 7618 22000
rect 5906 21542 6224 21570
rect 5906 21520 5962 21542
rect 4622 19612 4918 19632
rect 4678 19610 4702 19612
rect 4758 19610 4782 19612
rect 4838 19610 4862 19612
rect 4700 19558 4702 19610
rect 4764 19558 4776 19610
rect 4838 19558 4840 19610
rect 4678 19556 4702 19558
rect 4758 19556 4782 19558
rect 4838 19556 4862 19558
rect 4622 19536 4918 19556
rect 4080 19306 4292 19334
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4172 16998 4200 17682
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 11218 2636 11630
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10810 2636 11154
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 3620 10674 3648 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3804 10538 3832 10950
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1032 7948 1084 7954
rect 1032 7890 1084 7896
rect 110 7712 166 7721
rect 110 7647 166 7656
rect 20 7540 72 7546
rect 20 7482 72 7488
rect 124 7342 152 7647
rect 112 7336 164 7342
rect 112 7278 164 7284
rect 110 5536 166 5545
rect 110 5471 166 5480
rect 124 4593 152 5471
rect 110 4584 166 4593
rect 110 4519 166 4528
rect 662 82 718 480
rect 1044 82 1072 7890
rect 1596 7342 1624 8230
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1412 5166 1440 6122
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4758 1440 5102
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 1596 3777 1624 7142
rect 1688 7002 1716 9114
rect 1780 8974 1808 9862
rect 2516 9722 2544 10066
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1688 6254 1716 6938
rect 1768 6928 1820 6934
rect 1768 6870 1820 6876
rect 1780 6458 1808 6870
rect 1768 6452 1820 6458
rect 1820 6412 1900 6440
rect 1768 6394 1820 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5166 1716 6190
rect 1780 5778 1808 6258
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1688 4826 1716 5102
rect 1780 4826 1808 5714
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1582 3768 1638 3777
rect 1582 3703 1638 3712
rect 1688 3534 1716 4762
rect 1780 4154 1808 4762
rect 1872 4554 1900 6412
rect 1964 4622 1992 9318
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8022 2176 8774
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 2056 6458 2084 7414
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2148 6186 2176 7958
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7206 2268 7346
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2136 5024 2188 5030
rect 2240 5012 2268 7142
rect 2516 7002 2544 9658
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2516 6458 2544 6938
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5778 2360 6258
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2516 5778 2544 6122
rect 2608 5914 2636 9998
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9518 3004 9862
rect 3804 9654 3832 10474
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 9110 2728 9318
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2700 8498 2728 9046
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2884 8294 2912 8910
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2700 6866 2728 8230
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7342 2820 7822
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7410 2912 7686
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2792 6798 2820 7278
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2596 5908 2648 5914
rect 2648 5868 2728 5896
rect 2596 5850 2648 5856
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2516 5234 2544 5714
rect 2608 5370 2636 5714
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2188 4984 2268 5012
rect 2136 4966 2188 4972
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1964 4282 1992 4558
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1780 4146 1900 4154
rect 1780 4140 1912 4146
rect 1780 4126 1860 4140
rect 1860 4082 1912 4088
rect 1872 3942 1900 4082
rect 1860 3936 1912 3942
rect 1858 3904 1860 3913
rect 1952 3936 2004 3942
rect 1912 3904 1914 3913
rect 1952 3878 2004 3884
rect 1858 3839 1914 3848
rect 1872 3813 1900 3839
rect 1964 3602 1992 3878
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 3194 1716 3470
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1964 2650 1992 3538
rect 2148 3398 2176 4966
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2332 4282 2360 4490
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2332 3670 2360 4218
rect 2424 4010 2452 4694
rect 2700 4622 2728 5868
rect 2688 4616 2740 4622
rect 2740 4576 2820 4604
rect 2688 4558 2740 4564
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2320 3664 2372 3670
rect 2424 3641 2452 3946
rect 2792 3670 2820 4576
rect 2884 4146 2912 7210
rect 2976 7206 3004 9454
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8430 3832 8842
rect 3896 8838 3924 9998
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8430 3924 8774
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3344 7342 3372 8366
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 7546 3648 8230
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3712 7750 3740 8026
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3620 7342 3648 7482
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3344 7206 3372 7278
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6118 3004 6802
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 3620 5778 3648 7278
rect 3712 6662 3740 7686
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6322 3740 6598
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3804 5778 3832 8366
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3620 5370 3648 5714
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3804 4826 3832 5714
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2976 3738 3004 4082
rect 3804 4078 3832 4762
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3804 3738 3832 4014
rect 4080 3942 4108 4626
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3988 3738 4016 3878
rect 4172 3738 4200 16934
rect 4264 11218 4292 19306
rect 4622 18524 4918 18544
rect 4678 18522 4702 18524
rect 4758 18522 4782 18524
rect 4838 18522 4862 18524
rect 4700 18470 4702 18522
rect 4764 18470 4776 18522
rect 4838 18470 4840 18522
rect 4678 18468 4702 18470
rect 4758 18468 4782 18470
rect 4838 18468 4862 18470
rect 4622 18448 4918 18468
rect 6196 18426 6224 21542
rect 7392 21542 7618 21570
rect 7392 18426 7420 21542
rect 7562 21520 7618 21542
rect 8668 21548 8720 21554
rect 9218 21548 9274 22000
rect 9218 21520 9220 21548
rect 8668 21490 8720 21496
rect 9272 21520 9274 21548
rect 9680 21548 9732 21554
rect 9220 21490 9272 21496
rect 10966 21548 11022 22000
rect 12622 21570 12678 22000
rect 10966 21520 10968 21548
rect 9680 21490 9732 21496
rect 11020 21520 11022 21548
rect 12452 21542 12678 21570
rect 10968 21490 11020 21496
rect 8289 19068 8585 19088
rect 8345 19066 8369 19068
rect 8425 19066 8449 19068
rect 8505 19066 8529 19068
rect 8367 19014 8369 19066
rect 8431 19014 8443 19066
rect 8505 19014 8507 19066
rect 8345 19012 8369 19014
rect 8425 19012 8449 19014
rect 8505 19012 8529 19014
rect 8289 18992 8585 19012
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 6196 18222 6224 18362
rect 6184 18216 6236 18222
rect 4802 18184 4858 18193
rect 6184 18158 6236 18164
rect 4802 18119 4858 18128
rect 4816 17882 4844 18119
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4622 17436 4918 17456
rect 4678 17434 4702 17436
rect 4758 17434 4782 17436
rect 4838 17434 4862 17436
rect 4700 17382 4702 17434
rect 4764 17382 4776 17434
rect 4838 17382 4840 17434
rect 4678 17380 4702 17382
rect 4758 17380 4782 17382
rect 4838 17380 4862 17382
rect 4622 17360 4918 17380
rect 4622 16348 4918 16368
rect 4678 16346 4702 16348
rect 4758 16346 4782 16348
rect 4838 16346 4862 16348
rect 4700 16294 4702 16346
rect 4764 16294 4776 16346
rect 4838 16294 4840 16346
rect 4678 16292 4702 16294
rect 4758 16292 4782 16294
rect 4838 16292 4862 16294
rect 4622 16272 4918 16292
rect 4622 15260 4918 15280
rect 4678 15258 4702 15260
rect 4758 15258 4782 15260
rect 4838 15258 4862 15260
rect 4700 15206 4702 15258
rect 4764 15206 4776 15258
rect 4838 15206 4840 15258
rect 4678 15204 4702 15206
rect 4758 15204 4782 15206
rect 4838 15204 4862 15206
rect 4622 15184 4918 15204
rect 4622 14172 4918 14192
rect 4678 14170 4702 14172
rect 4758 14170 4782 14172
rect 4838 14170 4862 14172
rect 4700 14118 4702 14170
rect 4764 14118 4776 14170
rect 4838 14118 4840 14170
rect 4678 14116 4702 14118
rect 4758 14116 4782 14118
rect 4838 14116 4862 14118
rect 4622 14096 4918 14116
rect 4622 13084 4918 13104
rect 4678 13082 4702 13084
rect 4758 13082 4782 13084
rect 4838 13082 4862 13084
rect 4700 13030 4702 13082
rect 4764 13030 4776 13082
rect 4838 13030 4840 13082
rect 4678 13028 4702 13030
rect 4758 13028 4782 13030
rect 4838 13028 4862 13030
rect 4622 13008 4918 13028
rect 4622 11996 4918 12016
rect 4678 11994 4702 11996
rect 4758 11994 4782 11996
rect 4838 11994 4862 11996
rect 4700 11942 4702 11994
rect 4764 11942 4776 11994
rect 4838 11942 4840 11994
rect 4678 11940 4702 11942
rect 4758 11940 4782 11942
rect 4838 11940 4862 11942
rect 4622 11920 4918 11940
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4622 10908 4918 10928
rect 4678 10906 4702 10908
rect 4758 10906 4782 10908
rect 4838 10906 4862 10908
rect 4700 10854 4702 10906
rect 4764 10854 4776 10906
rect 4838 10854 4840 10906
rect 4678 10852 4702 10854
rect 4758 10852 4782 10854
rect 4838 10852 4862 10854
rect 4622 10832 4918 10852
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4448 10538 4476 10678
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4448 10198 4476 10474
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10198 5028 10406
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4264 9178 4292 10134
rect 4622 9820 4918 9840
rect 4678 9818 4702 9820
rect 4758 9818 4782 9820
rect 4838 9818 4862 9820
rect 4700 9766 4702 9818
rect 4764 9766 4776 9818
rect 4838 9766 4840 9818
rect 4678 9764 4702 9766
rect 4758 9764 4782 9766
rect 4838 9764 4862 9766
rect 4622 9744 4918 9764
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 9178 4568 9454
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4448 9042 4660 9058
rect 4448 9036 4672 9042
rect 4448 9030 4620 9036
rect 4448 8022 4476 9030
rect 4620 8978 4672 8984
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8430 4568 8910
rect 4622 8732 4918 8752
rect 4678 8730 4702 8732
rect 4758 8730 4782 8732
rect 4838 8730 4862 8732
rect 4700 8678 4702 8730
rect 4764 8678 4776 8730
rect 4838 8678 4840 8730
rect 4678 8676 4702 8678
rect 4758 8676 4782 8678
rect 4838 8676 4862 8678
rect 4622 8656 4918 8676
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4264 7750 4292 7958
rect 4540 7750 4568 8366
rect 4804 8288 4856 8294
rect 5000 8276 5028 8978
rect 5092 8945 5120 18022
rect 7562 13832 7618 13841
rect 7562 13767 7618 13776
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11354 7144 11494
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 5644 10470 5672 11154
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 9110 5580 9386
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 8430 5212 8842
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4856 8248 5028 8276
rect 4804 8230 4856 8236
rect 5092 8090 5120 8298
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4264 7206 4292 7686
rect 4540 7478 4568 7686
rect 4622 7644 4918 7664
rect 4678 7642 4702 7644
rect 4758 7642 4782 7644
rect 4838 7642 4862 7644
rect 4700 7590 4702 7642
rect 4764 7590 4776 7642
rect 4838 7590 4840 7642
rect 4678 7588 4702 7590
rect 4758 7588 4782 7590
rect 4838 7588 4862 7590
rect 4622 7568 4918 7588
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4264 5914 4292 6734
rect 5000 6662 5028 7890
rect 5184 6866 5212 8366
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5276 6916 5304 7278
rect 5356 6928 5408 6934
rect 5276 6888 5356 6916
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4622 6556 4918 6576
rect 4678 6554 4702 6556
rect 4758 6554 4782 6556
rect 4838 6554 4862 6556
rect 4700 6502 4702 6554
rect 4764 6502 4776 6554
rect 4838 6502 4840 6554
rect 4678 6500 4702 6502
rect 4758 6500 4782 6502
rect 4838 6500 4862 6502
rect 4622 6480 4918 6500
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5953 4844 6190
rect 4802 5944 4858 5953
rect 4252 5908 4304 5914
rect 4802 5879 4858 5888
rect 4252 5850 4304 5856
rect 4816 5846 4844 5879
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4622 5468 4918 5488
rect 4678 5466 4702 5468
rect 4758 5466 4782 5468
rect 4838 5466 4862 5468
rect 4700 5414 4702 5466
rect 4764 5414 4776 5466
rect 4838 5414 4840 5466
rect 4678 5412 4702 5414
rect 4758 5412 4782 5414
rect 4838 5412 4862 5414
rect 4622 5392 4918 5412
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4264 4826 4292 5034
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 2780 3664 2832 3670
rect 2320 3606 2372 3612
rect 2410 3632 2466 3641
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 3126 2176 3334
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2148 1737 2176 3062
rect 2332 2650 2360 3606
rect 2410 3567 2466 3576
rect 2686 3632 2742 3641
rect 2780 3606 2832 3612
rect 2686 3567 2742 3576
rect 2700 3398 2728 3567
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 3160 2990 3188 3674
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 2990 3372 3334
rect 3896 3126 3924 3402
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 2134 1728 2190 1737
rect 2134 1663 2190 1672
rect 662 54 1072 82
rect 1950 82 2006 480
rect 2240 82 2268 2518
rect 3528 2310 3556 2790
rect 3620 2378 3648 2858
rect 4172 2650 4200 3334
rect 4356 3194 4384 5170
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 4826 4936 5102
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4078 4476 4490
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 4072 4488 4078
rect 4540 4049 4568 4422
rect 4622 4380 4918 4400
rect 4678 4378 4702 4380
rect 4758 4378 4782 4380
rect 4838 4378 4862 4380
rect 4700 4326 4702 4378
rect 4764 4326 4776 4378
rect 4838 4326 4840 4378
rect 4678 4324 4702 4326
rect 4758 4324 4782 4326
rect 4838 4324 4862 4326
rect 4622 4304 4918 4324
rect 4436 4014 4488 4020
rect 4526 4040 4582 4049
rect 4526 3975 4582 3984
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4528 3936 4580 3942
rect 4724 3913 4752 3946
rect 4528 3878 4580 3884
rect 4710 3904 4766 3913
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4356 2650 4384 3130
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 1950 54 2268 82
rect 3238 82 3294 480
rect 3528 82 3556 2246
rect 3238 54 3556 82
rect 4264 82 4292 2518
rect 4540 2514 4568 3878
rect 4710 3839 4766 3848
rect 5000 3602 5028 6598
rect 5184 6118 5212 6802
rect 5276 6458 5304 6888
rect 5356 6870 5408 6876
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5092 5574 5120 5782
rect 5184 5778 5212 6054
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5092 5166 5120 5510
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 5184 5030 5212 5714
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4690 5212 4966
rect 5460 4729 5488 5102
rect 5446 4720 5502 4729
rect 5172 4684 5224 4690
rect 5446 4655 5502 4664
rect 5172 4626 5224 4632
rect 5184 3942 5212 4626
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4622 3292 4918 3312
rect 4678 3290 4702 3292
rect 4758 3290 4782 3292
rect 4838 3290 4862 3292
rect 4700 3238 4702 3290
rect 4764 3238 4776 3290
rect 4838 3238 4840 3290
rect 4678 3236 4702 3238
rect 4758 3236 4782 3238
rect 4838 3236 4862 3238
rect 4622 3216 4918 3236
rect 5000 2922 5028 3538
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 5092 2990 5120 3402
rect 5368 3398 5396 3946
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5092 2582 5120 2926
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5368 2514 5396 2926
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5460 2310 5488 2382
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 4622 2204 4918 2224
rect 4678 2202 4702 2204
rect 4758 2202 4782 2204
rect 4838 2202 4862 2204
rect 4700 2150 4702 2202
rect 4764 2150 4776 2202
rect 4838 2150 4840 2202
rect 4678 2148 4702 2150
rect 4758 2148 4782 2150
rect 4838 2148 4862 2150
rect 4622 2128 4918 2148
rect 4526 82 4582 480
rect 4264 54 4582 82
rect 5552 82 5580 3674
rect 5644 3505 5672 10406
rect 6012 10198 6040 10950
rect 6288 10810 6316 11018
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6288 10606 6316 10746
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6012 9178 6040 10134
rect 6288 9722 6316 10134
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6564 9178 6592 10950
rect 6656 10810 6684 11154
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10713 6684 10746
rect 6642 10704 6698 10713
rect 7116 10674 7144 11290
rect 7576 11218 7604 13767
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 6642 10639 6698 10648
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6932 10266 6960 10474
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6748 9110 6776 9590
rect 6932 9586 6960 10202
rect 7024 10198 7052 10474
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9586 7236 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 7208 8906 7236 9522
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 5736 7002 5764 8366
rect 6288 8022 6316 8366
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7478 5856 7890
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6118 6224 6734
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5846 6224 6054
rect 6288 5953 6316 7414
rect 6472 6866 6500 7822
rect 6564 7206 6592 8230
rect 7208 7886 7236 8842
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7342 6684 7686
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6840 6934 6868 7278
rect 7300 7002 7328 7958
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6288 5778 6316 5879
rect 6472 5778 6500 6802
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6748 5846 6776 6734
rect 7392 6254 7420 11018
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10198 7604 10610
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7576 9722 7604 10134
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7760 9382 7788 10134
rect 7944 10062 7972 10542
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8430 7604 8774
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7760 7546 7788 9318
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7852 7206 7880 7890
rect 7944 7818 7972 9998
rect 8036 9654 8064 18022
rect 8289 17980 8585 18000
rect 8345 17978 8369 17980
rect 8425 17978 8449 17980
rect 8505 17978 8529 17980
rect 8367 17926 8369 17978
rect 8431 17926 8443 17978
rect 8505 17926 8507 17978
rect 8345 17924 8369 17926
rect 8425 17924 8449 17926
rect 8505 17924 8529 17926
rect 8289 17904 8585 17924
rect 8289 16892 8585 16912
rect 8345 16890 8369 16892
rect 8425 16890 8449 16892
rect 8505 16890 8529 16892
rect 8367 16838 8369 16890
rect 8431 16838 8443 16890
rect 8505 16838 8507 16890
rect 8345 16836 8369 16838
rect 8425 16836 8449 16838
rect 8505 16836 8529 16838
rect 8289 16816 8585 16836
rect 8289 15804 8585 15824
rect 8345 15802 8369 15804
rect 8425 15802 8449 15804
rect 8505 15802 8529 15804
rect 8367 15750 8369 15802
rect 8431 15750 8443 15802
rect 8505 15750 8507 15802
rect 8345 15748 8369 15750
rect 8425 15748 8449 15750
rect 8505 15748 8529 15750
rect 8289 15728 8585 15748
rect 8289 14716 8585 14736
rect 8345 14714 8369 14716
rect 8425 14714 8449 14716
rect 8505 14714 8529 14716
rect 8367 14662 8369 14714
rect 8431 14662 8443 14714
rect 8505 14662 8507 14714
rect 8345 14660 8369 14662
rect 8425 14660 8449 14662
rect 8505 14660 8529 14662
rect 8289 14640 8585 14660
rect 8289 13628 8585 13648
rect 8345 13626 8369 13628
rect 8425 13626 8449 13628
rect 8505 13626 8529 13628
rect 8367 13574 8369 13626
rect 8431 13574 8443 13626
rect 8505 13574 8507 13626
rect 8345 13572 8369 13574
rect 8425 13572 8449 13574
rect 8505 13572 8529 13574
rect 8289 13552 8585 13572
rect 8289 12540 8585 12560
rect 8345 12538 8369 12540
rect 8425 12538 8449 12540
rect 8505 12538 8529 12540
rect 8367 12486 8369 12538
rect 8431 12486 8443 12538
rect 8505 12486 8507 12538
rect 8345 12484 8369 12486
rect 8425 12484 8449 12486
rect 8505 12484 8529 12486
rect 8289 12464 8585 12484
rect 8289 11452 8585 11472
rect 8345 11450 8369 11452
rect 8425 11450 8449 11452
rect 8505 11450 8529 11452
rect 8367 11398 8369 11450
rect 8431 11398 8443 11450
rect 8505 11398 8507 11450
rect 8345 11396 8369 11398
rect 8425 11396 8449 11398
rect 8505 11396 8529 11398
rect 8289 11376 8585 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10470 8248 11154
rect 8680 11082 8708 21490
rect 9232 21459 9260 21490
rect 9692 11558 9720 21490
rect 10980 21459 11008 21490
rect 11956 19612 12252 19632
rect 12012 19610 12036 19612
rect 12092 19610 12116 19612
rect 12172 19610 12196 19612
rect 12034 19558 12036 19610
rect 12098 19558 12110 19610
rect 12172 19558 12174 19610
rect 12012 19556 12036 19558
rect 12092 19556 12116 19558
rect 12172 19556 12196 19558
rect 11956 19536 12252 19556
rect 11956 18524 12252 18544
rect 12012 18522 12036 18524
rect 12092 18522 12116 18524
rect 12172 18522 12196 18524
rect 12034 18470 12036 18522
rect 12098 18470 12110 18522
rect 12172 18470 12174 18522
rect 12012 18468 12036 18470
rect 12092 18468 12116 18470
rect 12172 18468 12196 18470
rect 11956 18448 12252 18468
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8289 10364 8585 10384
rect 8345 10362 8369 10364
rect 8425 10362 8449 10364
rect 8505 10362 8529 10364
rect 8367 10310 8369 10362
rect 8431 10310 8443 10362
rect 8505 10310 8507 10362
rect 8345 10308 8369 10310
rect 8425 10308 8449 10310
rect 8505 10308 8529 10310
rect 8289 10288 8585 10308
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8289 9276 8585 9296
rect 8345 9274 8369 9276
rect 8425 9274 8449 9276
rect 8505 9274 8529 9276
rect 8367 9222 8369 9274
rect 8431 9222 8443 9274
rect 8505 9222 8507 9274
rect 8345 9220 8369 9222
rect 8425 9220 8449 9222
rect 8505 9220 8529 9222
rect 8289 9200 8585 9220
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8634 8064 9046
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8289 8188 8585 8208
rect 8345 8186 8369 8188
rect 8425 8186 8449 8188
rect 8505 8186 8529 8188
rect 8367 8134 8369 8186
rect 8431 8134 8443 8186
rect 8505 8134 8507 8186
rect 8345 8132 8369 8134
rect 8425 8132 8449 8134
rect 8505 8132 8529 8134
rect 8289 8112 8585 8132
rect 8772 7954 8800 8298
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 7002 7880 7142
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7852 6118 7880 6938
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4690 6408 5102
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5736 3602 5764 4558
rect 5920 4282 5948 4626
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5630 3496 5686 3505
rect 5630 3431 5686 3440
rect 5736 3194 5764 3538
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5632 2984 5684 2990
rect 5828 2972 5856 3538
rect 5920 3466 5948 3946
rect 6380 3602 6408 4626
rect 6564 3942 6592 4966
rect 6656 4758 6684 5170
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6748 4146 6776 5238
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5684 2944 5856 2972
rect 5632 2926 5684 2932
rect 5644 2854 5672 2926
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2514 5672 2790
rect 6196 2514 6224 3470
rect 6564 2582 6592 3878
rect 6840 3738 6868 4422
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6932 3058 6960 3130
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6932 2417 6960 2450
rect 6918 2408 6974 2417
rect 6918 2343 6974 2352
rect 5814 82 5870 480
rect 5552 54 5870 82
rect 7024 82 7052 6054
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 4826 7144 5510
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7208 4758 7236 5646
rect 7852 5098 7880 6054
rect 7944 5710 7972 7754
rect 8289 7100 8585 7120
rect 8345 7098 8369 7100
rect 8425 7098 8449 7100
rect 8505 7098 8529 7100
rect 8367 7046 8369 7098
rect 8431 7046 8443 7098
rect 8505 7046 8507 7098
rect 8345 7044 8369 7046
rect 8425 7044 8449 7046
rect 8505 7044 8529 7046
rect 8289 7024 8585 7044
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8036 5370 8064 6326
rect 8128 6254 8156 6666
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5642 8156 6190
rect 8289 6012 8585 6032
rect 8345 6010 8369 6012
rect 8425 6010 8449 6012
rect 8505 6010 8529 6012
rect 8367 5958 8369 6010
rect 8431 5958 8443 6010
rect 8505 5958 8507 6010
rect 8345 5956 8369 5958
rect 8425 5956 8449 5958
rect 8505 5956 8529 5958
rect 8289 5936 8585 5956
rect 8680 5846 8708 6598
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8772 5370 8800 6122
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7760 4758 7788 4966
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7576 4622 7604 4694
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7852 3942 7880 4762
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7760 3738 7788 3878
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3641 7880 3878
rect 7838 3632 7894 3641
rect 7838 3567 7894 3576
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3058 7696 3470
rect 7852 3058 7880 3567
rect 8036 3534 8064 4490
rect 8128 3942 8156 4966
rect 8220 4214 8248 5102
rect 8772 5098 8800 5306
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8289 4924 8585 4944
rect 8345 4922 8369 4924
rect 8425 4922 8449 4924
rect 8505 4922 8529 4924
rect 8367 4870 8369 4922
rect 8431 4870 8443 4922
rect 8505 4870 8507 4922
rect 8345 4868 8369 4870
rect 8425 4868 8449 4870
rect 8505 4868 8529 4870
rect 8289 4848 8585 4868
rect 8574 4584 8630 4593
rect 8574 4519 8630 4528
rect 8760 4548 8812 4554
rect 8588 4486 8616 4519
rect 8760 4490 8812 4496
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8680 4049 8708 4082
rect 8666 4040 8722 4049
rect 8772 4010 8800 4490
rect 8666 3975 8722 3984
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3584 8156 3878
rect 8289 3836 8585 3856
rect 8345 3834 8369 3836
rect 8425 3834 8449 3836
rect 8505 3834 8529 3836
rect 8367 3782 8369 3834
rect 8431 3782 8443 3834
rect 8505 3782 8507 3834
rect 8345 3780 8369 3782
rect 8425 3780 8449 3782
rect 8505 3780 8529 3782
rect 8289 3760 8585 3780
rect 8772 3670 8800 3946
rect 8760 3664 8812 3670
rect 8864 3641 8892 10406
rect 9048 9042 9076 11494
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 9586 9352 10950
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10266 10364 10406
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 9178 9352 9522
rect 9692 9450 9720 9998
rect 10244 9722 10272 10066
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9968 9110 9996 9386
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 7750 8984 8434
rect 9048 8294 9076 8978
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7410 8984 7686
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9048 4154 9076 8230
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7546 9168 7822
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 5166 9168 6598
rect 9232 6390 9260 7686
rect 9324 7274 9352 8774
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9324 7002 9352 7210
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9416 6458 9444 7210
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9232 4758 9260 6326
rect 9692 5846 9720 8842
rect 10244 8634 10272 9658
rect 10888 9586 10916 10202
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10980 9110 11008 9386
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10244 8294 10272 8570
rect 10520 8566 10548 9046
rect 10612 8634 10640 9046
rect 11164 9042 11192 9522
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11256 8634 11284 9862
rect 11532 9382 11560 10066
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10612 8090 10640 8570
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11164 8090 11192 8502
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10888 7410 10916 7958
rect 11256 7410 11284 8366
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10612 6798 10640 7210
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9784 6225 9812 6258
rect 10060 6254 10088 6598
rect 10048 6248 10100 6254
rect 9770 6216 9826 6225
rect 10048 6190 10100 6196
rect 9770 6151 9826 6160
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5302 9352 5510
rect 9692 5302 9720 5782
rect 10244 5370 10272 5850
rect 10612 5846 10640 6734
rect 10704 6254 10732 6870
rect 10980 6322 11008 7210
rect 11256 6934 11284 7346
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 11348 5914 11376 6802
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 11440 5710 11468 6054
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9692 4758 9720 5034
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 8944 4140 8996 4146
rect 9048 4126 9168 4154
rect 8944 4082 8996 4088
rect 8760 3606 8812 3612
rect 8850 3632 8906 3641
rect 8208 3596 8260 3602
rect 8128 3556 8208 3584
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7932 2916 7984 2922
rect 7932 2858 7984 2864
rect 7116 2514 7144 2858
rect 7944 2582 7972 2858
rect 8128 2854 8156 3556
rect 8850 3567 8906 3576
rect 8208 3538 8260 3544
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 2990 8248 3402
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 2582 8156 2790
rect 8220 2650 8248 2926
rect 8864 2854 8892 3567
rect 8956 3369 8984 4082
rect 8942 3360 8998 3369
rect 8942 3295 8998 3304
rect 8956 3194 8984 3295
rect 9140 3194 9168 4126
rect 9692 3942 9720 4694
rect 10336 4010 10364 5510
rect 10980 5098 11008 5646
rect 11440 5370 11468 5646
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4690 10640 4966
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10980 4282 11008 5034
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11164 4214 11192 5170
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11348 4622 11376 4762
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11256 4049 11284 4422
rect 11242 4040 11298 4049
rect 10324 4004 10376 4010
rect 11242 3975 11298 3984
rect 10324 3946 10376 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9692 2922 9720 3878
rect 11348 3738 11376 4558
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9956 3120 10008 3126
rect 9876 3080 9956 3108
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8289 2748 8585 2768
rect 8345 2746 8369 2748
rect 8425 2746 8449 2748
rect 8505 2746 8529 2748
rect 8367 2694 8369 2746
rect 8431 2694 8443 2746
rect 8505 2694 8507 2746
rect 8345 2692 8369 2694
rect 8425 2692 8449 2694
rect 8505 2692 8529 2694
rect 8289 2672 8585 2692
rect 9876 2650 9904 3080
rect 9956 3062 10008 3068
rect 10060 3058 10088 3606
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 2310 9260 2450
rect 10060 2446 10088 2518
rect 10520 2514 10548 3402
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10704 2514 10732 3130
rect 10796 2990 10824 3334
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10888 2650 10916 3130
rect 10980 2990 11008 3674
rect 11244 3460 11296 3466
rect 11440 3448 11468 4422
rect 11296 3420 11468 3448
rect 11244 3402 11296 3408
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 11256 2446 11284 2790
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9232 2106 9260 2246
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 7102 82 7158 480
rect 7024 54 7158 82
rect 662 0 718 54
rect 1950 0 2006 54
rect 3238 0 3294 54
rect 4526 0 4582 54
rect 5814 0 5870 54
rect 7102 0 7158 54
rect 8390 128 8446 480
rect 8390 76 8392 128
rect 8444 76 8446 128
rect 8390 0 8446 76
rect 9600 82 9628 2246
rect 9678 82 9734 480
rect 9600 54 9734 82
rect 9678 0 9734 54
rect 10966 82 11022 480
rect 11348 82 11376 2586
rect 11532 2106 11560 9318
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7478 11744 7890
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11716 7206 11744 7414
rect 11808 7324 11836 18158
rect 11956 17436 12252 17456
rect 12012 17434 12036 17436
rect 12092 17434 12116 17436
rect 12172 17434 12196 17436
rect 12034 17382 12036 17434
rect 12098 17382 12110 17434
rect 12172 17382 12174 17434
rect 12012 17380 12036 17382
rect 12092 17380 12116 17382
rect 12172 17380 12196 17382
rect 11956 17360 12252 17380
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 11956 16348 12252 16368
rect 12012 16346 12036 16348
rect 12092 16346 12116 16348
rect 12172 16346 12196 16348
rect 12034 16294 12036 16346
rect 12098 16294 12110 16346
rect 12172 16294 12174 16346
rect 12012 16292 12036 16294
rect 12092 16292 12116 16294
rect 12172 16292 12196 16294
rect 11956 16272 12252 16292
rect 11956 15260 12252 15280
rect 12012 15258 12036 15260
rect 12092 15258 12116 15260
rect 12172 15258 12196 15260
rect 12034 15206 12036 15258
rect 12098 15206 12110 15258
rect 12172 15206 12174 15258
rect 12012 15204 12036 15206
rect 12092 15204 12116 15206
rect 12172 15204 12196 15206
rect 11956 15184 12252 15204
rect 11956 14172 12252 14192
rect 12012 14170 12036 14172
rect 12092 14170 12116 14172
rect 12172 14170 12196 14172
rect 12034 14118 12036 14170
rect 12098 14118 12110 14170
rect 12172 14118 12174 14170
rect 12012 14116 12036 14118
rect 12092 14116 12116 14118
rect 12172 14116 12196 14118
rect 11956 14096 12252 14116
rect 11956 13084 12252 13104
rect 12012 13082 12036 13084
rect 12092 13082 12116 13084
rect 12172 13082 12196 13084
rect 12034 13030 12036 13082
rect 12098 13030 12110 13082
rect 12172 13030 12174 13082
rect 12012 13028 12036 13030
rect 12092 13028 12116 13030
rect 12172 13028 12196 13030
rect 11956 13008 12252 13028
rect 11956 11996 12252 12016
rect 12012 11994 12036 11996
rect 12092 11994 12116 11996
rect 12172 11994 12196 11996
rect 12034 11942 12036 11994
rect 12098 11942 12110 11994
rect 12172 11942 12174 11994
rect 12012 11940 12036 11942
rect 12092 11940 12116 11942
rect 12172 11940 12196 11942
rect 11956 11920 12252 11940
rect 11956 10908 12252 10928
rect 12012 10906 12036 10908
rect 12092 10906 12116 10908
rect 12172 10906 12196 10908
rect 12034 10854 12036 10906
rect 12098 10854 12110 10906
rect 12172 10854 12174 10906
rect 12012 10852 12036 10854
rect 12092 10852 12116 10854
rect 12172 10852 12196 10854
rect 11956 10832 12252 10852
rect 12164 10124 12216 10130
rect 12360 10112 12388 17070
rect 12452 11218 12480 21542
rect 12622 21520 12678 21542
rect 14370 21570 14426 22000
rect 14370 21542 14504 21570
rect 14370 21520 14426 21542
rect 14476 18426 14504 21542
rect 15200 21548 15252 21554
rect 16026 21548 16082 22000
rect 16026 21520 16028 21548
rect 15200 21490 15252 21496
rect 16080 21520 16082 21548
rect 16580 21548 16632 21554
rect 16028 21490 16080 21496
rect 17682 21548 17738 22000
rect 17682 21520 17684 21548
rect 16580 21490 16632 21496
rect 17736 21520 17738 21548
rect 19430 21570 19486 22000
rect 19430 21542 19656 21570
rect 19430 21520 19486 21542
rect 17684 21490 17736 21496
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12636 11257 12664 11290
rect 12622 11248 12678 11257
rect 12440 11212 12492 11218
rect 12622 11183 12678 11192
rect 12440 11154 12492 11160
rect 12452 10810 12480 11154
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12530 10568 12586 10577
rect 12452 10538 12530 10554
rect 12440 10532 12530 10538
rect 12492 10526 12530 10532
rect 12530 10503 12586 10512
rect 12440 10474 12492 10480
rect 15212 10266 15240 21490
rect 16040 21459 16068 21490
rect 15622 19068 15918 19088
rect 15678 19066 15702 19068
rect 15758 19066 15782 19068
rect 15838 19066 15862 19068
rect 15700 19014 15702 19066
rect 15764 19014 15776 19066
rect 15838 19014 15840 19066
rect 15678 19012 15702 19014
rect 15758 19012 15782 19014
rect 15838 19012 15862 19014
rect 15622 18992 15918 19012
rect 15622 17980 15918 18000
rect 15678 17978 15702 17980
rect 15758 17978 15782 17980
rect 15838 17978 15862 17980
rect 15700 17926 15702 17978
rect 15764 17926 15776 17978
rect 15838 17926 15840 17978
rect 15678 17924 15702 17926
rect 15758 17924 15782 17926
rect 15838 17924 15862 17926
rect 15622 17904 15918 17924
rect 15622 16892 15918 16912
rect 15678 16890 15702 16892
rect 15758 16890 15782 16892
rect 15838 16890 15862 16892
rect 15700 16838 15702 16890
rect 15764 16838 15776 16890
rect 15838 16838 15840 16890
rect 15678 16836 15702 16838
rect 15758 16836 15782 16838
rect 15838 16836 15862 16838
rect 15622 16816 15918 16836
rect 15622 15804 15918 15824
rect 15678 15802 15702 15804
rect 15758 15802 15782 15804
rect 15838 15802 15862 15804
rect 15700 15750 15702 15802
rect 15764 15750 15776 15802
rect 15838 15750 15840 15802
rect 15678 15748 15702 15750
rect 15758 15748 15782 15750
rect 15838 15748 15862 15750
rect 15622 15728 15918 15748
rect 15622 14716 15918 14736
rect 15678 14714 15702 14716
rect 15758 14714 15782 14716
rect 15838 14714 15862 14716
rect 15700 14662 15702 14714
rect 15764 14662 15776 14714
rect 15838 14662 15840 14714
rect 15678 14660 15702 14662
rect 15758 14660 15782 14662
rect 15838 14660 15862 14662
rect 15622 14640 15918 14660
rect 15622 13628 15918 13648
rect 15678 13626 15702 13628
rect 15758 13626 15782 13628
rect 15838 13626 15862 13628
rect 15700 13574 15702 13626
rect 15764 13574 15776 13626
rect 15838 13574 15840 13626
rect 15678 13572 15702 13574
rect 15758 13572 15782 13574
rect 15838 13572 15862 13574
rect 15622 13552 15918 13572
rect 15622 12540 15918 12560
rect 15678 12538 15702 12540
rect 15758 12538 15782 12540
rect 15838 12538 15862 12540
rect 15700 12486 15702 12538
rect 15764 12486 15776 12538
rect 15838 12486 15840 12538
rect 15678 12484 15702 12486
rect 15758 12484 15782 12486
rect 15838 12484 15862 12486
rect 15622 12464 15918 12484
rect 15622 11452 15918 11472
rect 15678 11450 15702 11452
rect 15758 11450 15782 11452
rect 15838 11450 15862 11452
rect 15700 11398 15702 11450
rect 15764 11398 15776 11450
rect 15838 11398 15840 11450
rect 15678 11396 15702 11398
rect 15758 11396 15782 11398
rect 15838 11396 15862 11398
rect 15622 11376 15918 11396
rect 15382 10704 15438 10713
rect 15382 10639 15438 10648
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15396 10130 15424 10639
rect 15622 10364 15918 10384
rect 15678 10362 15702 10364
rect 15758 10362 15782 10364
rect 15838 10362 15862 10364
rect 15700 10310 15702 10362
rect 15764 10310 15776 10362
rect 15838 10310 15840 10362
rect 15678 10308 15702 10310
rect 15758 10308 15782 10310
rect 15838 10308 15862 10310
rect 15622 10288 15918 10308
rect 12216 10084 12388 10112
rect 12532 10124 12584 10130
rect 12164 10066 12216 10072
rect 12532 10066 12584 10072
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 11956 9820 12252 9840
rect 12012 9818 12036 9820
rect 12092 9818 12116 9820
rect 12172 9818 12196 9820
rect 12034 9766 12036 9818
rect 12098 9766 12110 9818
rect 12172 9766 12174 9818
rect 12012 9764 12036 9766
rect 12092 9764 12116 9766
rect 12172 9764 12196 9766
rect 11956 9744 12252 9764
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 11956 8732 12252 8752
rect 12012 8730 12036 8732
rect 12092 8730 12116 8732
rect 12172 8730 12196 8732
rect 12034 8678 12036 8730
rect 12098 8678 12110 8730
rect 12172 8678 12174 8730
rect 12012 8676 12036 8678
rect 12092 8676 12116 8678
rect 12172 8676 12196 8678
rect 11956 8656 12252 8676
rect 12360 8634 12388 8978
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11900 7478 11928 7754
rect 11956 7644 12252 7664
rect 12012 7642 12036 7644
rect 12092 7642 12116 7644
rect 12172 7642 12196 7644
rect 12034 7590 12036 7642
rect 12098 7590 12110 7642
rect 12172 7590 12174 7642
rect 12012 7588 12036 7590
rect 12092 7588 12116 7590
rect 12172 7588 12196 7590
rect 11956 7568 12252 7588
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11808 7296 11928 7324
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11624 5030 11652 5782
rect 11716 5710 11744 6598
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11716 5234 11744 5646
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11808 4842 11836 5510
rect 11900 5137 11928 7296
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 11956 6556 12252 6576
rect 12012 6554 12036 6556
rect 12092 6554 12116 6556
rect 12172 6554 12196 6556
rect 12034 6502 12036 6554
rect 12098 6502 12110 6554
rect 12172 6502 12174 6554
rect 12012 6500 12036 6502
rect 12092 6500 12116 6502
rect 12172 6500 12196 6502
rect 11956 6480 12252 6500
rect 12360 6458 12388 6802
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12452 5778 12480 9590
rect 12544 9586 12572 10066
rect 12714 9616 12770 9625
rect 12532 9580 12584 9586
rect 12714 9551 12770 9560
rect 12532 9522 12584 9528
rect 12728 8430 12756 9551
rect 15396 9382 15424 10066
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 12716 8424 12768 8430
rect 12622 8392 12678 8401
rect 12716 8366 12768 8372
rect 12622 8327 12678 8336
rect 12636 7546 12664 8327
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12544 5914 12572 6190
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11956 5468 12252 5488
rect 12012 5466 12036 5468
rect 12092 5466 12116 5468
rect 12172 5466 12196 5468
rect 12034 5414 12036 5466
rect 12098 5414 12110 5466
rect 12172 5414 12174 5466
rect 12012 5412 12036 5414
rect 12092 5412 12116 5414
rect 12172 5412 12196 5414
rect 11956 5392 12252 5412
rect 11886 5128 11942 5137
rect 11886 5063 11942 5072
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11716 4814 11928 4842
rect 11716 4622 11744 4814
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11808 4010 11836 4694
rect 11900 4146 11928 4814
rect 11992 4622 12020 5034
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11956 4380 12252 4400
rect 12012 4378 12036 4380
rect 12092 4378 12116 4380
rect 12172 4378 12196 4380
rect 12034 4326 12036 4378
rect 12098 4326 12110 4378
rect 12172 4326 12174 4378
rect 12012 4324 12036 4326
rect 12092 4324 12116 4326
rect 12172 4324 12196 4326
rect 11956 4304 12252 4324
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 12348 3936 12400 3942
rect 12452 3924 12480 5034
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12544 4078 12572 4218
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12400 3896 12480 3924
rect 12348 3878 12400 3884
rect 12544 3738 12572 4014
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12636 3670 12664 7142
rect 12900 5908 12952 5914
rect 12952 5868 13032 5896
rect 12900 5850 12952 5856
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12912 5234 12940 5714
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 13004 4486 13032 5868
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4214 13032 4422
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 11624 3194 11652 3606
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 12624 3460 12676 3466
rect 12728 3448 12756 3674
rect 12676 3420 12756 3448
rect 12990 3496 13046 3505
rect 12990 3431 13046 3440
rect 12624 3402 12676 3408
rect 11808 3369 11836 3402
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 11956 3292 12252 3312
rect 12012 3290 12036 3292
rect 12092 3290 12116 3292
rect 12172 3290 12196 3292
rect 12034 3238 12036 3290
rect 12098 3238 12110 3290
rect 12172 3238 12174 3290
rect 12012 3236 12036 3238
rect 12092 3236 12116 3238
rect 12172 3236 12196 3238
rect 11956 3216 12252 3236
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 12636 3058 12664 3402
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3126 12848 3334
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 13004 3058 13032 3431
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12268 2417 12296 2450
rect 12254 2408 12310 2417
rect 12254 2343 12310 2352
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 11956 2204 12252 2224
rect 12012 2202 12036 2204
rect 12092 2202 12116 2204
rect 12172 2202 12196 2204
rect 12034 2150 12036 2202
rect 12098 2150 12110 2202
rect 12172 2150 12174 2202
rect 12012 2148 12036 2150
rect 12092 2148 12116 2150
rect 12172 2148 12196 2150
rect 11956 2128 12252 2148
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 11532 105 11560 2042
rect 10966 54 11376 82
rect 11518 96 11574 105
rect 10966 0 11022 54
rect 11518 31 11574 40
rect 12254 82 12310 480
rect 12636 82 12664 2042
rect 12820 134 12848 2246
rect 13096 2106 13124 7142
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13740 6118 13768 6802
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5681 13768 6054
rect 15396 5681 15424 9318
rect 15622 9276 15918 9296
rect 15678 9274 15702 9276
rect 15758 9274 15782 9276
rect 15838 9274 15862 9276
rect 15700 9222 15702 9274
rect 15764 9222 15776 9274
rect 15838 9222 15840 9274
rect 15678 9220 15702 9222
rect 15758 9220 15782 9222
rect 15838 9220 15862 9222
rect 15622 9200 15918 9220
rect 15622 8188 15918 8208
rect 15678 8186 15702 8188
rect 15758 8186 15782 8188
rect 15838 8186 15862 8188
rect 15700 8134 15702 8186
rect 15764 8134 15776 8186
rect 15838 8134 15840 8186
rect 15678 8132 15702 8134
rect 15758 8132 15782 8134
rect 15838 8132 15862 8134
rect 15622 8112 15918 8132
rect 15622 7100 15918 7120
rect 15678 7098 15702 7100
rect 15758 7098 15782 7100
rect 15838 7098 15862 7100
rect 15700 7046 15702 7098
rect 15764 7046 15776 7098
rect 15838 7046 15840 7098
rect 15678 7044 15702 7046
rect 15758 7044 15782 7046
rect 15838 7044 15862 7046
rect 15622 7024 15918 7044
rect 16592 6225 16620 21490
rect 17696 21459 17724 21490
rect 17222 20360 17278 20369
rect 17222 20295 17278 20304
rect 17236 10198 17264 20295
rect 19289 19612 19585 19632
rect 19345 19610 19369 19612
rect 19425 19610 19449 19612
rect 19505 19610 19529 19612
rect 19367 19558 19369 19610
rect 19431 19558 19443 19610
rect 19505 19558 19507 19610
rect 19345 19556 19369 19558
rect 19425 19556 19449 19558
rect 19505 19556 19529 19558
rect 19289 19536 19585 19556
rect 19289 18524 19585 18544
rect 19345 18522 19369 18524
rect 19425 18522 19449 18524
rect 19505 18522 19529 18524
rect 19367 18470 19369 18522
rect 19431 18470 19443 18522
rect 19505 18470 19507 18522
rect 19345 18468 19369 18470
rect 19425 18468 19449 18470
rect 19505 18468 19529 18470
rect 19289 18448 19585 18468
rect 19289 17436 19585 17456
rect 19345 17434 19369 17436
rect 19425 17434 19449 17436
rect 19505 17434 19529 17436
rect 19367 17382 19369 17434
rect 19431 17382 19443 17434
rect 19505 17382 19507 17434
rect 19345 17380 19369 17382
rect 19425 17380 19449 17382
rect 19505 17380 19529 17382
rect 19289 17360 19585 17380
rect 19289 16348 19585 16368
rect 19345 16346 19369 16348
rect 19425 16346 19449 16348
rect 19505 16346 19529 16348
rect 19367 16294 19369 16346
rect 19431 16294 19443 16346
rect 19505 16294 19507 16346
rect 19345 16292 19369 16294
rect 19425 16292 19449 16294
rect 19505 16292 19529 16294
rect 19289 16272 19585 16292
rect 19062 15464 19118 15473
rect 19062 15399 19118 15408
rect 19076 14482 19104 15399
rect 19289 15260 19585 15280
rect 19345 15258 19369 15260
rect 19425 15258 19449 15260
rect 19505 15258 19529 15260
rect 19367 15206 19369 15258
rect 19431 15206 19443 15258
rect 19505 15206 19507 15258
rect 19345 15204 19369 15206
rect 19425 15204 19449 15206
rect 19505 15204 19529 15206
rect 19289 15184 19585 15204
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 14074 19104 14418
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19168 13705 19196 14214
rect 19289 14172 19585 14192
rect 19345 14170 19369 14172
rect 19425 14170 19449 14172
rect 19505 14170 19529 14172
rect 19367 14118 19369 14170
rect 19431 14118 19443 14170
rect 19505 14118 19507 14170
rect 19345 14116 19369 14118
rect 19425 14116 19449 14118
rect 19505 14116 19529 14118
rect 19289 14096 19585 14116
rect 19154 13696 19210 13705
rect 19154 13631 19210 13640
rect 19289 13084 19585 13104
rect 19345 13082 19369 13084
rect 19425 13082 19449 13084
rect 19505 13082 19529 13084
rect 19367 13030 19369 13082
rect 19431 13030 19443 13082
rect 19505 13030 19507 13082
rect 19345 13028 19369 13030
rect 19425 13028 19449 13030
rect 19505 13028 19529 13030
rect 19289 13008 19585 13028
rect 19289 11996 19585 12016
rect 19345 11994 19369 11996
rect 19425 11994 19449 11996
rect 19505 11994 19529 11996
rect 19367 11942 19369 11994
rect 19431 11942 19443 11994
rect 19505 11942 19507 11994
rect 19345 11940 19369 11942
rect 19425 11940 19449 11942
rect 19505 11940 19529 11942
rect 19289 11920 19585 11940
rect 19289 10908 19585 10928
rect 19345 10906 19369 10908
rect 19425 10906 19449 10908
rect 19505 10906 19529 10908
rect 19367 10854 19369 10906
rect 19431 10854 19443 10906
rect 19505 10854 19507 10906
rect 19345 10852 19369 10854
rect 19425 10852 19449 10854
rect 19505 10852 19529 10854
rect 19289 10832 19585 10852
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 19289 9820 19585 9840
rect 19345 9818 19369 9820
rect 19425 9818 19449 9820
rect 19505 9818 19529 9820
rect 19367 9766 19369 9818
rect 19431 9766 19443 9818
rect 19505 9766 19507 9818
rect 19345 9764 19369 9766
rect 19425 9764 19449 9766
rect 19505 9764 19529 9766
rect 19289 9744 19585 9764
rect 19628 9625 19656 21542
rect 19708 21548 19760 21554
rect 21086 21548 21142 22000
rect 21086 21520 21088 21548
rect 19708 21490 19760 21496
rect 21140 21520 21142 21548
rect 21088 21490 21140 21496
rect 19720 10577 19748 21490
rect 21100 21459 21128 21490
rect 19890 17912 19946 17921
rect 19890 17847 19946 17856
rect 19904 17338 19932 17847
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19706 10568 19762 10577
rect 19706 10503 19762 10512
rect 19614 9616 19670 9625
rect 19614 9551 19670 9560
rect 19289 8732 19585 8752
rect 19345 8730 19369 8732
rect 19425 8730 19449 8732
rect 19505 8730 19529 8732
rect 19367 8678 19369 8730
rect 19431 8678 19443 8730
rect 19505 8678 19507 8730
rect 19345 8676 19369 8678
rect 19425 8676 19449 8678
rect 19505 8676 19529 8678
rect 19289 8656 19585 8676
rect 19289 7644 19585 7664
rect 19345 7642 19369 7644
rect 19425 7642 19449 7644
rect 19505 7642 19529 7644
rect 19367 7590 19369 7642
rect 19431 7590 19443 7642
rect 19505 7590 19507 7642
rect 19345 7588 19369 7590
rect 19425 7588 19449 7590
rect 19505 7588 19529 7590
rect 19289 7568 19585 7588
rect 19289 6556 19585 6576
rect 19345 6554 19369 6556
rect 19425 6554 19449 6556
rect 19505 6554 19529 6556
rect 19367 6502 19369 6554
rect 19431 6502 19443 6554
rect 19505 6502 19507 6554
rect 19345 6500 19369 6502
rect 19425 6500 19449 6502
rect 19505 6500 19529 6502
rect 19289 6480 19585 6500
rect 16578 6216 16634 6225
rect 16578 6151 16634 6160
rect 15622 6012 15918 6032
rect 15678 6010 15702 6012
rect 15758 6010 15782 6012
rect 15838 6010 15862 6012
rect 15700 5958 15702 6010
rect 15764 5958 15776 6010
rect 15838 5958 15840 6010
rect 15678 5956 15702 5958
rect 15758 5956 15782 5958
rect 15838 5956 15862 5958
rect 15622 5936 15918 5956
rect 13726 5672 13782 5681
rect 13726 5607 13782 5616
rect 15382 5672 15438 5681
rect 15382 5607 15438 5616
rect 19289 5468 19585 5488
rect 19345 5466 19369 5468
rect 19425 5466 19449 5468
rect 19505 5466 19529 5468
rect 19367 5414 19369 5466
rect 19431 5414 19443 5466
rect 19505 5414 19507 5466
rect 19345 5412 19369 5414
rect 19425 5412 19449 5414
rect 19505 5412 19529 5414
rect 19289 5392 19585 5412
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13188 3602 13216 4218
rect 13372 4154 13400 5170
rect 13556 5137 13584 5170
rect 13542 5128 13598 5137
rect 13542 5063 13598 5072
rect 15622 4924 15918 4944
rect 15678 4922 15702 4924
rect 15758 4922 15782 4924
rect 15838 4922 15862 4924
rect 15700 4870 15702 4922
rect 15764 4870 15776 4922
rect 15838 4870 15840 4922
rect 15678 4868 15702 4870
rect 15758 4868 15782 4870
rect 15838 4868 15862 4870
rect 15622 4848 15918 4868
rect 13450 4720 13506 4729
rect 13450 4655 13452 4664
rect 13504 4655 13506 4664
rect 13636 4684 13688 4690
rect 13452 4626 13504 4632
rect 13636 4626 13688 4632
rect 13464 4282 13492 4626
rect 13648 4593 13676 4626
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 13820 4548 13872 4554
rect 13648 4282 13676 4519
rect 13820 4490 13872 4496
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13372 4126 13492 4154
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 2582 13400 3334
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 12254 54 12664 82
rect 12808 128 12860 134
rect 12808 70 12860 76
rect 13464 82 13492 4126
rect 13832 4078 13860 4490
rect 19289 4380 19585 4400
rect 19345 4378 19369 4380
rect 19425 4378 19449 4380
rect 19505 4378 19529 4380
rect 19367 4326 19369 4378
rect 19431 4326 19443 4378
rect 19505 4326 19507 4378
rect 19345 4324 19369 4326
rect 19425 4324 19449 4326
rect 19505 4324 19529 4326
rect 19289 4304 19585 4324
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 15622 3836 15918 3856
rect 15678 3834 15702 3836
rect 15758 3834 15782 3836
rect 15838 3834 15862 3836
rect 15700 3782 15702 3834
rect 15764 3782 15776 3834
rect 15838 3782 15840 3834
rect 15678 3780 15702 3782
rect 15758 3780 15782 3782
rect 15838 3780 15862 3782
rect 15622 3760 15918 3780
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 13556 3194 13584 3538
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 3194 13676 3402
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 14016 2854 14044 3470
rect 15212 2854 15240 3538
rect 17130 3496 17186 3505
rect 17130 3431 17186 3440
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14016 2650 14044 2790
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14568 2310 14596 2790
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 13542 82 13598 480
rect 13464 54 13598 82
rect 14568 82 14596 2246
rect 15488 2106 15516 2926
rect 15622 2748 15918 2768
rect 15678 2746 15702 2748
rect 15758 2746 15782 2748
rect 15838 2746 15862 2748
rect 15700 2694 15702 2746
rect 15764 2694 15776 2746
rect 15838 2694 15840 2746
rect 15678 2692 15702 2694
rect 15758 2692 15782 2694
rect 15838 2692 15862 2694
rect 15622 2672 15918 2692
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 14830 82 14886 480
rect 14568 54 14886 82
rect 15948 82 15976 3062
rect 17144 2650 17172 3431
rect 19289 3292 19585 3312
rect 19345 3290 19369 3292
rect 19425 3290 19449 3292
rect 19505 3290 19529 3292
rect 19367 3238 19369 3290
rect 19431 3238 19443 3290
rect 19505 3238 19507 3290
rect 19345 3236 19369 3238
rect 19425 3236 19449 3238
rect 19505 3236 19529 3238
rect 19289 3216 19585 3236
rect 18418 3088 18474 3097
rect 18418 3023 18474 3032
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 16118 82 16174 480
rect 15948 54 16174 82
rect 17144 82 17172 2314
rect 17406 82 17462 480
rect 17144 54 17462 82
rect 18432 82 18460 3023
rect 19289 2204 19585 2224
rect 19345 2202 19369 2204
rect 19425 2202 19449 2204
rect 19505 2202 19529 2204
rect 19367 2150 19369 2202
rect 19431 2150 19443 2202
rect 19505 2150 19507 2202
rect 19345 2148 19369 2150
rect 19425 2148 19449 2150
rect 19505 2148 19529 2150
rect 19289 2128 19585 2148
rect 19706 1592 19762 1601
rect 19706 1527 19762 1536
rect 18694 82 18750 480
rect 18432 54 18750 82
rect 19720 82 19748 1527
rect 19982 82 20038 480
rect 19720 54 20038 82
rect 21008 82 21036 3878
rect 21546 1320 21602 1329
rect 21546 1255 21602 1264
rect 21270 82 21326 480
rect 21560 105 21588 1255
rect 21008 54 21326 82
rect 12254 0 12310 54
rect 13542 0 13598 54
rect 14830 0 14886 54
rect 16118 0 16174 54
rect 17406 0 17462 54
rect 18694 0 18750 54
rect 19982 0 20038 54
rect 21270 0 21326 54
rect 21546 96 21602 105
rect 21546 31 21602 40
<< via2 >>
rect 1398 20304 1454 20360
rect 1306 15952 1362 16008
rect 1582 11872 1638 11928
rect 1398 10376 1454 10432
rect 4622 19610 4678 19612
rect 4702 19610 4758 19612
rect 4782 19610 4838 19612
rect 4862 19610 4918 19612
rect 4622 19558 4648 19610
rect 4648 19558 4678 19610
rect 4702 19558 4712 19610
rect 4712 19558 4758 19610
rect 4782 19558 4828 19610
rect 4828 19558 4838 19610
rect 4862 19558 4892 19610
rect 4892 19558 4918 19610
rect 4622 19556 4678 19558
rect 4702 19556 4758 19558
rect 4782 19556 4838 19558
rect 4862 19556 4918 19558
rect 110 7656 166 7712
rect 110 5480 166 5536
rect 110 4528 166 4584
rect 1582 3712 1638 3768
rect 1858 3884 1860 3904
rect 1860 3884 1912 3904
rect 1912 3884 1914 3904
rect 1858 3848 1914 3884
rect 4622 18522 4678 18524
rect 4702 18522 4758 18524
rect 4782 18522 4838 18524
rect 4862 18522 4918 18524
rect 4622 18470 4648 18522
rect 4648 18470 4678 18522
rect 4702 18470 4712 18522
rect 4712 18470 4758 18522
rect 4782 18470 4828 18522
rect 4828 18470 4838 18522
rect 4862 18470 4892 18522
rect 4892 18470 4918 18522
rect 4622 18468 4678 18470
rect 4702 18468 4758 18470
rect 4782 18468 4838 18470
rect 4862 18468 4918 18470
rect 8289 19066 8345 19068
rect 8369 19066 8425 19068
rect 8449 19066 8505 19068
rect 8529 19066 8585 19068
rect 8289 19014 8315 19066
rect 8315 19014 8345 19066
rect 8369 19014 8379 19066
rect 8379 19014 8425 19066
rect 8449 19014 8495 19066
rect 8495 19014 8505 19066
rect 8529 19014 8559 19066
rect 8559 19014 8585 19066
rect 8289 19012 8345 19014
rect 8369 19012 8425 19014
rect 8449 19012 8505 19014
rect 8529 19012 8585 19014
rect 4802 18128 4858 18184
rect 4622 17434 4678 17436
rect 4702 17434 4758 17436
rect 4782 17434 4838 17436
rect 4862 17434 4918 17436
rect 4622 17382 4648 17434
rect 4648 17382 4678 17434
rect 4702 17382 4712 17434
rect 4712 17382 4758 17434
rect 4782 17382 4828 17434
rect 4828 17382 4838 17434
rect 4862 17382 4892 17434
rect 4892 17382 4918 17434
rect 4622 17380 4678 17382
rect 4702 17380 4758 17382
rect 4782 17380 4838 17382
rect 4862 17380 4918 17382
rect 4622 16346 4678 16348
rect 4702 16346 4758 16348
rect 4782 16346 4838 16348
rect 4862 16346 4918 16348
rect 4622 16294 4648 16346
rect 4648 16294 4678 16346
rect 4702 16294 4712 16346
rect 4712 16294 4758 16346
rect 4782 16294 4828 16346
rect 4828 16294 4838 16346
rect 4862 16294 4892 16346
rect 4892 16294 4918 16346
rect 4622 16292 4678 16294
rect 4702 16292 4758 16294
rect 4782 16292 4838 16294
rect 4862 16292 4918 16294
rect 4622 15258 4678 15260
rect 4702 15258 4758 15260
rect 4782 15258 4838 15260
rect 4862 15258 4918 15260
rect 4622 15206 4648 15258
rect 4648 15206 4678 15258
rect 4702 15206 4712 15258
rect 4712 15206 4758 15258
rect 4782 15206 4828 15258
rect 4828 15206 4838 15258
rect 4862 15206 4892 15258
rect 4892 15206 4918 15258
rect 4622 15204 4678 15206
rect 4702 15204 4758 15206
rect 4782 15204 4838 15206
rect 4862 15204 4918 15206
rect 4622 14170 4678 14172
rect 4702 14170 4758 14172
rect 4782 14170 4838 14172
rect 4862 14170 4918 14172
rect 4622 14118 4648 14170
rect 4648 14118 4678 14170
rect 4702 14118 4712 14170
rect 4712 14118 4758 14170
rect 4782 14118 4828 14170
rect 4828 14118 4838 14170
rect 4862 14118 4892 14170
rect 4892 14118 4918 14170
rect 4622 14116 4678 14118
rect 4702 14116 4758 14118
rect 4782 14116 4838 14118
rect 4862 14116 4918 14118
rect 4622 13082 4678 13084
rect 4702 13082 4758 13084
rect 4782 13082 4838 13084
rect 4862 13082 4918 13084
rect 4622 13030 4648 13082
rect 4648 13030 4678 13082
rect 4702 13030 4712 13082
rect 4712 13030 4758 13082
rect 4782 13030 4828 13082
rect 4828 13030 4838 13082
rect 4862 13030 4892 13082
rect 4892 13030 4918 13082
rect 4622 13028 4678 13030
rect 4702 13028 4758 13030
rect 4782 13028 4838 13030
rect 4862 13028 4918 13030
rect 4622 11994 4678 11996
rect 4702 11994 4758 11996
rect 4782 11994 4838 11996
rect 4862 11994 4918 11996
rect 4622 11942 4648 11994
rect 4648 11942 4678 11994
rect 4702 11942 4712 11994
rect 4712 11942 4758 11994
rect 4782 11942 4828 11994
rect 4828 11942 4838 11994
rect 4862 11942 4892 11994
rect 4892 11942 4918 11994
rect 4622 11940 4678 11942
rect 4702 11940 4758 11942
rect 4782 11940 4838 11942
rect 4862 11940 4918 11942
rect 4622 10906 4678 10908
rect 4702 10906 4758 10908
rect 4782 10906 4838 10908
rect 4862 10906 4918 10908
rect 4622 10854 4648 10906
rect 4648 10854 4678 10906
rect 4702 10854 4712 10906
rect 4712 10854 4758 10906
rect 4782 10854 4828 10906
rect 4828 10854 4838 10906
rect 4862 10854 4892 10906
rect 4892 10854 4918 10906
rect 4622 10852 4678 10854
rect 4702 10852 4758 10854
rect 4782 10852 4838 10854
rect 4862 10852 4918 10854
rect 4622 9818 4678 9820
rect 4702 9818 4758 9820
rect 4782 9818 4838 9820
rect 4862 9818 4918 9820
rect 4622 9766 4648 9818
rect 4648 9766 4678 9818
rect 4702 9766 4712 9818
rect 4712 9766 4758 9818
rect 4782 9766 4828 9818
rect 4828 9766 4838 9818
rect 4862 9766 4892 9818
rect 4892 9766 4918 9818
rect 4622 9764 4678 9766
rect 4702 9764 4758 9766
rect 4782 9764 4838 9766
rect 4862 9764 4918 9766
rect 4622 8730 4678 8732
rect 4702 8730 4758 8732
rect 4782 8730 4838 8732
rect 4862 8730 4918 8732
rect 4622 8678 4648 8730
rect 4648 8678 4678 8730
rect 4702 8678 4712 8730
rect 4712 8678 4758 8730
rect 4782 8678 4828 8730
rect 4828 8678 4838 8730
rect 4862 8678 4892 8730
rect 4892 8678 4918 8730
rect 4622 8676 4678 8678
rect 4702 8676 4758 8678
rect 4782 8676 4838 8678
rect 4862 8676 4918 8678
rect 7562 13776 7618 13832
rect 5078 8880 5134 8936
rect 4622 7642 4678 7644
rect 4702 7642 4758 7644
rect 4782 7642 4838 7644
rect 4862 7642 4918 7644
rect 4622 7590 4648 7642
rect 4648 7590 4678 7642
rect 4702 7590 4712 7642
rect 4712 7590 4758 7642
rect 4782 7590 4828 7642
rect 4828 7590 4838 7642
rect 4862 7590 4892 7642
rect 4892 7590 4918 7642
rect 4622 7588 4678 7590
rect 4702 7588 4758 7590
rect 4782 7588 4838 7590
rect 4862 7588 4918 7590
rect 4622 6554 4678 6556
rect 4702 6554 4758 6556
rect 4782 6554 4838 6556
rect 4862 6554 4918 6556
rect 4622 6502 4648 6554
rect 4648 6502 4678 6554
rect 4702 6502 4712 6554
rect 4712 6502 4758 6554
rect 4782 6502 4828 6554
rect 4828 6502 4838 6554
rect 4862 6502 4892 6554
rect 4892 6502 4918 6554
rect 4622 6500 4678 6502
rect 4702 6500 4758 6502
rect 4782 6500 4838 6502
rect 4862 6500 4918 6502
rect 4802 5888 4858 5944
rect 4622 5466 4678 5468
rect 4702 5466 4758 5468
rect 4782 5466 4838 5468
rect 4862 5466 4918 5468
rect 4622 5414 4648 5466
rect 4648 5414 4678 5466
rect 4702 5414 4712 5466
rect 4712 5414 4758 5466
rect 4782 5414 4828 5466
rect 4828 5414 4838 5466
rect 4862 5414 4892 5466
rect 4892 5414 4918 5466
rect 4622 5412 4678 5414
rect 4702 5412 4758 5414
rect 4782 5412 4838 5414
rect 4862 5412 4918 5414
rect 2410 3576 2466 3632
rect 2686 3576 2742 3632
rect 2134 1672 2190 1728
rect 4622 4378 4678 4380
rect 4702 4378 4758 4380
rect 4782 4378 4838 4380
rect 4862 4378 4918 4380
rect 4622 4326 4648 4378
rect 4648 4326 4678 4378
rect 4702 4326 4712 4378
rect 4712 4326 4758 4378
rect 4782 4326 4828 4378
rect 4828 4326 4838 4378
rect 4862 4326 4892 4378
rect 4892 4326 4918 4378
rect 4622 4324 4678 4326
rect 4702 4324 4758 4326
rect 4782 4324 4838 4326
rect 4862 4324 4918 4326
rect 4526 3984 4582 4040
rect 4710 3848 4766 3904
rect 5446 4664 5502 4720
rect 4622 3290 4678 3292
rect 4702 3290 4758 3292
rect 4782 3290 4838 3292
rect 4862 3290 4918 3292
rect 4622 3238 4648 3290
rect 4648 3238 4678 3290
rect 4702 3238 4712 3290
rect 4712 3238 4758 3290
rect 4782 3238 4828 3290
rect 4828 3238 4838 3290
rect 4862 3238 4892 3290
rect 4892 3238 4918 3290
rect 4622 3236 4678 3238
rect 4702 3236 4758 3238
rect 4782 3236 4838 3238
rect 4862 3236 4918 3238
rect 4622 2202 4678 2204
rect 4702 2202 4758 2204
rect 4782 2202 4838 2204
rect 4862 2202 4918 2204
rect 4622 2150 4648 2202
rect 4648 2150 4678 2202
rect 4702 2150 4712 2202
rect 4712 2150 4758 2202
rect 4782 2150 4828 2202
rect 4828 2150 4838 2202
rect 4862 2150 4892 2202
rect 4892 2150 4918 2202
rect 4622 2148 4678 2150
rect 4702 2148 4758 2150
rect 4782 2148 4838 2150
rect 4862 2148 4918 2150
rect 6642 10648 6698 10704
rect 6274 5888 6330 5944
rect 8289 17978 8345 17980
rect 8369 17978 8425 17980
rect 8449 17978 8505 17980
rect 8529 17978 8585 17980
rect 8289 17926 8315 17978
rect 8315 17926 8345 17978
rect 8369 17926 8379 17978
rect 8379 17926 8425 17978
rect 8449 17926 8495 17978
rect 8495 17926 8505 17978
rect 8529 17926 8559 17978
rect 8559 17926 8585 17978
rect 8289 17924 8345 17926
rect 8369 17924 8425 17926
rect 8449 17924 8505 17926
rect 8529 17924 8585 17926
rect 8289 16890 8345 16892
rect 8369 16890 8425 16892
rect 8449 16890 8505 16892
rect 8529 16890 8585 16892
rect 8289 16838 8315 16890
rect 8315 16838 8345 16890
rect 8369 16838 8379 16890
rect 8379 16838 8425 16890
rect 8449 16838 8495 16890
rect 8495 16838 8505 16890
rect 8529 16838 8559 16890
rect 8559 16838 8585 16890
rect 8289 16836 8345 16838
rect 8369 16836 8425 16838
rect 8449 16836 8505 16838
rect 8529 16836 8585 16838
rect 8289 15802 8345 15804
rect 8369 15802 8425 15804
rect 8449 15802 8505 15804
rect 8529 15802 8585 15804
rect 8289 15750 8315 15802
rect 8315 15750 8345 15802
rect 8369 15750 8379 15802
rect 8379 15750 8425 15802
rect 8449 15750 8495 15802
rect 8495 15750 8505 15802
rect 8529 15750 8559 15802
rect 8559 15750 8585 15802
rect 8289 15748 8345 15750
rect 8369 15748 8425 15750
rect 8449 15748 8505 15750
rect 8529 15748 8585 15750
rect 8289 14714 8345 14716
rect 8369 14714 8425 14716
rect 8449 14714 8505 14716
rect 8529 14714 8585 14716
rect 8289 14662 8315 14714
rect 8315 14662 8345 14714
rect 8369 14662 8379 14714
rect 8379 14662 8425 14714
rect 8449 14662 8495 14714
rect 8495 14662 8505 14714
rect 8529 14662 8559 14714
rect 8559 14662 8585 14714
rect 8289 14660 8345 14662
rect 8369 14660 8425 14662
rect 8449 14660 8505 14662
rect 8529 14660 8585 14662
rect 8289 13626 8345 13628
rect 8369 13626 8425 13628
rect 8449 13626 8505 13628
rect 8529 13626 8585 13628
rect 8289 13574 8315 13626
rect 8315 13574 8345 13626
rect 8369 13574 8379 13626
rect 8379 13574 8425 13626
rect 8449 13574 8495 13626
rect 8495 13574 8505 13626
rect 8529 13574 8559 13626
rect 8559 13574 8585 13626
rect 8289 13572 8345 13574
rect 8369 13572 8425 13574
rect 8449 13572 8505 13574
rect 8529 13572 8585 13574
rect 8289 12538 8345 12540
rect 8369 12538 8425 12540
rect 8449 12538 8505 12540
rect 8529 12538 8585 12540
rect 8289 12486 8315 12538
rect 8315 12486 8345 12538
rect 8369 12486 8379 12538
rect 8379 12486 8425 12538
rect 8449 12486 8495 12538
rect 8495 12486 8505 12538
rect 8529 12486 8559 12538
rect 8559 12486 8585 12538
rect 8289 12484 8345 12486
rect 8369 12484 8425 12486
rect 8449 12484 8505 12486
rect 8529 12484 8585 12486
rect 8289 11450 8345 11452
rect 8369 11450 8425 11452
rect 8449 11450 8505 11452
rect 8529 11450 8585 11452
rect 8289 11398 8315 11450
rect 8315 11398 8345 11450
rect 8369 11398 8379 11450
rect 8379 11398 8425 11450
rect 8449 11398 8495 11450
rect 8495 11398 8505 11450
rect 8529 11398 8559 11450
rect 8559 11398 8585 11450
rect 8289 11396 8345 11398
rect 8369 11396 8425 11398
rect 8449 11396 8505 11398
rect 8529 11396 8585 11398
rect 11956 19610 12012 19612
rect 12036 19610 12092 19612
rect 12116 19610 12172 19612
rect 12196 19610 12252 19612
rect 11956 19558 11982 19610
rect 11982 19558 12012 19610
rect 12036 19558 12046 19610
rect 12046 19558 12092 19610
rect 12116 19558 12162 19610
rect 12162 19558 12172 19610
rect 12196 19558 12226 19610
rect 12226 19558 12252 19610
rect 11956 19556 12012 19558
rect 12036 19556 12092 19558
rect 12116 19556 12172 19558
rect 12196 19556 12252 19558
rect 11956 18522 12012 18524
rect 12036 18522 12092 18524
rect 12116 18522 12172 18524
rect 12196 18522 12252 18524
rect 11956 18470 11982 18522
rect 11982 18470 12012 18522
rect 12036 18470 12046 18522
rect 12046 18470 12092 18522
rect 12116 18470 12162 18522
rect 12162 18470 12172 18522
rect 12196 18470 12226 18522
rect 12226 18470 12252 18522
rect 11956 18468 12012 18470
rect 12036 18468 12092 18470
rect 12116 18468 12172 18470
rect 12196 18468 12252 18470
rect 8289 10362 8345 10364
rect 8369 10362 8425 10364
rect 8449 10362 8505 10364
rect 8529 10362 8585 10364
rect 8289 10310 8315 10362
rect 8315 10310 8345 10362
rect 8369 10310 8379 10362
rect 8379 10310 8425 10362
rect 8449 10310 8495 10362
rect 8495 10310 8505 10362
rect 8529 10310 8559 10362
rect 8559 10310 8585 10362
rect 8289 10308 8345 10310
rect 8369 10308 8425 10310
rect 8449 10308 8505 10310
rect 8529 10308 8585 10310
rect 8289 9274 8345 9276
rect 8369 9274 8425 9276
rect 8449 9274 8505 9276
rect 8529 9274 8585 9276
rect 8289 9222 8315 9274
rect 8315 9222 8345 9274
rect 8369 9222 8379 9274
rect 8379 9222 8425 9274
rect 8449 9222 8495 9274
rect 8495 9222 8505 9274
rect 8529 9222 8559 9274
rect 8559 9222 8585 9274
rect 8289 9220 8345 9222
rect 8369 9220 8425 9222
rect 8449 9220 8505 9222
rect 8529 9220 8585 9222
rect 8289 8186 8345 8188
rect 8369 8186 8425 8188
rect 8449 8186 8505 8188
rect 8529 8186 8585 8188
rect 8289 8134 8315 8186
rect 8315 8134 8345 8186
rect 8369 8134 8379 8186
rect 8379 8134 8425 8186
rect 8449 8134 8495 8186
rect 8495 8134 8505 8186
rect 8529 8134 8559 8186
rect 8559 8134 8585 8186
rect 8289 8132 8345 8134
rect 8369 8132 8425 8134
rect 8449 8132 8505 8134
rect 8529 8132 8585 8134
rect 5630 3440 5686 3496
rect 6918 2352 6974 2408
rect 8289 7098 8345 7100
rect 8369 7098 8425 7100
rect 8449 7098 8505 7100
rect 8529 7098 8585 7100
rect 8289 7046 8315 7098
rect 8315 7046 8345 7098
rect 8369 7046 8379 7098
rect 8379 7046 8425 7098
rect 8449 7046 8495 7098
rect 8495 7046 8505 7098
rect 8529 7046 8559 7098
rect 8559 7046 8585 7098
rect 8289 7044 8345 7046
rect 8369 7044 8425 7046
rect 8449 7044 8505 7046
rect 8529 7044 8585 7046
rect 8289 6010 8345 6012
rect 8369 6010 8425 6012
rect 8449 6010 8505 6012
rect 8529 6010 8585 6012
rect 8289 5958 8315 6010
rect 8315 5958 8345 6010
rect 8369 5958 8379 6010
rect 8379 5958 8425 6010
rect 8449 5958 8495 6010
rect 8495 5958 8505 6010
rect 8529 5958 8559 6010
rect 8559 5958 8585 6010
rect 8289 5956 8345 5958
rect 8369 5956 8425 5958
rect 8449 5956 8505 5958
rect 8529 5956 8585 5958
rect 7838 3576 7894 3632
rect 8289 4922 8345 4924
rect 8369 4922 8425 4924
rect 8449 4922 8505 4924
rect 8529 4922 8585 4924
rect 8289 4870 8315 4922
rect 8315 4870 8345 4922
rect 8369 4870 8379 4922
rect 8379 4870 8425 4922
rect 8449 4870 8495 4922
rect 8495 4870 8505 4922
rect 8529 4870 8559 4922
rect 8559 4870 8585 4922
rect 8289 4868 8345 4870
rect 8369 4868 8425 4870
rect 8449 4868 8505 4870
rect 8529 4868 8585 4870
rect 8574 4528 8630 4584
rect 8666 3984 8722 4040
rect 8289 3834 8345 3836
rect 8369 3834 8425 3836
rect 8449 3834 8505 3836
rect 8529 3834 8585 3836
rect 8289 3782 8315 3834
rect 8315 3782 8345 3834
rect 8369 3782 8379 3834
rect 8379 3782 8425 3834
rect 8449 3782 8495 3834
rect 8495 3782 8505 3834
rect 8529 3782 8559 3834
rect 8559 3782 8585 3834
rect 8289 3780 8345 3782
rect 8369 3780 8425 3782
rect 8449 3780 8505 3782
rect 8529 3780 8585 3782
rect 9770 6160 9826 6216
rect 8850 3576 8906 3632
rect 8942 3304 8998 3360
rect 11242 3984 11298 4040
rect 8289 2746 8345 2748
rect 8369 2746 8425 2748
rect 8449 2746 8505 2748
rect 8529 2746 8585 2748
rect 8289 2694 8315 2746
rect 8315 2694 8345 2746
rect 8369 2694 8379 2746
rect 8379 2694 8425 2746
rect 8449 2694 8495 2746
rect 8495 2694 8505 2746
rect 8529 2694 8559 2746
rect 8559 2694 8585 2746
rect 8289 2692 8345 2694
rect 8369 2692 8425 2694
rect 8449 2692 8505 2694
rect 8529 2692 8585 2694
rect 11956 17434 12012 17436
rect 12036 17434 12092 17436
rect 12116 17434 12172 17436
rect 12196 17434 12252 17436
rect 11956 17382 11982 17434
rect 11982 17382 12012 17434
rect 12036 17382 12046 17434
rect 12046 17382 12092 17434
rect 12116 17382 12162 17434
rect 12162 17382 12172 17434
rect 12196 17382 12226 17434
rect 12226 17382 12252 17434
rect 11956 17380 12012 17382
rect 12036 17380 12092 17382
rect 12116 17380 12172 17382
rect 12196 17380 12252 17382
rect 11956 16346 12012 16348
rect 12036 16346 12092 16348
rect 12116 16346 12172 16348
rect 12196 16346 12252 16348
rect 11956 16294 11982 16346
rect 11982 16294 12012 16346
rect 12036 16294 12046 16346
rect 12046 16294 12092 16346
rect 12116 16294 12162 16346
rect 12162 16294 12172 16346
rect 12196 16294 12226 16346
rect 12226 16294 12252 16346
rect 11956 16292 12012 16294
rect 12036 16292 12092 16294
rect 12116 16292 12172 16294
rect 12196 16292 12252 16294
rect 11956 15258 12012 15260
rect 12036 15258 12092 15260
rect 12116 15258 12172 15260
rect 12196 15258 12252 15260
rect 11956 15206 11982 15258
rect 11982 15206 12012 15258
rect 12036 15206 12046 15258
rect 12046 15206 12092 15258
rect 12116 15206 12162 15258
rect 12162 15206 12172 15258
rect 12196 15206 12226 15258
rect 12226 15206 12252 15258
rect 11956 15204 12012 15206
rect 12036 15204 12092 15206
rect 12116 15204 12172 15206
rect 12196 15204 12252 15206
rect 11956 14170 12012 14172
rect 12036 14170 12092 14172
rect 12116 14170 12172 14172
rect 12196 14170 12252 14172
rect 11956 14118 11982 14170
rect 11982 14118 12012 14170
rect 12036 14118 12046 14170
rect 12046 14118 12092 14170
rect 12116 14118 12162 14170
rect 12162 14118 12172 14170
rect 12196 14118 12226 14170
rect 12226 14118 12252 14170
rect 11956 14116 12012 14118
rect 12036 14116 12092 14118
rect 12116 14116 12172 14118
rect 12196 14116 12252 14118
rect 11956 13082 12012 13084
rect 12036 13082 12092 13084
rect 12116 13082 12172 13084
rect 12196 13082 12252 13084
rect 11956 13030 11982 13082
rect 11982 13030 12012 13082
rect 12036 13030 12046 13082
rect 12046 13030 12092 13082
rect 12116 13030 12162 13082
rect 12162 13030 12172 13082
rect 12196 13030 12226 13082
rect 12226 13030 12252 13082
rect 11956 13028 12012 13030
rect 12036 13028 12092 13030
rect 12116 13028 12172 13030
rect 12196 13028 12252 13030
rect 11956 11994 12012 11996
rect 12036 11994 12092 11996
rect 12116 11994 12172 11996
rect 12196 11994 12252 11996
rect 11956 11942 11982 11994
rect 11982 11942 12012 11994
rect 12036 11942 12046 11994
rect 12046 11942 12092 11994
rect 12116 11942 12162 11994
rect 12162 11942 12172 11994
rect 12196 11942 12226 11994
rect 12226 11942 12252 11994
rect 11956 11940 12012 11942
rect 12036 11940 12092 11942
rect 12116 11940 12172 11942
rect 12196 11940 12252 11942
rect 11956 10906 12012 10908
rect 12036 10906 12092 10908
rect 12116 10906 12172 10908
rect 12196 10906 12252 10908
rect 11956 10854 11982 10906
rect 11982 10854 12012 10906
rect 12036 10854 12046 10906
rect 12046 10854 12092 10906
rect 12116 10854 12162 10906
rect 12162 10854 12172 10906
rect 12196 10854 12226 10906
rect 12226 10854 12252 10906
rect 11956 10852 12012 10854
rect 12036 10852 12092 10854
rect 12116 10852 12172 10854
rect 12196 10852 12252 10854
rect 12622 11192 12678 11248
rect 12530 10512 12586 10568
rect 15622 19066 15678 19068
rect 15702 19066 15758 19068
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15622 19014 15648 19066
rect 15648 19014 15678 19066
rect 15702 19014 15712 19066
rect 15712 19014 15758 19066
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15918 19066
rect 15622 19012 15678 19014
rect 15702 19012 15758 19014
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 15622 17978 15678 17980
rect 15702 17978 15758 17980
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15622 17926 15648 17978
rect 15648 17926 15678 17978
rect 15702 17926 15712 17978
rect 15712 17926 15758 17978
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15918 17978
rect 15622 17924 15678 17926
rect 15702 17924 15758 17926
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 15622 16890 15678 16892
rect 15702 16890 15758 16892
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15622 16838 15648 16890
rect 15648 16838 15678 16890
rect 15702 16838 15712 16890
rect 15712 16838 15758 16890
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15918 16890
rect 15622 16836 15678 16838
rect 15702 16836 15758 16838
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15622 15802 15678 15804
rect 15702 15802 15758 15804
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15622 15750 15648 15802
rect 15648 15750 15678 15802
rect 15702 15750 15712 15802
rect 15712 15750 15758 15802
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15918 15802
rect 15622 15748 15678 15750
rect 15702 15748 15758 15750
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15622 14714 15678 14716
rect 15702 14714 15758 14716
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15622 14662 15648 14714
rect 15648 14662 15678 14714
rect 15702 14662 15712 14714
rect 15712 14662 15758 14714
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15918 14714
rect 15622 14660 15678 14662
rect 15702 14660 15758 14662
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15622 13626 15678 13628
rect 15702 13626 15758 13628
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15622 13574 15648 13626
rect 15648 13574 15678 13626
rect 15702 13574 15712 13626
rect 15712 13574 15758 13626
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15918 13626
rect 15622 13572 15678 13574
rect 15702 13572 15758 13574
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15622 12538 15678 12540
rect 15702 12538 15758 12540
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15622 12486 15648 12538
rect 15648 12486 15678 12538
rect 15702 12486 15712 12538
rect 15712 12486 15758 12538
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15918 12538
rect 15622 12484 15678 12486
rect 15702 12484 15758 12486
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15622 11450 15678 11452
rect 15702 11450 15758 11452
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15622 11398 15648 11450
rect 15648 11398 15678 11450
rect 15702 11398 15712 11450
rect 15712 11398 15758 11450
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15918 11450
rect 15622 11396 15678 11398
rect 15702 11396 15758 11398
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15382 10648 15438 10704
rect 15622 10362 15678 10364
rect 15702 10362 15758 10364
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15622 10310 15648 10362
rect 15648 10310 15678 10362
rect 15702 10310 15712 10362
rect 15712 10310 15758 10362
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15918 10362
rect 15622 10308 15678 10310
rect 15702 10308 15758 10310
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 11956 9818 12012 9820
rect 12036 9818 12092 9820
rect 12116 9818 12172 9820
rect 12196 9818 12252 9820
rect 11956 9766 11982 9818
rect 11982 9766 12012 9818
rect 12036 9766 12046 9818
rect 12046 9766 12092 9818
rect 12116 9766 12162 9818
rect 12162 9766 12172 9818
rect 12196 9766 12226 9818
rect 12226 9766 12252 9818
rect 11956 9764 12012 9766
rect 12036 9764 12092 9766
rect 12116 9764 12172 9766
rect 12196 9764 12252 9766
rect 11956 8730 12012 8732
rect 12036 8730 12092 8732
rect 12116 8730 12172 8732
rect 12196 8730 12252 8732
rect 11956 8678 11982 8730
rect 11982 8678 12012 8730
rect 12036 8678 12046 8730
rect 12046 8678 12092 8730
rect 12116 8678 12162 8730
rect 12162 8678 12172 8730
rect 12196 8678 12226 8730
rect 12226 8678 12252 8730
rect 11956 8676 12012 8678
rect 12036 8676 12092 8678
rect 12116 8676 12172 8678
rect 12196 8676 12252 8678
rect 11956 7642 12012 7644
rect 12036 7642 12092 7644
rect 12116 7642 12172 7644
rect 12196 7642 12252 7644
rect 11956 7590 11982 7642
rect 11982 7590 12012 7642
rect 12036 7590 12046 7642
rect 12046 7590 12092 7642
rect 12116 7590 12162 7642
rect 12162 7590 12172 7642
rect 12196 7590 12226 7642
rect 12226 7590 12252 7642
rect 11956 7588 12012 7590
rect 12036 7588 12092 7590
rect 12116 7588 12172 7590
rect 12196 7588 12252 7590
rect 11956 6554 12012 6556
rect 12036 6554 12092 6556
rect 12116 6554 12172 6556
rect 12196 6554 12252 6556
rect 11956 6502 11982 6554
rect 11982 6502 12012 6554
rect 12036 6502 12046 6554
rect 12046 6502 12092 6554
rect 12116 6502 12162 6554
rect 12162 6502 12172 6554
rect 12196 6502 12226 6554
rect 12226 6502 12252 6554
rect 11956 6500 12012 6502
rect 12036 6500 12092 6502
rect 12116 6500 12172 6502
rect 12196 6500 12252 6502
rect 12714 9560 12770 9616
rect 12622 8336 12678 8392
rect 11956 5466 12012 5468
rect 12036 5466 12092 5468
rect 12116 5466 12172 5468
rect 12196 5466 12252 5468
rect 11956 5414 11982 5466
rect 11982 5414 12012 5466
rect 12036 5414 12046 5466
rect 12046 5414 12092 5466
rect 12116 5414 12162 5466
rect 12162 5414 12172 5466
rect 12196 5414 12226 5466
rect 12226 5414 12252 5466
rect 11956 5412 12012 5414
rect 12036 5412 12092 5414
rect 12116 5412 12172 5414
rect 12196 5412 12252 5414
rect 11886 5072 11942 5128
rect 11956 4378 12012 4380
rect 12036 4378 12092 4380
rect 12116 4378 12172 4380
rect 12196 4378 12252 4380
rect 11956 4326 11982 4378
rect 11982 4326 12012 4378
rect 12036 4326 12046 4378
rect 12046 4326 12092 4378
rect 12116 4326 12162 4378
rect 12162 4326 12172 4378
rect 12196 4326 12226 4378
rect 12226 4326 12252 4378
rect 11956 4324 12012 4326
rect 12036 4324 12092 4326
rect 12116 4324 12172 4326
rect 12196 4324 12252 4326
rect 12990 3440 13046 3496
rect 11794 3304 11850 3360
rect 11956 3290 12012 3292
rect 12036 3290 12092 3292
rect 12116 3290 12172 3292
rect 12196 3290 12252 3292
rect 11956 3238 11982 3290
rect 11982 3238 12012 3290
rect 12036 3238 12046 3290
rect 12046 3238 12092 3290
rect 12116 3238 12162 3290
rect 12162 3238 12172 3290
rect 12196 3238 12226 3290
rect 12226 3238 12252 3290
rect 11956 3236 12012 3238
rect 12036 3236 12092 3238
rect 12116 3236 12172 3238
rect 12196 3236 12252 3238
rect 12254 2352 12310 2408
rect 11956 2202 12012 2204
rect 12036 2202 12092 2204
rect 12116 2202 12172 2204
rect 12196 2202 12252 2204
rect 11956 2150 11982 2202
rect 11982 2150 12012 2202
rect 12036 2150 12046 2202
rect 12046 2150 12092 2202
rect 12116 2150 12162 2202
rect 12162 2150 12172 2202
rect 12196 2150 12226 2202
rect 12226 2150 12252 2202
rect 11956 2148 12012 2150
rect 12036 2148 12092 2150
rect 12116 2148 12172 2150
rect 12196 2148 12252 2150
rect 11518 40 11574 96
rect 15622 9274 15678 9276
rect 15702 9274 15758 9276
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15622 9222 15648 9274
rect 15648 9222 15678 9274
rect 15702 9222 15712 9274
rect 15712 9222 15758 9274
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15918 9274
rect 15622 9220 15678 9222
rect 15702 9220 15758 9222
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15622 8186 15678 8188
rect 15702 8186 15758 8188
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15622 8134 15648 8186
rect 15648 8134 15678 8186
rect 15702 8134 15712 8186
rect 15712 8134 15758 8186
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15918 8186
rect 15622 8132 15678 8134
rect 15702 8132 15758 8134
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15622 7098 15678 7100
rect 15702 7098 15758 7100
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15622 7046 15648 7098
rect 15648 7046 15678 7098
rect 15702 7046 15712 7098
rect 15712 7046 15758 7098
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15918 7098
rect 15622 7044 15678 7046
rect 15702 7044 15758 7046
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 17222 20304 17278 20360
rect 19289 19610 19345 19612
rect 19369 19610 19425 19612
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19289 19558 19315 19610
rect 19315 19558 19345 19610
rect 19369 19558 19379 19610
rect 19379 19558 19425 19610
rect 19449 19558 19495 19610
rect 19495 19558 19505 19610
rect 19529 19558 19559 19610
rect 19559 19558 19585 19610
rect 19289 19556 19345 19558
rect 19369 19556 19425 19558
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19289 18522 19345 18524
rect 19369 18522 19425 18524
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19289 18470 19315 18522
rect 19315 18470 19345 18522
rect 19369 18470 19379 18522
rect 19379 18470 19425 18522
rect 19449 18470 19495 18522
rect 19495 18470 19505 18522
rect 19529 18470 19559 18522
rect 19559 18470 19585 18522
rect 19289 18468 19345 18470
rect 19369 18468 19425 18470
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19289 17434 19345 17436
rect 19369 17434 19425 17436
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19289 17382 19315 17434
rect 19315 17382 19345 17434
rect 19369 17382 19379 17434
rect 19379 17382 19425 17434
rect 19449 17382 19495 17434
rect 19495 17382 19505 17434
rect 19529 17382 19559 17434
rect 19559 17382 19585 17434
rect 19289 17380 19345 17382
rect 19369 17380 19425 17382
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19289 16346 19345 16348
rect 19369 16346 19425 16348
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19289 16294 19315 16346
rect 19315 16294 19345 16346
rect 19369 16294 19379 16346
rect 19379 16294 19425 16346
rect 19449 16294 19495 16346
rect 19495 16294 19505 16346
rect 19529 16294 19559 16346
rect 19559 16294 19585 16346
rect 19289 16292 19345 16294
rect 19369 16292 19425 16294
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19062 15408 19118 15464
rect 19289 15258 19345 15260
rect 19369 15258 19425 15260
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19289 15206 19315 15258
rect 19315 15206 19345 15258
rect 19369 15206 19379 15258
rect 19379 15206 19425 15258
rect 19449 15206 19495 15258
rect 19495 15206 19505 15258
rect 19529 15206 19559 15258
rect 19559 15206 19585 15258
rect 19289 15204 19345 15206
rect 19369 15204 19425 15206
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19289 14170 19345 14172
rect 19369 14170 19425 14172
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19289 14118 19315 14170
rect 19315 14118 19345 14170
rect 19369 14118 19379 14170
rect 19379 14118 19425 14170
rect 19449 14118 19495 14170
rect 19495 14118 19505 14170
rect 19529 14118 19559 14170
rect 19559 14118 19585 14170
rect 19289 14116 19345 14118
rect 19369 14116 19425 14118
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19154 13640 19210 13696
rect 19289 13082 19345 13084
rect 19369 13082 19425 13084
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19289 13030 19315 13082
rect 19315 13030 19345 13082
rect 19369 13030 19379 13082
rect 19379 13030 19425 13082
rect 19449 13030 19495 13082
rect 19495 13030 19505 13082
rect 19529 13030 19559 13082
rect 19559 13030 19585 13082
rect 19289 13028 19345 13030
rect 19369 13028 19425 13030
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19289 11994 19345 11996
rect 19369 11994 19425 11996
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19289 11942 19315 11994
rect 19315 11942 19345 11994
rect 19369 11942 19379 11994
rect 19379 11942 19425 11994
rect 19449 11942 19495 11994
rect 19495 11942 19505 11994
rect 19529 11942 19559 11994
rect 19559 11942 19585 11994
rect 19289 11940 19345 11942
rect 19369 11940 19425 11942
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19289 10906 19345 10908
rect 19369 10906 19425 10908
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19289 10854 19315 10906
rect 19315 10854 19345 10906
rect 19369 10854 19379 10906
rect 19379 10854 19425 10906
rect 19449 10854 19495 10906
rect 19495 10854 19505 10906
rect 19529 10854 19559 10906
rect 19559 10854 19585 10906
rect 19289 10852 19345 10854
rect 19369 10852 19425 10854
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19289 9818 19345 9820
rect 19369 9818 19425 9820
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19289 9766 19315 9818
rect 19315 9766 19345 9818
rect 19369 9766 19379 9818
rect 19379 9766 19425 9818
rect 19449 9766 19495 9818
rect 19495 9766 19505 9818
rect 19529 9766 19559 9818
rect 19559 9766 19585 9818
rect 19289 9764 19345 9766
rect 19369 9764 19425 9766
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19890 17856 19946 17912
rect 19706 10512 19762 10568
rect 19614 9560 19670 9616
rect 19289 8730 19345 8732
rect 19369 8730 19425 8732
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19289 8678 19315 8730
rect 19315 8678 19345 8730
rect 19369 8678 19379 8730
rect 19379 8678 19425 8730
rect 19449 8678 19495 8730
rect 19495 8678 19505 8730
rect 19529 8678 19559 8730
rect 19559 8678 19585 8730
rect 19289 8676 19345 8678
rect 19369 8676 19425 8678
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19289 7642 19345 7644
rect 19369 7642 19425 7644
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19289 7590 19315 7642
rect 19315 7590 19345 7642
rect 19369 7590 19379 7642
rect 19379 7590 19425 7642
rect 19449 7590 19495 7642
rect 19495 7590 19505 7642
rect 19529 7590 19559 7642
rect 19559 7590 19585 7642
rect 19289 7588 19345 7590
rect 19369 7588 19425 7590
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19289 6554 19345 6556
rect 19369 6554 19425 6556
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19289 6502 19315 6554
rect 19315 6502 19345 6554
rect 19369 6502 19379 6554
rect 19379 6502 19425 6554
rect 19449 6502 19495 6554
rect 19495 6502 19505 6554
rect 19529 6502 19559 6554
rect 19559 6502 19585 6554
rect 19289 6500 19345 6502
rect 19369 6500 19425 6502
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 16578 6160 16634 6216
rect 15622 6010 15678 6012
rect 15702 6010 15758 6012
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15622 5958 15648 6010
rect 15648 5958 15678 6010
rect 15702 5958 15712 6010
rect 15712 5958 15758 6010
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15918 6010
rect 15622 5956 15678 5958
rect 15702 5956 15758 5958
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 13726 5616 13782 5672
rect 15382 5616 15438 5672
rect 19289 5466 19345 5468
rect 19369 5466 19425 5468
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19289 5414 19315 5466
rect 19315 5414 19345 5466
rect 19369 5414 19379 5466
rect 19379 5414 19425 5466
rect 19449 5414 19495 5466
rect 19495 5414 19505 5466
rect 19529 5414 19559 5466
rect 19559 5414 19585 5466
rect 19289 5412 19345 5414
rect 19369 5412 19425 5414
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 13542 5072 13598 5128
rect 15622 4922 15678 4924
rect 15702 4922 15758 4924
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15622 4870 15648 4922
rect 15648 4870 15678 4922
rect 15702 4870 15712 4922
rect 15712 4870 15758 4922
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15918 4922
rect 15622 4868 15678 4870
rect 15702 4868 15758 4870
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 13450 4684 13506 4720
rect 13450 4664 13452 4684
rect 13452 4664 13504 4684
rect 13504 4664 13506 4684
rect 13634 4528 13690 4584
rect 19289 4378 19345 4380
rect 19369 4378 19425 4380
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19289 4326 19315 4378
rect 19315 4326 19345 4378
rect 19369 4326 19379 4378
rect 19379 4326 19425 4378
rect 19449 4326 19495 4378
rect 19495 4326 19505 4378
rect 19529 4326 19559 4378
rect 19559 4326 19585 4378
rect 19289 4324 19345 4326
rect 19369 4324 19425 4326
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 15622 3834 15678 3836
rect 15702 3834 15758 3836
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15622 3782 15648 3834
rect 15648 3782 15678 3834
rect 15702 3782 15712 3834
rect 15712 3782 15758 3834
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15918 3834
rect 15622 3780 15678 3782
rect 15702 3780 15758 3782
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 17130 3440 17186 3496
rect 15622 2746 15678 2748
rect 15702 2746 15758 2748
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15622 2694 15648 2746
rect 15648 2694 15678 2746
rect 15702 2694 15712 2746
rect 15712 2694 15758 2746
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15918 2746
rect 15622 2692 15678 2694
rect 15702 2692 15758 2694
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 19289 3290 19345 3292
rect 19369 3290 19425 3292
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19289 3238 19315 3290
rect 19315 3238 19345 3290
rect 19369 3238 19379 3290
rect 19379 3238 19425 3290
rect 19449 3238 19495 3290
rect 19495 3238 19505 3290
rect 19529 3238 19559 3290
rect 19559 3238 19585 3290
rect 19289 3236 19345 3238
rect 19369 3236 19425 3238
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 18418 3032 18474 3088
rect 19289 2202 19345 2204
rect 19369 2202 19425 2204
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19289 2150 19315 2202
rect 19315 2150 19345 2202
rect 19369 2150 19379 2202
rect 19379 2150 19425 2202
rect 19449 2150 19495 2202
rect 19495 2150 19505 2202
rect 19529 2150 19559 2202
rect 19559 2150 19585 2202
rect 19289 2148 19345 2150
rect 19369 2148 19425 2150
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 19706 1536 19762 1592
rect 21546 1264 21602 1320
rect 21546 40 21602 96
<< metal3 >>
rect 0 20816 480 20936
rect 21520 20816 22000 20936
rect 62 20362 122 20816
rect 1393 20362 1459 20365
rect 62 20360 1459 20362
rect 62 20304 1398 20360
rect 1454 20304 1459 20360
rect 62 20302 1459 20304
rect 1393 20299 1459 20302
rect 17217 20362 17283 20365
rect 21590 20362 21650 20816
rect 17217 20360 21650 20362
rect 17217 20304 17222 20360
rect 17278 20304 21650 20360
rect 17217 20302 21650 20304
rect 17217 20299 17283 20302
rect 4610 19616 4930 19617
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4930 19616
rect 4610 19551 4930 19552
rect 11944 19616 12264 19617
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 19551 12264 19552
rect 19277 19616 19597 19617
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 19551 19597 19552
rect 8277 19072 8597 19073
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 19007 8597 19008
rect 15610 19072 15930 19073
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 19007 15930 19008
rect 0 18640 480 18760
rect 62 18186 122 18640
rect 4610 18528 4930 18529
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4930 18528
rect 4610 18463 4930 18464
rect 11944 18528 12264 18529
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 18463 12264 18464
rect 19277 18528 19597 18529
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 18463 19597 18464
rect 21520 18368 22000 18488
rect 4797 18186 4863 18189
rect 62 18184 4863 18186
rect 62 18128 4802 18184
rect 4858 18128 4863 18184
rect 62 18126 4863 18128
rect 4797 18123 4863 18126
rect 8277 17984 8597 17985
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 17919 8597 17920
rect 15610 17984 15930 17985
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 17919 15930 17920
rect 19885 17914 19951 17917
rect 21590 17914 21650 18368
rect 19885 17912 21650 17914
rect 19885 17856 19890 17912
rect 19946 17856 21650 17912
rect 19885 17854 21650 17856
rect 19885 17851 19951 17854
rect 4610 17440 4930 17441
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4930 17440
rect 4610 17375 4930 17376
rect 11944 17440 12264 17441
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 17375 12264 17376
rect 19277 17440 19597 17441
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 17375 19597 17376
rect 8277 16896 8597 16897
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 16831 8597 16832
rect 15610 16896 15930 16897
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 16831 15930 16832
rect 0 16464 480 16584
rect 62 16010 122 16464
rect 4610 16352 4930 16353
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4930 16352
rect 4610 16287 4930 16288
rect 11944 16352 12264 16353
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 16287 12264 16288
rect 19277 16352 19597 16353
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 16287 19597 16288
rect 1301 16010 1367 16013
rect 62 16008 1367 16010
rect 62 15952 1306 16008
rect 1362 15952 1367 16008
rect 62 15950 1367 15952
rect 1301 15947 1367 15950
rect 21520 15920 22000 16040
rect 8277 15808 8597 15809
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 15743 8597 15744
rect 15610 15808 15930 15809
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 15743 15930 15744
rect 19057 15466 19123 15469
rect 21590 15466 21650 15920
rect 19057 15464 21650 15466
rect 19057 15408 19062 15464
rect 19118 15408 21650 15464
rect 19057 15406 21650 15408
rect 19057 15403 19123 15406
rect 4610 15264 4930 15265
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4930 15264
rect 4610 15199 4930 15200
rect 11944 15264 12264 15265
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 15199 12264 15200
rect 19277 15264 19597 15265
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 15199 19597 15200
rect 8277 14720 8597 14721
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 14655 8597 14656
rect 15610 14720 15930 14721
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 14655 15930 14656
rect 0 14288 480 14408
rect 62 13834 122 14288
rect 4610 14176 4930 14177
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4930 14176
rect 4610 14111 4930 14112
rect 11944 14176 12264 14177
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 14111 12264 14112
rect 19277 14176 19597 14177
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 14111 19597 14112
rect 7557 13834 7623 13837
rect 21582 13834 21588 13836
rect 62 13832 7623 13834
rect 62 13776 7562 13832
rect 7618 13776 7623 13832
rect 62 13774 7623 13776
rect 7557 13771 7623 13774
rect 19290 13774 21588 13834
rect 19149 13698 19215 13701
rect 19290 13698 19350 13774
rect 21582 13772 21588 13774
rect 21652 13772 21658 13836
rect 19149 13696 19350 13698
rect 19149 13640 19154 13696
rect 19210 13640 19350 13696
rect 19149 13638 19350 13640
rect 19149 13635 19215 13638
rect 8277 13632 8597 13633
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 13567 8597 13568
rect 15610 13632 15930 13633
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 13567 15930 13568
rect 21520 13564 22000 13592
rect 21520 13562 21588 13564
rect 21460 13502 21588 13562
rect 21520 13500 21588 13502
rect 21652 13500 22000 13564
rect 21520 13472 22000 13500
rect 4610 13088 4930 13089
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4930 13088
rect 4610 13023 4930 13024
rect 11944 13088 12264 13089
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 13023 12264 13024
rect 19277 13088 19597 13089
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 13023 19597 13024
rect 8277 12544 8597 12545
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 12479 8597 12480
rect 15610 12544 15930 12545
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 12479 15930 12480
rect 0 12112 480 12232
rect 62 11930 122 12112
rect 4610 12000 4930 12001
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4930 12000
rect 4610 11935 4930 11936
rect 11944 12000 12264 12001
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 11935 12264 11936
rect 19277 12000 19597 12001
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 11935 19597 11936
rect 1577 11930 1643 11933
rect 62 11928 1643 11930
rect 62 11872 1582 11928
rect 1638 11872 1643 11928
rect 62 11870 1643 11872
rect 1577 11867 1643 11870
rect 8277 11456 8597 11457
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 11391 8597 11392
rect 15610 11456 15930 11457
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 11391 15930 11392
rect 12617 11250 12683 11253
rect 21398 11250 21404 11252
rect 12617 11248 21404 11250
rect 12617 11192 12622 11248
rect 12678 11192 21404 11248
rect 12617 11190 21404 11192
rect 12617 11187 12683 11190
rect 21398 11188 21404 11190
rect 21468 11188 21474 11252
rect 21520 11116 22000 11144
rect 21520 11114 21588 11116
rect 21460 11054 21588 11114
rect 21520 11052 21588 11054
rect 21652 11052 22000 11116
rect 21520 11024 22000 11052
rect 4610 10912 4930 10913
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4930 10912
rect 4610 10847 4930 10848
rect 11944 10912 12264 10913
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 10847 12264 10848
rect 19277 10912 19597 10913
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 10847 19597 10848
rect 6637 10706 6703 10709
rect 15377 10706 15443 10709
rect 6637 10704 15443 10706
rect 6637 10648 6642 10704
rect 6698 10648 15382 10704
rect 15438 10648 15443 10704
rect 6637 10646 15443 10648
rect 6637 10643 6703 10646
rect 15377 10643 15443 10646
rect 12525 10570 12591 10573
rect 19701 10570 19767 10573
rect 12525 10568 19767 10570
rect 12525 10512 12530 10568
rect 12586 10512 19706 10568
rect 19762 10512 19767 10568
rect 12525 10510 19767 10512
rect 12525 10507 12591 10510
rect 19701 10507 19767 10510
rect 1393 10434 1459 10437
rect 62 10432 1459 10434
rect 62 10376 1398 10432
rect 1454 10376 1459 10432
rect 62 10374 1459 10376
rect 62 9920 122 10374
rect 1393 10371 1459 10374
rect 8277 10368 8597 10369
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 10303 8597 10304
rect 15610 10368 15930 10369
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 10303 15930 10304
rect 0 9800 480 9920
rect 4610 9824 4930 9825
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4930 9824
rect 4610 9759 4930 9760
rect 11944 9824 12264 9825
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 9759 12264 9760
rect 19277 9824 19597 9825
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 9759 19597 9760
rect 12709 9618 12775 9621
rect 19609 9618 19675 9621
rect 12709 9616 19675 9618
rect 12709 9560 12714 9616
rect 12770 9560 19614 9616
rect 19670 9560 19675 9616
rect 12709 9558 19675 9560
rect 12709 9555 12775 9558
rect 19609 9555 19675 9558
rect 8277 9280 8597 9281
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 8277 9215 8597 9216
rect 15610 9280 15930 9281
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 9215 15930 9216
rect 5073 8938 5139 8941
rect 5206 8938 5212 8940
rect 5073 8936 5212 8938
rect 5073 8880 5078 8936
rect 5134 8880 5212 8936
rect 5073 8878 5212 8880
rect 5073 8875 5139 8878
rect 5206 8876 5212 8878
rect 5276 8876 5282 8940
rect 4610 8736 4930 8737
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4930 8736
rect 4610 8671 4930 8672
rect 11944 8736 12264 8737
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 8671 12264 8672
rect 19277 8736 19597 8737
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 8671 19597 8672
rect 21520 8576 22000 8696
rect 12617 8394 12683 8397
rect 21590 8394 21650 8576
rect 12617 8392 21650 8394
rect 12617 8336 12622 8392
rect 12678 8336 21650 8392
rect 12617 8334 21650 8336
rect 12617 8331 12683 8334
rect 8277 8192 8597 8193
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 8127 8597 8128
rect 15610 8192 15930 8193
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 8127 15930 8128
rect 0 7712 480 7744
rect 0 7656 110 7712
rect 166 7656 480 7712
rect 0 7624 480 7656
rect 4610 7648 4930 7649
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4930 7648
rect 4610 7583 4930 7584
rect 11944 7648 12264 7649
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 7583 12264 7584
rect 19277 7648 19597 7649
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 7583 19597 7584
rect 8277 7104 8597 7105
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 7039 8597 7040
rect 15610 7104 15930 7105
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 7039 15930 7040
rect 4610 6560 4930 6561
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4930 6560
rect 4610 6495 4930 6496
rect 11944 6560 12264 6561
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 6495 12264 6496
rect 19277 6560 19597 6561
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 6495 19597 6496
rect 9765 6218 9831 6221
rect 16573 6218 16639 6221
rect 9765 6216 16639 6218
rect 9765 6160 9770 6216
rect 9826 6160 16578 6216
rect 16634 6160 16639 6216
rect 9765 6158 16639 6160
rect 9765 6155 9831 6158
rect 16573 6155 16639 6158
rect 21520 6128 22000 6248
rect 8277 6016 8597 6017
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 5951 8597 5952
rect 15610 6016 15930 6017
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 5951 15930 5952
rect 4797 5946 4863 5949
rect 6269 5946 6335 5949
rect 4797 5944 6335 5946
rect 4797 5888 4802 5944
rect 4858 5888 6274 5944
rect 6330 5888 6335 5944
rect 4797 5886 6335 5888
rect 4797 5883 4863 5886
rect 6269 5883 6335 5886
rect 13721 5674 13787 5677
rect 15377 5674 15443 5677
rect 21590 5674 21650 6128
rect 13721 5672 21650 5674
rect 13721 5616 13726 5672
rect 13782 5616 15382 5672
rect 15438 5616 21650 5672
rect 13721 5614 21650 5616
rect 13721 5611 13787 5614
rect 15377 5611 15443 5614
rect 0 5536 480 5568
rect 0 5480 110 5536
rect 166 5480 480 5536
rect 0 5448 480 5480
rect 4610 5472 4930 5473
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4930 5472
rect 4610 5407 4930 5408
rect 11944 5472 12264 5473
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 5407 12264 5408
rect 19277 5472 19597 5473
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 5407 19597 5408
rect 11881 5130 11947 5133
rect 13537 5130 13603 5133
rect 4110 5128 13603 5130
rect 4110 5072 11886 5128
rect 11942 5072 13542 5128
rect 13598 5072 13603 5128
rect 4110 5070 13603 5072
rect 105 4586 171 4589
rect 4110 4586 4170 5070
rect 11881 5067 11947 5070
rect 13537 5067 13603 5070
rect 8277 4928 8597 4929
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 4863 8597 4864
rect 15610 4928 15930 4929
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 4863 15930 4864
rect 5441 4722 5507 4725
rect 13445 4722 13511 4725
rect 5441 4720 13511 4722
rect 5441 4664 5446 4720
rect 5502 4664 13450 4720
rect 13506 4664 13511 4720
rect 5441 4662 13511 4664
rect 5441 4659 5507 4662
rect 13445 4659 13511 4662
rect 105 4584 4170 4586
rect 105 4528 110 4584
rect 166 4528 4170 4584
rect 105 4526 4170 4528
rect 8569 4586 8635 4589
rect 13629 4586 13695 4589
rect 8569 4584 13695 4586
rect 8569 4528 8574 4584
rect 8630 4528 13634 4584
rect 13690 4528 13695 4584
rect 8569 4526 13695 4528
rect 105 4523 171 4526
rect 8569 4523 8635 4526
rect 13629 4523 13695 4526
rect 4610 4384 4930 4385
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4930 4384
rect 4610 4319 4930 4320
rect 11944 4384 12264 4385
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 4319 12264 4320
rect 19277 4384 19597 4385
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 4319 19597 4320
rect 4521 4042 4587 4045
rect 8661 4042 8727 4045
rect 11237 4042 11303 4045
rect 4521 4040 11303 4042
rect 4521 3984 4526 4040
rect 4582 3984 8666 4040
rect 8722 3984 11242 4040
rect 11298 3984 11303 4040
rect 4521 3982 11303 3984
rect 4521 3979 4587 3982
rect 8661 3979 8727 3982
rect 11237 3979 11303 3982
rect 1853 3906 1919 3909
rect 62 3904 1919 3906
rect 62 3848 1858 3904
rect 1914 3848 1919 3904
rect 62 3846 1919 3848
rect 62 3392 122 3846
rect 1853 3843 1919 3846
rect 4705 3906 4771 3909
rect 4705 3904 8034 3906
rect 4705 3848 4710 3904
rect 4766 3848 8034 3904
rect 4705 3846 8034 3848
rect 4705 3843 4771 3846
rect 1577 3770 1643 3773
rect 4102 3770 4108 3772
rect 1577 3768 4108 3770
rect 1577 3712 1582 3768
rect 1638 3712 4108 3768
rect 1577 3710 4108 3712
rect 1577 3707 1643 3710
rect 4102 3708 4108 3710
rect 4172 3708 4178 3772
rect 2405 3634 2471 3637
rect 2681 3634 2747 3637
rect 7833 3634 7899 3637
rect 2405 3632 7899 3634
rect 2405 3576 2410 3632
rect 2466 3576 2686 3632
rect 2742 3576 7838 3632
rect 7894 3576 7899 3632
rect 2405 3574 7899 3576
rect 7974 3634 8034 3846
rect 8277 3840 8597 3841
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 3775 8597 3776
rect 15610 3840 15930 3841
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 3775 15930 3776
rect 21520 3680 22000 3800
rect 8845 3634 8911 3637
rect 7974 3632 8911 3634
rect 7974 3576 8850 3632
rect 8906 3576 8911 3632
rect 7974 3574 8911 3576
rect 2405 3571 2471 3574
rect 2681 3571 2747 3574
rect 7833 3571 7899 3574
rect 8845 3571 8911 3574
rect 5625 3498 5691 3501
rect 12985 3498 13051 3501
rect 5625 3496 13051 3498
rect 5625 3440 5630 3496
rect 5686 3440 12990 3496
rect 13046 3440 13051 3496
rect 5625 3438 13051 3440
rect 5625 3435 5691 3438
rect 12985 3435 13051 3438
rect 17125 3498 17191 3501
rect 21590 3498 21650 3680
rect 17125 3496 21650 3498
rect 17125 3440 17130 3496
rect 17186 3440 21650 3496
rect 17125 3438 21650 3440
rect 17125 3435 17191 3438
rect 0 3272 480 3392
rect 8937 3362 9003 3365
rect 11789 3362 11855 3365
rect 8937 3360 11855 3362
rect 8937 3304 8942 3360
rect 8998 3304 11794 3360
rect 11850 3304 11855 3360
rect 8937 3302 11855 3304
rect 8937 3299 9003 3302
rect 11789 3299 11855 3302
rect 4610 3296 4930 3297
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4930 3296
rect 4610 3231 4930 3232
rect 11944 3296 12264 3297
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 3231 12264 3232
rect 19277 3296 19597 3297
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 19277 3231 19597 3232
rect 18270 3028 18276 3092
rect 18340 3090 18346 3092
rect 18413 3090 18479 3093
rect 18340 3088 18479 3090
rect 18340 3032 18418 3088
rect 18474 3032 18479 3088
rect 18340 3030 18479 3032
rect 18340 3028 18346 3030
rect 18413 3027 18479 3030
rect 8277 2752 8597 2753
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2687 8597 2688
rect 15610 2752 15930 2753
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2687 15930 2688
rect 6913 2410 6979 2413
rect 12249 2410 12315 2413
rect 6913 2408 12315 2410
rect 6913 2352 6918 2408
rect 6974 2352 12254 2408
rect 12310 2352 12315 2408
rect 6913 2350 12315 2352
rect 6913 2347 6979 2350
rect 12249 2347 12315 2350
rect 4610 2208 4930 2209
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4930 2208
rect 4610 2143 4930 2144
rect 11944 2208 12264 2209
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2143 12264 2144
rect 19277 2208 19597 2209
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2143 19597 2144
rect 2129 1730 2195 1733
rect 62 1728 2195 1730
rect 62 1672 2134 1728
rect 2190 1672 2195 1728
rect 62 1670 2195 1672
rect 62 1216 122 1670
rect 2129 1667 2195 1670
rect 5206 1532 5212 1596
rect 5276 1594 5282 1596
rect 19701 1594 19767 1597
rect 5276 1592 19767 1594
rect 5276 1536 19706 1592
rect 19762 1536 19767 1592
rect 5276 1534 19767 1536
rect 5276 1532 5282 1534
rect 19701 1531 19767 1534
rect 21520 1322 22000 1352
rect 21460 1320 22000 1322
rect 21460 1264 21546 1320
rect 21602 1264 22000 1320
rect 21460 1262 22000 1264
rect 21520 1232 22000 1262
rect 0 1096 480 1216
rect 11513 98 11579 101
rect 21541 98 21607 101
rect 11513 96 21607 98
rect 11513 40 11518 96
rect 11574 40 21546 96
rect 21602 40 21607 96
rect 11513 38 21607 40
rect 11513 35 11579 38
rect 21541 35 21607 38
<< via3 >>
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 4698 19612 4762 19616
rect 4698 19556 4702 19612
rect 4702 19556 4758 19612
rect 4758 19556 4762 19612
rect 4698 19552 4762 19556
rect 4778 19612 4842 19616
rect 4778 19556 4782 19612
rect 4782 19556 4838 19612
rect 4838 19556 4842 19612
rect 4778 19552 4842 19556
rect 4858 19612 4922 19616
rect 4858 19556 4862 19612
rect 4862 19556 4918 19612
rect 4918 19556 4922 19612
rect 4858 19552 4922 19556
rect 11952 19612 12016 19616
rect 11952 19556 11956 19612
rect 11956 19556 12012 19612
rect 12012 19556 12016 19612
rect 11952 19552 12016 19556
rect 12032 19612 12096 19616
rect 12032 19556 12036 19612
rect 12036 19556 12092 19612
rect 12092 19556 12096 19612
rect 12032 19552 12096 19556
rect 12112 19612 12176 19616
rect 12112 19556 12116 19612
rect 12116 19556 12172 19612
rect 12172 19556 12176 19612
rect 12112 19552 12176 19556
rect 12192 19612 12256 19616
rect 12192 19556 12196 19612
rect 12196 19556 12252 19612
rect 12252 19556 12256 19612
rect 12192 19552 12256 19556
rect 19285 19612 19349 19616
rect 19285 19556 19289 19612
rect 19289 19556 19345 19612
rect 19345 19556 19349 19612
rect 19285 19552 19349 19556
rect 19365 19612 19429 19616
rect 19365 19556 19369 19612
rect 19369 19556 19425 19612
rect 19425 19556 19429 19612
rect 19365 19552 19429 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 8285 19068 8349 19072
rect 8285 19012 8289 19068
rect 8289 19012 8345 19068
rect 8345 19012 8349 19068
rect 8285 19008 8349 19012
rect 8365 19068 8429 19072
rect 8365 19012 8369 19068
rect 8369 19012 8425 19068
rect 8425 19012 8429 19068
rect 8365 19008 8429 19012
rect 8445 19068 8509 19072
rect 8445 19012 8449 19068
rect 8449 19012 8505 19068
rect 8505 19012 8509 19068
rect 8445 19008 8509 19012
rect 8525 19068 8589 19072
rect 8525 19012 8529 19068
rect 8529 19012 8585 19068
rect 8585 19012 8589 19068
rect 8525 19008 8589 19012
rect 15618 19068 15682 19072
rect 15618 19012 15622 19068
rect 15622 19012 15678 19068
rect 15678 19012 15682 19068
rect 15618 19008 15682 19012
rect 15698 19068 15762 19072
rect 15698 19012 15702 19068
rect 15702 19012 15758 19068
rect 15758 19012 15762 19068
rect 15698 19008 15762 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 4698 18524 4762 18528
rect 4698 18468 4702 18524
rect 4702 18468 4758 18524
rect 4758 18468 4762 18524
rect 4698 18464 4762 18468
rect 4778 18524 4842 18528
rect 4778 18468 4782 18524
rect 4782 18468 4838 18524
rect 4838 18468 4842 18524
rect 4778 18464 4842 18468
rect 4858 18524 4922 18528
rect 4858 18468 4862 18524
rect 4862 18468 4918 18524
rect 4918 18468 4922 18524
rect 4858 18464 4922 18468
rect 11952 18524 12016 18528
rect 11952 18468 11956 18524
rect 11956 18468 12012 18524
rect 12012 18468 12016 18524
rect 11952 18464 12016 18468
rect 12032 18524 12096 18528
rect 12032 18468 12036 18524
rect 12036 18468 12092 18524
rect 12092 18468 12096 18524
rect 12032 18464 12096 18468
rect 12112 18524 12176 18528
rect 12112 18468 12116 18524
rect 12116 18468 12172 18524
rect 12172 18468 12176 18524
rect 12112 18464 12176 18468
rect 12192 18524 12256 18528
rect 12192 18468 12196 18524
rect 12196 18468 12252 18524
rect 12252 18468 12256 18524
rect 12192 18464 12256 18468
rect 19285 18524 19349 18528
rect 19285 18468 19289 18524
rect 19289 18468 19345 18524
rect 19345 18468 19349 18524
rect 19285 18464 19349 18468
rect 19365 18524 19429 18528
rect 19365 18468 19369 18524
rect 19369 18468 19425 18524
rect 19425 18468 19429 18524
rect 19365 18464 19429 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 8285 17980 8349 17984
rect 8285 17924 8289 17980
rect 8289 17924 8345 17980
rect 8345 17924 8349 17980
rect 8285 17920 8349 17924
rect 8365 17980 8429 17984
rect 8365 17924 8369 17980
rect 8369 17924 8425 17980
rect 8425 17924 8429 17980
rect 8365 17920 8429 17924
rect 8445 17980 8509 17984
rect 8445 17924 8449 17980
rect 8449 17924 8505 17980
rect 8505 17924 8509 17980
rect 8445 17920 8509 17924
rect 8525 17980 8589 17984
rect 8525 17924 8529 17980
rect 8529 17924 8585 17980
rect 8585 17924 8589 17980
rect 8525 17920 8589 17924
rect 15618 17980 15682 17984
rect 15618 17924 15622 17980
rect 15622 17924 15678 17980
rect 15678 17924 15682 17980
rect 15618 17920 15682 17924
rect 15698 17980 15762 17984
rect 15698 17924 15702 17980
rect 15702 17924 15758 17980
rect 15758 17924 15762 17980
rect 15698 17920 15762 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 4698 17436 4762 17440
rect 4698 17380 4702 17436
rect 4702 17380 4758 17436
rect 4758 17380 4762 17436
rect 4698 17376 4762 17380
rect 4778 17436 4842 17440
rect 4778 17380 4782 17436
rect 4782 17380 4838 17436
rect 4838 17380 4842 17436
rect 4778 17376 4842 17380
rect 4858 17436 4922 17440
rect 4858 17380 4862 17436
rect 4862 17380 4918 17436
rect 4918 17380 4922 17436
rect 4858 17376 4922 17380
rect 11952 17436 12016 17440
rect 11952 17380 11956 17436
rect 11956 17380 12012 17436
rect 12012 17380 12016 17436
rect 11952 17376 12016 17380
rect 12032 17436 12096 17440
rect 12032 17380 12036 17436
rect 12036 17380 12092 17436
rect 12092 17380 12096 17436
rect 12032 17376 12096 17380
rect 12112 17436 12176 17440
rect 12112 17380 12116 17436
rect 12116 17380 12172 17436
rect 12172 17380 12176 17436
rect 12112 17376 12176 17380
rect 12192 17436 12256 17440
rect 12192 17380 12196 17436
rect 12196 17380 12252 17436
rect 12252 17380 12256 17436
rect 12192 17376 12256 17380
rect 19285 17436 19349 17440
rect 19285 17380 19289 17436
rect 19289 17380 19345 17436
rect 19345 17380 19349 17436
rect 19285 17376 19349 17380
rect 19365 17436 19429 17440
rect 19365 17380 19369 17436
rect 19369 17380 19425 17436
rect 19425 17380 19429 17436
rect 19365 17376 19429 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 8285 16892 8349 16896
rect 8285 16836 8289 16892
rect 8289 16836 8345 16892
rect 8345 16836 8349 16892
rect 8285 16832 8349 16836
rect 8365 16892 8429 16896
rect 8365 16836 8369 16892
rect 8369 16836 8425 16892
rect 8425 16836 8429 16892
rect 8365 16832 8429 16836
rect 8445 16892 8509 16896
rect 8445 16836 8449 16892
rect 8449 16836 8505 16892
rect 8505 16836 8509 16892
rect 8445 16832 8509 16836
rect 8525 16892 8589 16896
rect 8525 16836 8529 16892
rect 8529 16836 8585 16892
rect 8585 16836 8589 16892
rect 8525 16832 8589 16836
rect 15618 16892 15682 16896
rect 15618 16836 15622 16892
rect 15622 16836 15678 16892
rect 15678 16836 15682 16892
rect 15618 16832 15682 16836
rect 15698 16892 15762 16896
rect 15698 16836 15702 16892
rect 15702 16836 15758 16892
rect 15758 16836 15762 16892
rect 15698 16832 15762 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 4698 16348 4762 16352
rect 4698 16292 4702 16348
rect 4702 16292 4758 16348
rect 4758 16292 4762 16348
rect 4698 16288 4762 16292
rect 4778 16348 4842 16352
rect 4778 16292 4782 16348
rect 4782 16292 4838 16348
rect 4838 16292 4842 16348
rect 4778 16288 4842 16292
rect 4858 16348 4922 16352
rect 4858 16292 4862 16348
rect 4862 16292 4918 16348
rect 4918 16292 4922 16348
rect 4858 16288 4922 16292
rect 11952 16348 12016 16352
rect 11952 16292 11956 16348
rect 11956 16292 12012 16348
rect 12012 16292 12016 16348
rect 11952 16288 12016 16292
rect 12032 16348 12096 16352
rect 12032 16292 12036 16348
rect 12036 16292 12092 16348
rect 12092 16292 12096 16348
rect 12032 16288 12096 16292
rect 12112 16348 12176 16352
rect 12112 16292 12116 16348
rect 12116 16292 12172 16348
rect 12172 16292 12176 16348
rect 12112 16288 12176 16292
rect 12192 16348 12256 16352
rect 12192 16292 12196 16348
rect 12196 16292 12252 16348
rect 12252 16292 12256 16348
rect 12192 16288 12256 16292
rect 19285 16348 19349 16352
rect 19285 16292 19289 16348
rect 19289 16292 19345 16348
rect 19345 16292 19349 16348
rect 19285 16288 19349 16292
rect 19365 16348 19429 16352
rect 19365 16292 19369 16348
rect 19369 16292 19425 16348
rect 19425 16292 19429 16348
rect 19365 16288 19429 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 8285 15804 8349 15808
rect 8285 15748 8289 15804
rect 8289 15748 8345 15804
rect 8345 15748 8349 15804
rect 8285 15744 8349 15748
rect 8365 15804 8429 15808
rect 8365 15748 8369 15804
rect 8369 15748 8425 15804
rect 8425 15748 8429 15804
rect 8365 15744 8429 15748
rect 8445 15804 8509 15808
rect 8445 15748 8449 15804
rect 8449 15748 8505 15804
rect 8505 15748 8509 15804
rect 8445 15744 8509 15748
rect 8525 15804 8589 15808
rect 8525 15748 8529 15804
rect 8529 15748 8585 15804
rect 8585 15748 8589 15804
rect 8525 15744 8589 15748
rect 15618 15804 15682 15808
rect 15618 15748 15622 15804
rect 15622 15748 15678 15804
rect 15678 15748 15682 15804
rect 15618 15744 15682 15748
rect 15698 15804 15762 15808
rect 15698 15748 15702 15804
rect 15702 15748 15758 15804
rect 15758 15748 15762 15804
rect 15698 15744 15762 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 4698 15260 4762 15264
rect 4698 15204 4702 15260
rect 4702 15204 4758 15260
rect 4758 15204 4762 15260
rect 4698 15200 4762 15204
rect 4778 15260 4842 15264
rect 4778 15204 4782 15260
rect 4782 15204 4838 15260
rect 4838 15204 4842 15260
rect 4778 15200 4842 15204
rect 4858 15260 4922 15264
rect 4858 15204 4862 15260
rect 4862 15204 4918 15260
rect 4918 15204 4922 15260
rect 4858 15200 4922 15204
rect 11952 15260 12016 15264
rect 11952 15204 11956 15260
rect 11956 15204 12012 15260
rect 12012 15204 12016 15260
rect 11952 15200 12016 15204
rect 12032 15260 12096 15264
rect 12032 15204 12036 15260
rect 12036 15204 12092 15260
rect 12092 15204 12096 15260
rect 12032 15200 12096 15204
rect 12112 15260 12176 15264
rect 12112 15204 12116 15260
rect 12116 15204 12172 15260
rect 12172 15204 12176 15260
rect 12112 15200 12176 15204
rect 12192 15260 12256 15264
rect 12192 15204 12196 15260
rect 12196 15204 12252 15260
rect 12252 15204 12256 15260
rect 12192 15200 12256 15204
rect 19285 15260 19349 15264
rect 19285 15204 19289 15260
rect 19289 15204 19345 15260
rect 19345 15204 19349 15260
rect 19285 15200 19349 15204
rect 19365 15260 19429 15264
rect 19365 15204 19369 15260
rect 19369 15204 19425 15260
rect 19425 15204 19429 15260
rect 19365 15200 19429 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 8285 14716 8349 14720
rect 8285 14660 8289 14716
rect 8289 14660 8345 14716
rect 8345 14660 8349 14716
rect 8285 14656 8349 14660
rect 8365 14716 8429 14720
rect 8365 14660 8369 14716
rect 8369 14660 8425 14716
rect 8425 14660 8429 14716
rect 8365 14656 8429 14660
rect 8445 14716 8509 14720
rect 8445 14660 8449 14716
rect 8449 14660 8505 14716
rect 8505 14660 8509 14716
rect 8445 14656 8509 14660
rect 8525 14716 8589 14720
rect 8525 14660 8529 14716
rect 8529 14660 8585 14716
rect 8585 14660 8589 14716
rect 8525 14656 8589 14660
rect 15618 14716 15682 14720
rect 15618 14660 15622 14716
rect 15622 14660 15678 14716
rect 15678 14660 15682 14716
rect 15618 14656 15682 14660
rect 15698 14716 15762 14720
rect 15698 14660 15702 14716
rect 15702 14660 15758 14716
rect 15758 14660 15762 14716
rect 15698 14656 15762 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 4698 14172 4762 14176
rect 4698 14116 4702 14172
rect 4702 14116 4758 14172
rect 4758 14116 4762 14172
rect 4698 14112 4762 14116
rect 4778 14172 4842 14176
rect 4778 14116 4782 14172
rect 4782 14116 4838 14172
rect 4838 14116 4842 14172
rect 4778 14112 4842 14116
rect 4858 14172 4922 14176
rect 4858 14116 4862 14172
rect 4862 14116 4918 14172
rect 4918 14116 4922 14172
rect 4858 14112 4922 14116
rect 11952 14172 12016 14176
rect 11952 14116 11956 14172
rect 11956 14116 12012 14172
rect 12012 14116 12016 14172
rect 11952 14112 12016 14116
rect 12032 14172 12096 14176
rect 12032 14116 12036 14172
rect 12036 14116 12092 14172
rect 12092 14116 12096 14172
rect 12032 14112 12096 14116
rect 12112 14172 12176 14176
rect 12112 14116 12116 14172
rect 12116 14116 12172 14172
rect 12172 14116 12176 14172
rect 12112 14112 12176 14116
rect 12192 14172 12256 14176
rect 12192 14116 12196 14172
rect 12196 14116 12252 14172
rect 12252 14116 12256 14172
rect 12192 14112 12256 14116
rect 19285 14172 19349 14176
rect 19285 14116 19289 14172
rect 19289 14116 19345 14172
rect 19345 14116 19349 14172
rect 19285 14112 19349 14116
rect 19365 14172 19429 14176
rect 19365 14116 19369 14172
rect 19369 14116 19425 14172
rect 19425 14116 19429 14172
rect 19365 14112 19429 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 21588 13772 21652 13836
rect 8285 13628 8349 13632
rect 8285 13572 8289 13628
rect 8289 13572 8345 13628
rect 8345 13572 8349 13628
rect 8285 13568 8349 13572
rect 8365 13628 8429 13632
rect 8365 13572 8369 13628
rect 8369 13572 8425 13628
rect 8425 13572 8429 13628
rect 8365 13568 8429 13572
rect 8445 13628 8509 13632
rect 8445 13572 8449 13628
rect 8449 13572 8505 13628
rect 8505 13572 8509 13628
rect 8445 13568 8509 13572
rect 8525 13628 8589 13632
rect 8525 13572 8529 13628
rect 8529 13572 8585 13628
rect 8585 13572 8589 13628
rect 8525 13568 8589 13572
rect 15618 13628 15682 13632
rect 15618 13572 15622 13628
rect 15622 13572 15678 13628
rect 15678 13572 15682 13628
rect 15618 13568 15682 13572
rect 15698 13628 15762 13632
rect 15698 13572 15702 13628
rect 15702 13572 15758 13628
rect 15758 13572 15762 13628
rect 15698 13568 15762 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 21588 13500 21652 13564
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 4698 13084 4762 13088
rect 4698 13028 4702 13084
rect 4702 13028 4758 13084
rect 4758 13028 4762 13084
rect 4698 13024 4762 13028
rect 4778 13084 4842 13088
rect 4778 13028 4782 13084
rect 4782 13028 4838 13084
rect 4838 13028 4842 13084
rect 4778 13024 4842 13028
rect 4858 13084 4922 13088
rect 4858 13028 4862 13084
rect 4862 13028 4918 13084
rect 4918 13028 4922 13084
rect 4858 13024 4922 13028
rect 11952 13084 12016 13088
rect 11952 13028 11956 13084
rect 11956 13028 12012 13084
rect 12012 13028 12016 13084
rect 11952 13024 12016 13028
rect 12032 13084 12096 13088
rect 12032 13028 12036 13084
rect 12036 13028 12092 13084
rect 12092 13028 12096 13084
rect 12032 13024 12096 13028
rect 12112 13084 12176 13088
rect 12112 13028 12116 13084
rect 12116 13028 12172 13084
rect 12172 13028 12176 13084
rect 12112 13024 12176 13028
rect 12192 13084 12256 13088
rect 12192 13028 12196 13084
rect 12196 13028 12252 13084
rect 12252 13028 12256 13084
rect 12192 13024 12256 13028
rect 19285 13084 19349 13088
rect 19285 13028 19289 13084
rect 19289 13028 19345 13084
rect 19345 13028 19349 13084
rect 19285 13024 19349 13028
rect 19365 13084 19429 13088
rect 19365 13028 19369 13084
rect 19369 13028 19425 13084
rect 19425 13028 19429 13084
rect 19365 13024 19429 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 8285 12540 8349 12544
rect 8285 12484 8289 12540
rect 8289 12484 8345 12540
rect 8345 12484 8349 12540
rect 8285 12480 8349 12484
rect 8365 12540 8429 12544
rect 8365 12484 8369 12540
rect 8369 12484 8425 12540
rect 8425 12484 8429 12540
rect 8365 12480 8429 12484
rect 8445 12540 8509 12544
rect 8445 12484 8449 12540
rect 8449 12484 8505 12540
rect 8505 12484 8509 12540
rect 8445 12480 8509 12484
rect 8525 12540 8589 12544
rect 8525 12484 8529 12540
rect 8529 12484 8585 12540
rect 8585 12484 8589 12540
rect 8525 12480 8589 12484
rect 15618 12540 15682 12544
rect 15618 12484 15622 12540
rect 15622 12484 15678 12540
rect 15678 12484 15682 12540
rect 15618 12480 15682 12484
rect 15698 12540 15762 12544
rect 15698 12484 15702 12540
rect 15702 12484 15758 12540
rect 15758 12484 15762 12540
rect 15698 12480 15762 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 4698 11996 4762 12000
rect 4698 11940 4702 11996
rect 4702 11940 4758 11996
rect 4758 11940 4762 11996
rect 4698 11936 4762 11940
rect 4778 11996 4842 12000
rect 4778 11940 4782 11996
rect 4782 11940 4838 11996
rect 4838 11940 4842 11996
rect 4778 11936 4842 11940
rect 4858 11996 4922 12000
rect 4858 11940 4862 11996
rect 4862 11940 4918 11996
rect 4918 11940 4922 11996
rect 4858 11936 4922 11940
rect 11952 11996 12016 12000
rect 11952 11940 11956 11996
rect 11956 11940 12012 11996
rect 12012 11940 12016 11996
rect 11952 11936 12016 11940
rect 12032 11996 12096 12000
rect 12032 11940 12036 11996
rect 12036 11940 12092 11996
rect 12092 11940 12096 11996
rect 12032 11936 12096 11940
rect 12112 11996 12176 12000
rect 12112 11940 12116 11996
rect 12116 11940 12172 11996
rect 12172 11940 12176 11996
rect 12112 11936 12176 11940
rect 12192 11996 12256 12000
rect 12192 11940 12196 11996
rect 12196 11940 12252 11996
rect 12252 11940 12256 11996
rect 12192 11936 12256 11940
rect 19285 11996 19349 12000
rect 19285 11940 19289 11996
rect 19289 11940 19345 11996
rect 19345 11940 19349 11996
rect 19285 11936 19349 11940
rect 19365 11996 19429 12000
rect 19365 11940 19369 11996
rect 19369 11940 19425 11996
rect 19425 11940 19429 11996
rect 19365 11936 19429 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 8285 11452 8349 11456
rect 8285 11396 8289 11452
rect 8289 11396 8345 11452
rect 8345 11396 8349 11452
rect 8285 11392 8349 11396
rect 8365 11452 8429 11456
rect 8365 11396 8369 11452
rect 8369 11396 8425 11452
rect 8425 11396 8429 11452
rect 8365 11392 8429 11396
rect 8445 11452 8509 11456
rect 8445 11396 8449 11452
rect 8449 11396 8505 11452
rect 8505 11396 8509 11452
rect 8445 11392 8509 11396
rect 8525 11452 8589 11456
rect 8525 11396 8529 11452
rect 8529 11396 8585 11452
rect 8585 11396 8589 11452
rect 8525 11392 8589 11396
rect 15618 11452 15682 11456
rect 15618 11396 15622 11452
rect 15622 11396 15678 11452
rect 15678 11396 15682 11452
rect 15618 11392 15682 11396
rect 15698 11452 15762 11456
rect 15698 11396 15702 11452
rect 15702 11396 15758 11452
rect 15758 11396 15762 11452
rect 15698 11392 15762 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 21404 11188 21468 11252
rect 21588 11052 21652 11116
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 4698 10908 4762 10912
rect 4698 10852 4702 10908
rect 4702 10852 4758 10908
rect 4758 10852 4762 10908
rect 4698 10848 4762 10852
rect 4778 10908 4842 10912
rect 4778 10852 4782 10908
rect 4782 10852 4838 10908
rect 4838 10852 4842 10908
rect 4778 10848 4842 10852
rect 4858 10908 4922 10912
rect 4858 10852 4862 10908
rect 4862 10852 4918 10908
rect 4918 10852 4922 10908
rect 4858 10848 4922 10852
rect 11952 10908 12016 10912
rect 11952 10852 11956 10908
rect 11956 10852 12012 10908
rect 12012 10852 12016 10908
rect 11952 10848 12016 10852
rect 12032 10908 12096 10912
rect 12032 10852 12036 10908
rect 12036 10852 12092 10908
rect 12092 10852 12096 10908
rect 12032 10848 12096 10852
rect 12112 10908 12176 10912
rect 12112 10852 12116 10908
rect 12116 10852 12172 10908
rect 12172 10852 12176 10908
rect 12112 10848 12176 10852
rect 12192 10908 12256 10912
rect 12192 10852 12196 10908
rect 12196 10852 12252 10908
rect 12252 10852 12256 10908
rect 12192 10848 12256 10852
rect 19285 10908 19349 10912
rect 19285 10852 19289 10908
rect 19289 10852 19345 10908
rect 19345 10852 19349 10908
rect 19285 10848 19349 10852
rect 19365 10908 19429 10912
rect 19365 10852 19369 10908
rect 19369 10852 19425 10908
rect 19425 10852 19429 10908
rect 19365 10848 19429 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 8285 10364 8349 10368
rect 8285 10308 8289 10364
rect 8289 10308 8345 10364
rect 8345 10308 8349 10364
rect 8285 10304 8349 10308
rect 8365 10364 8429 10368
rect 8365 10308 8369 10364
rect 8369 10308 8425 10364
rect 8425 10308 8429 10364
rect 8365 10304 8429 10308
rect 8445 10364 8509 10368
rect 8445 10308 8449 10364
rect 8449 10308 8505 10364
rect 8505 10308 8509 10364
rect 8445 10304 8509 10308
rect 8525 10364 8589 10368
rect 8525 10308 8529 10364
rect 8529 10308 8585 10364
rect 8585 10308 8589 10364
rect 8525 10304 8589 10308
rect 15618 10364 15682 10368
rect 15618 10308 15622 10364
rect 15622 10308 15678 10364
rect 15678 10308 15682 10364
rect 15618 10304 15682 10308
rect 15698 10364 15762 10368
rect 15698 10308 15702 10364
rect 15702 10308 15758 10364
rect 15758 10308 15762 10364
rect 15698 10304 15762 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 4698 9820 4762 9824
rect 4698 9764 4702 9820
rect 4702 9764 4758 9820
rect 4758 9764 4762 9820
rect 4698 9760 4762 9764
rect 4778 9820 4842 9824
rect 4778 9764 4782 9820
rect 4782 9764 4838 9820
rect 4838 9764 4842 9820
rect 4778 9760 4842 9764
rect 4858 9820 4922 9824
rect 4858 9764 4862 9820
rect 4862 9764 4918 9820
rect 4918 9764 4922 9820
rect 4858 9760 4922 9764
rect 11952 9820 12016 9824
rect 11952 9764 11956 9820
rect 11956 9764 12012 9820
rect 12012 9764 12016 9820
rect 11952 9760 12016 9764
rect 12032 9820 12096 9824
rect 12032 9764 12036 9820
rect 12036 9764 12092 9820
rect 12092 9764 12096 9820
rect 12032 9760 12096 9764
rect 12112 9820 12176 9824
rect 12112 9764 12116 9820
rect 12116 9764 12172 9820
rect 12172 9764 12176 9820
rect 12112 9760 12176 9764
rect 12192 9820 12256 9824
rect 12192 9764 12196 9820
rect 12196 9764 12252 9820
rect 12252 9764 12256 9820
rect 12192 9760 12256 9764
rect 19285 9820 19349 9824
rect 19285 9764 19289 9820
rect 19289 9764 19345 9820
rect 19345 9764 19349 9820
rect 19285 9760 19349 9764
rect 19365 9820 19429 9824
rect 19365 9764 19369 9820
rect 19369 9764 19425 9820
rect 19425 9764 19429 9820
rect 19365 9760 19429 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 8285 9276 8349 9280
rect 8285 9220 8289 9276
rect 8289 9220 8345 9276
rect 8345 9220 8349 9276
rect 8285 9216 8349 9220
rect 8365 9276 8429 9280
rect 8365 9220 8369 9276
rect 8369 9220 8425 9276
rect 8425 9220 8429 9276
rect 8365 9216 8429 9220
rect 8445 9276 8509 9280
rect 8445 9220 8449 9276
rect 8449 9220 8505 9276
rect 8505 9220 8509 9276
rect 8445 9216 8509 9220
rect 8525 9276 8589 9280
rect 8525 9220 8529 9276
rect 8529 9220 8585 9276
rect 8585 9220 8589 9276
rect 8525 9216 8589 9220
rect 15618 9276 15682 9280
rect 15618 9220 15622 9276
rect 15622 9220 15678 9276
rect 15678 9220 15682 9276
rect 15618 9216 15682 9220
rect 15698 9276 15762 9280
rect 15698 9220 15702 9276
rect 15702 9220 15758 9276
rect 15758 9220 15762 9276
rect 15698 9216 15762 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 5212 8876 5276 8940
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 4698 8732 4762 8736
rect 4698 8676 4702 8732
rect 4702 8676 4758 8732
rect 4758 8676 4762 8732
rect 4698 8672 4762 8676
rect 4778 8732 4842 8736
rect 4778 8676 4782 8732
rect 4782 8676 4838 8732
rect 4838 8676 4842 8732
rect 4778 8672 4842 8676
rect 4858 8732 4922 8736
rect 4858 8676 4862 8732
rect 4862 8676 4918 8732
rect 4918 8676 4922 8732
rect 4858 8672 4922 8676
rect 11952 8732 12016 8736
rect 11952 8676 11956 8732
rect 11956 8676 12012 8732
rect 12012 8676 12016 8732
rect 11952 8672 12016 8676
rect 12032 8732 12096 8736
rect 12032 8676 12036 8732
rect 12036 8676 12092 8732
rect 12092 8676 12096 8732
rect 12032 8672 12096 8676
rect 12112 8732 12176 8736
rect 12112 8676 12116 8732
rect 12116 8676 12172 8732
rect 12172 8676 12176 8732
rect 12112 8672 12176 8676
rect 12192 8732 12256 8736
rect 12192 8676 12196 8732
rect 12196 8676 12252 8732
rect 12252 8676 12256 8732
rect 12192 8672 12256 8676
rect 19285 8732 19349 8736
rect 19285 8676 19289 8732
rect 19289 8676 19345 8732
rect 19345 8676 19349 8732
rect 19285 8672 19349 8676
rect 19365 8732 19429 8736
rect 19365 8676 19369 8732
rect 19369 8676 19425 8732
rect 19425 8676 19429 8732
rect 19365 8672 19429 8676
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 8285 8188 8349 8192
rect 8285 8132 8289 8188
rect 8289 8132 8345 8188
rect 8345 8132 8349 8188
rect 8285 8128 8349 8132
rect 8365 8188 8429 8192
rect 8365 8132 8369 8188
rect 8369 8132 8425 8188
rect 8425 8132 8429 8188
rect 8365 8128 8429 8132
rect 8445 8188 8509 8192
rect 8445 8132 8449 8188
rect 8449 8132 8505 8188
rect 8505 8132 8509 8188
rect 8445 8128 8509 8132
rect 8525 8188 8589 8192
rect 8525 8132 8529 8188
rect 8529 8132 8585 8188
rect 8585 8132 8589 8188
rect 8525 8128 8589 8132
rect 15618 8188 15682 8192
rect 15618 8132 15622 8188
rect 15622 8132 15678 8188
rect 15678 8132 15682 8188
rect 15618 8128 15682 8132
rect 15698 8188 15762 8192
rect 15698 8132 15702 8188
rect 15702 8132 15758 8188
rect 15758 8132 15762 8188
rect 15698 8128 15762 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 4698 7644 4762 7648
rect 4698 7588 4702 7644
rect 4702 7588 4758 7644
rect 4758 7588 4762 7644
rect 4698 7584 4762 7588
rect 4778 7644 4842 7648
rect 4778 7588 4782 7644
rect 4782 7588 4838 7644
rect 4838 7588 4842 7644
rect 4778 7584 4842 7588
rect 4858 7644 4922 7648
rect 4858 7588 4862 7644
rect 4862 7588 4918 7644
rect 4918 7588 4922 7644
rect 4858 7584 4922 7588
rect 11952 7644 12016 7648
rect 11952 7588 11956 7644
rect 11956 7588 12012 7644
rect 12012 7588 12016 7644
rect 11952 7584 12016 7588
rect 12032 7644 12096 7648
rect 12032 7588 12036 7644
rect 12036 7588 12092 7644
rect 12092 7588 12096 7644
rect 12032 7584 12096 7588
rect 12112 7644 12176 7648
rect 12112 7588 12116 7644
rect 12116 7588 12172 7644
rect 12172 7588 12176 7644
rect 12112 7584 12176 7588
rect 12192 7644 12256 7648
rect 12192 7588 12196 7644
rect 12196 7588 12252 7644
rect 12252 7588 12256 7644
rect 12192 7584 12256 7588
rect 19285 7644 19349 7648
rect 19285 7588 19289 7644
rect 19289 7588 19345 7644
rect 19345 7588 19349 7644
rect 19285 7584 19349 7588
rect 19365 7644 19429 7648
rect 19365 7588 19369 7644
rect 19369 7588 19425 7644
rect 19425 7588 19429 7644
rect 19365 7584 19429 7588
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 8285 7100 8349 7104
rect 8285 7044 8289 7100
rect 8289 7044 8345 7100
rect 8345 7044 8349 7100
rect 8285 7040 8349 7044
rect 8365 7100 8429 7104
rect 8365 7044 8369 7100
rect 8369 7044 8425 7100
rect 8425 7044 8429 7100
rect 8365 7040 8429 7044
rect 8445 7100 8509 7104
rect 8445 7044 8449 7100
rect 8449 7044 8505 7100
rect 8505 7044 8509 7100
rect 8445 7040 8509 7044
rect 8525 7100 8589 7104
rect 8525 7044 8529 7100
rect 8529 7044 8585 7100
rect 8585 7044 8589 7100
rect 8525 7040 8589 7044
rect 15618 7100 15682 7104
rect 15618 7044 15622 7100
rect 15622 7044 15678 7100
rect 15678 7044 15682 7100
rect 15618 7040 15682 7044
rect 15698 7100 15762 7104
rect 15698 7044 15702 7100
rect 15702 7044 15758 7100
rect 15758 7044 15762 7100
rect 15698 7040 15762 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 4698 6556 4762 6560
rect 4698 6500 4702 6556
rect 4702 6500 4758 6556
rect 4758 6500 4762 6556
rect 4698 6496 4762 6500
rect 4778 6556 4842 6560
rect 4778 6500 4782 6556
rect 4782 6500 4838 6556
rect 4838 6500 4842 6556
rect 4778 6496 4842 6500
rect 4858 6556 4922 6560
rect 4858 6500 4862 6556
rect 4862 6500 4918 6556
rect 4918 6500 4922 6556
rect 4858 6496 4922 6500
rect 11952 6556 12016 6560
rect 11952 6500 11956 6556
rect 11956 6500 12012 6556
rect 12012 6500 12016 6556
rect 11952 6496 12016 6500
rect 12032 6556 12096 6560
rect 12032 6500 12036 6556
rect 12036 6500 12092 6556
rect 12092 6500 12096 6556
rect 12032 6496 12096 6500
rect 12112 6556 12176 6560
rect 12112 6500 12116 6556
rect 12116 6500 12172 6556
rect 12172 6500 12176 6556
rect 12112 6496 12176 6500
rect 12192 6556 12256 6560
rect 12192 6500 12196 6556
rect 12196 6500 12252 6556
rect 12252 6500 12256 6556
rect 12192 6496 12256 6500
rect 19285 6556 19349 6560
rect 19285 6500 19289 6556
rect 19289 6500 19345 6556
rect 19345 6500 19349 6556
rect 19285 6496 19349 6500
rect 19365 6556 19429 6560
rect 19365 6500 19369 6556
rect 19369 6500 19425 6556
rect 19425 6500 19429 6556
rect 19365 6496 19429 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 8285 6012 8349 6016
rect 8285 5956 8289 6012
rect 8289 5956 8345 6012
rect 8345 5956 8349 6012
rect 8285 5952 8349 5956
rect 8365 6012 8429 6016
rect 8365 5956 8369 6012
rect 8369 5956 8425 6012
rect 8425 5956 8429 6012
rect 8365 5952 8429 5956
rect 8445 6012 8509 6016
rect 8445 5956 8449 6012
rect 8449 5956 8505 6012
rect 8505 5956 8509 6012
rect 8445 5952 8509 5956
rect 8525 6012 8589 6016
rect 8525 5956 8529 6012
rect 8529 5956 8585 6012
rect 8585 5956 8589 6012
rect 8525 5952 8589 5956
rect 15618 6012 15682 6016
rect 15618 5956 15622 6012
rect 15622 5956 15678 6012
rect 15678 5956 15682 6012
rect 15618 5952 15682 5956
rect 15698 6012 15762 6016
rect 15698 5956 15702 6012
rect 15702 5956 15758 6012
rect 15758 5956 15762 6012
rect 15698 5952 15762 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 4698 5468 4762 5472
rect 4698 5412 4702 5468
rect 4702 5412 4758 5468
rect 4758 5412 4762 5468
rect 4698 5408 4762 5412
rect 4778 5468 4842 5472
rect 4778 5412 4782 5468
rect 4782 5412 4838 5468
rect 4838 5412 4842 5468
rect 4778 5408 4842 5412
rect 4858 5468 4922 5472
rect 4858 5412 4862 5468
rect 4862 5412 4918 5468
rect 4918 5412 4922 5468
rect 4858 5408 4922 5412
rect 11952 5468 12016 5472
rect 11952 5412 11956 5468
rect 11956 5412 12012 5468
rect 12012 5412 12016 5468
rect 11952 5408 12016 5412
rect 12032 5468 12096 5472
rect 12032 5412 12036 5468
rect 12036 5412 12092 5468
rect 12092 5412 12096 5468
rect 12032 5408 12096 5412
rect 12112 5468 12176 5472
rect 12112 5412 12116 5468
rect 12116 5412 12172 5468
rect 12172 5412 12176 5468
rect 12112 5408 12176 5412
rect 12192 5468 12256 5472
rect 12192 5412 12196 5468
rect 12196 5412 12252 5468
rect 12252 5412 12256 5468
rect 12192 5408 12256 5412
rect 19285 5468 19349 5472
rect 19285 5412 19289 5468
rect 19289 5412 19345 5468
rect 19345 5412 19349 5468
rect 19285 5408 19349 5412
rect 19365 5468 19429 5472
rect 19365 5412 19369 5468
rect 19369 5412 19425 5468
rect 19425 5412 19429 5468
rect 19365 5408 19429 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 8285 4924 8349 4928
rect 8285 4868 8289 4924
rect 8289 4868 8345 4924
rect 8345 4868 8349 4924
rect 8285 4864 8349 4868
rect 8365 4924 8429 4928
rect 8365 4868 8369 4924
rect 8369 4868 8425 4924
rect 8425 4868 8429 4924
rect 8365 4864 8429 4868
rect 8445 4924 8509 4928
rect 8445 4868 8449 4924
rect 8449 4868 8505 4924
rect 8505 4868 8509 4924
rect 8445 4864 8509 4868
rect 8525 4924 8589 4928
rect 8525 4868 8529 4924
rect 8529 4868 8585 4924
rect 8585 4868 8589 4924
rect 8525 4864 8589 4868
rect 15618 4924 15682 4928
rect 15618 4868 15622 4924
rect 15622 4868 15678 4924
rect 15678 4868 15682 4924
rect 15618 4864 15682 4868
rect 15698 4924 15762 4928
rect 15698 4868 15702 4924
rect 15702 4868 15758 4924
rect 15758 4868 15762 4924
rect 15698 4864 15762 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 4698 4380 4762 4384
rect 4698 4324 4702 4380
rect 4702 4324 4758 4380
rect 4758 4324 4762 4380
rect 4698 4320 4762 4324
rect 4778 4380 4842 4384
rect 4778 4324 4782 4380
rect 4782 4324 4838 4380
rect 4838 4324 4842 4380
rect 4778 4320 4842 4324
rect 4858 4380 4922 4384
rect 4858 4324 4862 4380
rect 4862 4324 4918 4380
rect 4918 4324 4922 4380
rect 4858 4320 4922 4324
rect 11952 4380 12016 4384
rect 11952 4324 11956 4380
rect 11956 4324 12012 4380
rect 12012 4324 12016 4380
rect 11952 4320 12016 4324
rect 12032 4380 12096 4384
rect 12032 4324 12036 4380
rect 12036 4324 12092 4380
rect 12092 4324 12096 4380
rect 12032 4320 12096 4324
rect 12112 4380 12176 4384
rect 12112 4324 12116 4380
rect 12116 4324 12172 4380
rect 12172 4324 12176 4380
rect 12112 4320 12176 4324
rect 12192 4380 12256 4384
rect 12192 4324 12196 4380
rect 12196 4324 12252 4380
rect 12252 4324 12256 4380
rect 12192 4320 12256 4324
rect 19285 4380 19349 4384
rect 19285 4324 19289 4380
rect 19289 4324 19345 4380
rect 19345 4324 19349 4380
rect 19285 4320 19349 4324
rect 19365 4380 19429 4384
rect 19365 4324 19369 4380
rect 19369 4324 19425 4380
rect 19425 4324 19429 4380
rect 19365 4320 19429 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 4108 3708 4172 3772
rect 8285 3836 8349 3840
rect 8285 3780 8289 3836
rect 8289 3780 8345 3836
rect 8345 3780 8349 3836
rect 8285 3776 8349 3780
rect 8365 3836 8429 3840
rect 8365 3780 8369 3836
rect 8369 3780 8425 3836
rect 8425 3780 8429 3836
rect 8365 3776 8429 3780
rect 8445 3836 8509 3840
rect 8445 3780 8449 3836
rect 8449 3780 8505 3836
rect 8505 3780 8509 3836
rect 8445 3776 8509 3780
rect 8525 3836 8589 3840
rect 8525 3780 8529 3836
rect 8529 3780 8585 3836
rect 8585 3780 8589 3836
rect 8525 3776 8589 3780
rect 15618 3836 15682 3840
rect 15618 3780 15622 3836
rect 15622 3780 15678 3836
rect 15678 3780 15682 3836
rect 15618 3776 15682 3780
rect 15698 3836 15762 3840
rect 15698 3780 15702 3836
rect 15702 3780 15758 3836
rect 15758 3780 15762 3836
rect 15698 3776 15762 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 4698 3292 4762 3296
rect 4698 3236 4702 3292
rect 4702 3236 4758 3292
rect 4758 3236 4762 3292
rect 4698 3232 4762 3236
rect 4778 3292 4842 3296
rect 4778 3236 4782 3292
rect 4782 3236 4838 3292
rect 4838 3236 4842 3292
rect 4778 3232 4842 3236
rect 4858 3292 4922 3296
rect 4858 3236 4862 3292
rect 4862 3236 4918 3292
rect 4918 3236 4922 3292
rect 4858 3232 4922 3236
rect 11952 3292 12016 3296
rect 11952 3236 11956 3292
rect 11956 3236 12012 3292
rect 12012 3236 12016 3292
rect 11952 3232 12016 3236
rect 12032 3292 12096 3296
rect 12032 3236 12036 3292
rect 12036 3236 12092 3292
rect 12092 3236 12096 3292
rect 12032 3232 12096 3236
rect 12112 3292 12176 3296
rect 12112 3236 12116 3292
rect 12116 3236 12172 3292
rect 12172 3236 12176 3292
rect 12112 3232 12176 3236
rect 12192 3292 12256 3296
rect 12192 3236 12196 3292
rect 12196 3236 12252 3292
rect 12252 3236 12256 3292
rect 12192 3232 12256 3236
rect 19285 3292 19349 3296
rect 19285 3236 19289 3292
rect 19289 3236 19345 3292
rect 19345 3236 19349 3292
rect 19285 3232 19349 3236
rect 19365 3292 19429 3296
rect 19365 3236 19369 3292
rect 19369 3236 19425 3292
rect 19425 3236 19429 3292
rect 19365 3232 19429 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 18276 3028 18340 3092
rect 8285 2748 8349 2752
rect 8285 2692 8289 2748
rect 8289 2692 8345 2748
rect 8345 2692 8349 2748
rect 8285 2688 8349 2692
rect 8365 2748 8429 2752
rect 8365 2692 8369 2748
rect 8369 2692 8425 2748
rect 8425 2692 8429 2748
rect 8365 2688 8429 2692
rect 8445 2748 8509 2752
rect 8445 2692 8449 2748
rect 8449 2692 8505 2748
rect 8505 2692 8509 2748
rect 8445 2688 8509 2692
rect 8525 2748 8589 2752
rect 8525 2692 8529 2748
rect 8529 2692 8585 2748
rect 8585 2692 8589 2748
rect 8525 2688 8589 2692
rect 15618 2748 15682 2752
rect 15618 2692 15622 2748
rect 15622 2692 15678 2748
rect 15678 2692 15682 2748
rect 15618 2688 15682 2692
rect 15698 2748 15762 2752
rect 15698 2692 15702 2748
rect 15702 2692 15758 2748
rect 15758 2692 15762 2748
rect 15698 2688 15762 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 4698 2204 4762 2208
rect 4698 2148 4702 2204
rect 4702 2148 4758 2204
rect 4758 2148 4762 2204
rect 4698 2144 4762 2148
rect 4778 2204 4842 2208
rect 4778 2148 4782 2204
rect 4782 2148 4838 2204
rect 4838 2148 4842 2204
rect 4778 2144 4842 2148
rect 4858 2204 4922 2208
rect 4858 2148 4862 2204
rect 4862 2148 4918 2204
rect 4918 2148 4922 2204
rect 4858 2144 4922 2148
rect 11952 2204 12016 2208
rect 11952 2148 11956 2204
rect 11956 2148 12012 2204
rect 12012 2148 12016 2204
rect 11952 2144 12016 2148
rect 12032 2204 12096 2208
rect 12032 2148 12036 2204
rect 12036 2148 12092 2204
rect 12092 2148 12096 2204
rect 12032 2144 12096 2148
rect 12112 2204 12176 2208
rect 12112 2148 12116 2204
rect 12116 2148 12172 2204
rect 12172 2148 12176 2204
rect 12112 2144 12176 2148
rect 12192 2204 12256 2208
rect 12192 2148 12196 2204
rect 12196 2148 12252 2204
rect 12252 2148 12256 2204
rect 12192 2144 12256 2148
rect 19285 2204 19349 2208
rect 19285 2148 19289 2204
rect 19289 2148 19345 2204
rect 19345 2148 19349 2204
rect 19285 2144 19349 2148
rect 19365 2204 19429 2208
rect 19365 2148 19369 2204
rect 19369 2148 19425 2204
rect 19425 2148 19429 2204
rect 19365 2144 19429 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 5212 1532 5276 1596
<< metal4 >>
rect 4610 19616 4931 19632
rect 4610 19552 4618 19616
rect 4682 19552 4698 19616
rect 4762 19552 4778 19616
rect 4842 19552 4858 19616
rect 4922 19552 4931 19616
rect 4610 18528 4931 19552
rect 4610 18464 4618 18528
rect 4682 18464 4698 18528
rect 4762 18464 4778 18528
rect 4842 18464 4858 18528
rect 4922 18464 4931 18528
rect 4610 17440 4931 18464
rect 4610 17376 4618 17440
rect 4682 17376 4698 17440
rect 4762 17376 4778 17440
rect 4842 17376 4858 17440
rect 4922 17376 4931 17440
rect 4610 16352 4931 17376
rect 4610 16288 4618 16352
rect 4682 16288 4698 16352
rect 4762 16288 4778 16352
rect 4842 16288 4858 16352
rect 4922 16288 4931 16352
rect 4610 15264 4931 16288
rect 4610 15200 4618 15264
rect 4682 15200 4698 15264
rect 4762 15200 4778 15264
rect 4842 15200 4858 15264
rect 4922 15200 4931 15264
rect 4610 14176 4931 15200
rect 4610 14112 4618 14176
rect 4682 14112 4698 14176
rect 4762 14112 4778 14176
rect 4842 14112 4858 14176
rect 4922 14112 4931 14176
rect 4610 13088 4931 14112
rect 4610 13024 4618 13088
rect 4682 13024 4698 13088
rect 4762 13024 4778 13088
rect 4842 13024 4858 13088
rect 4922 13024 4931 13088
rect 4610 12000 4931 13024
rect 4610 11936 4618 12000
rect 4682 11936 4698 12000
rect 4762 11936 4778 12000
rect 4842 11936 4858 12000
rect 4922 11936 4931 12000
rect 4610 10912 4931 11936
rect 4610 10848 4618 10912
rect 4682 10848 4698 10912
rect 4762 10848 4778 10912
rect 4842 10848 4858 10912
rect 4922 10848 4931 10912
rect 4610 9824 4931 10848
rect 4610 9760 4618 9824
rect 4682 9760 4698 9824
rect 4762 9760 4778 9824
rect 4842 9760 4858 9824
rect 4922 9760 4931 9824
rect 4610 8736 4931 9760
rect 8277 19072 8597 19632
rect 8277 19008 8285 19072
rect 8349 19008 8365 19072
rect 8429 19008 8445 19072
rect 8509 19008 8525 19072
rect 8589 19008 8597 19072
rect 8277 17984 8597 19008
rect 8277 17920 8285 17984
rect 8349 17920 8365 17984
rect 8429 17920 8445 17984
rect 8509 17920 8525 17984
rect 8589 17920 8597 17984
rect 8277 16896 8597 17920
rect 8277 16832 8285 16896
rect 8349 16832 8365 16896
rect 8429 16832 8445 16896
rect 8509 16832 8525 16896
rect 8589 16832 8597 16896
rect 8277 15808 8597 16832
rect 8277 15744 8285 15808
rect 8349 15744 8365 15808
rect 8429 15744 8445 15808
rect 8509 15744 8525 15808
rect 8589 15744 8597 15808
rect 8277 14720 8597 15744
rect 8277 14656 8285 14720
rect 8349 14656 8365 14720
rect 8429 14656 8445 14720
rect 8509 14656 8525 14720
rect 8589 14656 8597 14720
rect 8277 13632 8597 14656
rect 8277 13568 8285 13632
rect 8349 13568 8365 13632
rect 8429 13568 8445 13632
rect 8509 13568 8525 13632
rect 8589 13568 8597 13632
rect 8277 12544 8597 13568
rect 8277 12480 8285 12544
rect 8349 12480 8365 12544
rect 8429 12480 8445 12544
rect 8509 12480 8525 12544
rect 8589 12480 8597 12544
rect 8277 11456 8597 12480
rect 8277 11392 8285 11456
rect 8349 11392 8365 11456
rect 8429 11392 8445 11456
rect 8509 11392 8525 11456
rect 8589 11392 8597 11456
rect 8277 10368 8597 11392
rect 8277 10304 8285 10368
rect 8349 10304 8365 10368
rect 8429 10304 8445 10368
rect 8509 10304 8525 10368
rect 8589 10304 8597 10368
rect 8277 9280 8597 10304
rect 8277 9216 8285 9280
rect 8349 9216 8365 9280
rect 8429 9216 8445 9280
rect 8509 9216 8525 9280
rect 8589 9216 8597 9280
rect 5211 8940 5277 8941
rect 5211 8876 5212 8940
rect 5276 8876 5277 8940
rect 5211 8875 5277 8876
rect 4610 8672 4618 8736
rect 4682 8672 4698 8736
rect 4762 8672 4778 8736
rect 4842 8672 4858 8736
rect 4922 8672 4931 8736
rect 4610 7648 4931 8672
rect 4610 7584 4618 7648
rect 4682 7584 4698 7648
rect 4762 7584 4778 7648
rect 4842 7584 4858 7648
rect 4922 7584 4931 7648
rect 4610 6560 4931 7584
rect 4610 6496 4618 6560
rect 4682 6496 4698 6560
rect 4762 6496 4778 6560
rect 4842 6496 4858 6560
rect 4922 6496 4931 6560
rect 4610 5472 4931 6496
rect 4610 5408 4618 5472
rect 4682 5408 4698 5472
rect 4762 5408 4778 5472
rect 4842 5408 4858 5472
rect 4922 5408 4931 5472
rect 4610 4384 4931 5408
rect 4610 4320 4618 4384
rect 4682 4320 4698 4384
rect 4762 4320 4778 4384
rect 4842 4320 4858 4384
rect 4922 4320 4931 4384
rect 4107 3772 4173 3773
rect 4107 3708 4108 3772
rect 4172 3708 4173 3772
rect 4107 3707 4173 3708
rect 4110 3178 4170 3707
rect 4610 3296 4931 4320
rect 4610 3232 4618 3296
rect 4682 3232 4698 3296
rect 4762 3232 4778 3296
rect 4842 3232 4858 3296
rect 4922 3232 4931 3296
rect 4610 2208 4931 3232
rect 4610 2144 4618 2208
rect 4682 2144 4698 2208
rect 4762 2144 4778 2208
rect 4842 2144 4858 2208
rect 4922 2144 4931 2208
rect 4610 2128 4931 2144
rect 5214 1597 5274 8875
rect 8277 8192 8597 9216
rect 8277 8128 8285 8192
rect 8349 8128 8365 8192
rect 8429 8128 8445 8192
rect 8509 8128 8525 8192
rect 8589 8128 8597 8192
rect 8277 7104 8597 8128
rect 8277 7040 8285 7104
rect 8349 7040 8365 7104
rect 8429 7040 8445 7104
rect 8509 7040 8525 7104
rect 8589 7040 8597 7104
rect 8277 6016 8597 7040
rect 8277 5952 8285 6016
rect 8349 5952 8365 6016
rect 8429 5952 8445 6016
rect 8509 5952 8525 6016
rect 8589 5952 8597 6016
rect 8277 4928 8597 5952
rect 8277 4864 8285 4928
rect 8349 4864 8365 4928
rect 8429 4864 8445 4928
rect 8509 4864 8525 4928
rect 8589 4864 8597 4928
rect 8277 3840 8597 4864
rect 8277 3776 8285 3840
rect 8349 3776 8365 3840
rect 8429 3776 8445 3840
rect 8509 3776 8525 3840
rect 8589 3776 8597 3840
rect 8277 2752 8597 3776
rect 8277 2688 8285 2752
rect 8349 2688 8365 2752
rect 8429 2688 8445 2752
rect 8509 2688 8525 2752
rect 8589 2688 8597 2752
rect 8277 2128 8597 2688
rect 11944 19616 12264 19632
rect 11944 19552 11952 19616
rect 12016 19552 12032 19616
rect 12096 19552 12112 19616
rect 12176 19552 12192 19616
rect 12256 19552 12264 19616
rect 11944 18528 12264 19552
rect 11944 18464 11952 18528
rect 12016 18464 12032 18528
rect 12096 18464 12112 18528
rect 12176 18464 12192 18528
rect 12256 18464 12264 18528
rect 11944 17440 12264 18464
rect 11944 17376 11952 17440
rect 12016 17376 12032 17440
rect 12096 17376 12112 17440
rect 12176 17376 12192 17440
rect 12256 17376 12264 17440
rect 11944 16352 12264 17376
rect 11944 16288 11952 16352
rect 12016 16288 12032 16352
rect 12096 16288 12112 16352
rect 12176 16288 12192 16352
rect 12256 16288 12264 16352
rect 11944 15264 12264 16288
rect 11944 15200 11952 15264
rect 12016 15200 12032 15264
rect 12096 15200 12112 15264
rect 12176 15200 12192 15264
rect 12256 15200 12264 15264
rect 11944 14176 12264 15200
rect 11944 14112 11952 14176
rect 12016 14112 12032 14176
rect 12096 14112 12112 14176
rect 12176 14112 12192 14176
rect 12256 14112 12264 14176
rect 11944 13088 12264 14112
rect 11944 13024 11952 13088
rect 12016 13024 12032 13088
rect 12096 13024 12112 13088
rect 12176 13024 12192 13088
rect 12256 13024 12264 13088
rect 11944 12000 12264 13024
rect 11944 11936 11952 12000
rect 12016 11936 12032 12000
rect 12096 11936 12112 12000
rect 12176 11936 12192 12000
rect 12256 11936 12264 12000
rect 11944 10912 12264 11936
rect 11944 10848 11952 10912
rect 12016 10848 12032 10912
rect 12096 10848 12112 10912
rect 12176 10848 12192 10912
rect 12256 10848 12264 10912
rect 11944 9824 12264 10848
rect 11944 9760 11952 9824
rect 12016 9760 12032 9824
rect 12096 9760 12112 9824
rect 12176 9760 12192 9824
rect 12256 9760 12264 9824
rect 11944 8736 12264 9760
rect 11944 8672 11952 8736
rect 12016 8672 12032 8736
rect 12096 8672 12112 8736
rect 12176 8672 12192 8736
rect 12256 8672 12264 8736
rect 11944 7648 12264 8672
rect 11944 7584 11952 7648
rect 12016 7584 12032 7648
rect 12096 7584 12112 7648
rect 12176 7584 12192 7648
rect 12256 7584 12264 7648
rect 11944 6560 12264 7584
rect 11944 6496 11952 6560
rect 12016 6496 12032 6560
rect 12096 6496 12112 6560
rect 12176 6496 12192 6560
rect 12256 6496 12264 6560
rect 11944 5472 12264 6496
rect 11944 5408 11952 5472
rect 12016 5408 12032 5472
rect 12096 5408 12112 5472
rect 12176 5408 12192 5472
rect 12256 5408 12264 5472
rect 11944 4384 12264 5408
rect 11944 4320 11952 4384
rect 12016 4320 12032 4384
rect 12096 4320 12112 4384
rect 12176 4320 12192 4384
rect 12256 4320 12264 4384
rect 11944 3296 12264 4320
rect 11944 3232 11952 3296
rect 12016 3232 12032 3296
rect 12096 3232 12112 3296
rect 12176 3232 12192 3296
rect 12256 3232 12264 3296
rect 11944 2208 12264 3232
rect 11944 2144 11952 2208
rect 12016 2144 12032 2208
rect 12096 2144 12112 2208
rect 12176 2144 12192 2208
rect 12256 2144 12264 2208
rect 11944 2128 12264 2144
rect 15610 19072 15930 19632
rect 15610 19008 15618 19072
rect 15682 19008 15698 19072
rect 15762 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15930 19072
rect 15610 17984 15930 19008
rect 15610 17920 15618 17984
rect 15682 17920 15698 17984
rect 15762 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15930 17984
rect 15610 16896 15930 17920
rect 15610 16832 15618 16896
rect 15682 16832 15698 16896
rect 15762 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15930 16896
rect 15610 15808 15930 16832
rect 15610 15744 15618 15808
rect 15682 15744 15698 15808
rect 15762 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15930 15808
rect 15610 14720 15930 15744
rect 15610 14656 15618 14720
rect 15682 14656 15698 14720
rect 15762 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15930 14720
rect 15610 13632 15930 14656
rect 15610 13568 15618 13632
rect 15682 13568 15698 13632
rect 15762 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15930 13632
rect 15610 12544 15930 13568
rect 15610 12480 15618 12544
rect 15682 12480 15698 12544
rect 15762 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15930 12544
rect 15610 11456 15930 12480
rect 15610 11392 15618 11456
rect 15682 11392 15698 11456
rect 15762 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15930 11456
rect 15610 10368 15930 11392
rect 15610 10304 15618 10368
rect 15682 10304 15698 10368
rect 15762 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15930 10368
rect 15610 9280 15930 10304
rect 15610 9216 15618 9280
rect 15682 9216 15698 9280
rect 15762 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15930 9280
rect 15610 8192 15930 9216
rect 15610 8128 15618 8192
rect 15682 8128 15698 8192
rect 15762 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15930 8192
rect 15610 7104 15930 8128
rect 15610 7040 15618 7104
rect 15682 7040 15698 7104
rect 15762 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15930 7104
rect 15610 6016 15930 7040
rect 15610 5952 15618 6016
rect 15682 5952 15698 6016
rect 15762 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15930 6016
rect 15610 4928 15930 5952
rect 15610 4864 15618 4928
rect 15682 4864 15698 4928
rect 15762 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15930 4928
rect 15610 3840 15930 4864
rect 15610 3776 15618 3840
rect 15682 3776 15698 3840
rect 15762 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15930 3840
rect 15610 2752 15930 3776
rect 19277 19616 19597 19632
rect 19277 19552 19285 19616
rect 19349 19552 19365 19616
rect 19429 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19597 19616
rect 19277 18528 19597 19552
rect 19277 18464 19285 18528
rect 19349 18464 19365 18528
rect 19429 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19597 18528
rect 19277 17440 19597 18464
rect 19277 17376 19285 17440
rect 19349 17376 19365 17440
rect 19429 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19597 17440
rect 19277 16352 19597 17376
rect 19277 16288 19285 16352
rect 19349 16288 19365 16352
rect 19429 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19597 16352
rect 19277 15264 19597 16288
rect 19277 15200 19285 15264
rect 19349 15200 19365 15264
rect 19429 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19597 15264
rect 19277 14176 19597 15200
rect 19277 14112 19285 14176
rect 19349 14112 19365 14176
rect 19429 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19597 14176
rect 19277 13088 19597 14112
rect 21587 13836 21653 13837
rect 21587 13772 21588 13836
rect 21652 13772 21653 13836
rect 21587 13771 21653 13772
rect 21590 13565 21650 13771
rect 21587 13564 21653 13565
rect 21587 13500 21588 13564
rect 21652 13500 21653 13564
rect 21587 13499 21653 13500
rect 19277 13024 19285 13088
rect 19349 13024 19365 13088
rect 19429 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19597 13088
rect 19277 12000 19597 13024
rect 19277 11936 19285 12000
rect 19349 11936 19365 12000
rect 19429 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19597 12000
rect 19277 10912 19597 11936
rect 21403 11252 21469 11253
rect 21403 11188 21404 11252
rect 21468 11250 21469 11252
rect 21468 11190 21650 11250
rect 21468 11188 21469 11190
rect 21403 11187 21469 11188
rect 21590 11117 21650 11190
rect 21587 11116 21653 11117
rect 21587 11052 21588 11116
rect 21652 11052 21653 11116
rect 21587 11051 21653 11052
rect 19277 10848 19285 10912
rect 19349 10848 19365 10912
rect 19429 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19597 10912
rect 19277 9824 19597 10848
rect 19277 9760 19285 9824
rect 19349 9760 19365 9824
rect 19429 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19597 9824
rect 19277 8736 19597 9760
rect 19277 8672 19285 8736
rect 19349 8672 19365 8736
rect 19429 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19597 8736
rect 19277 7648 19597 8672
rect 19277 7584 19285 7648
rect 19349 7584 19365 7648
rect 19429 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19597 7648
rect 19277 6560 19597 7584
rect 19277 6496 19285 6560
rect 19349 6496 19365 6560
rect 19429 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19597 6560
rect 19277 5472 19597 6496
rect 19277 5408 19285 5472
rect 19349 5408 19365 5472
rect 19429 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19597 5472
rect 19277 4384 19597 5408
rect 19277 4320 19285 4384
rect 19349 4320 19365 4384
rect 19429 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19597 4384
rect 19277 3296 19597 4320
rect 19277 3232 19285 3296
rect 19349 3232 19365 3296
rect 19429 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19597 3296
rect 15610 2688 15618 2752
rect 15682 2688 15698 2752
rect 15762 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15930 2752
rect 15610 2128 15930 2688
rect 19277 2208 19597 3232
rect 19277 2144 19285 2208
rect 19349 2144 19365 2208
rect 19429 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19597 2208
rect 19277 2128 19597 2144
rect 5211 1596 5277 1597
rect 5211 1532 5212 1596
rect 5276 1532 5277 1596
rect 5211 1531 5277 1532
<< via4 >>
rect 4022 2942 4258 3178
rect 18190 3092 18426 3178
rect 18190 3028 18276 3092
rect 18276 3028 18340 3092
rect 18340 3028 18426 3092
rect 18190 2942 18426 3028
<< metal5 >>
rect 3980 3178 18468 3220
rect 3980 2942 4022 3178
rect 4258 2942 18190 3178
rect 18426 2942 18468 3178
rect 3980 2900 18468 2942
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__44__D
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor4_4  _49_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_28
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__47__B
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__C
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__C
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _48_
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 1602 592
use scs8hd_nor4_4  _50_
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__C
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__B
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__D
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__D
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__B
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _68_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_145 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_163 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_177 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_165 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_183
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 20884 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 20884 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 406 592
use scs8hd_or4_4  _44_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__B
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_13
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__C
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _47_
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__48__B
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__44__C
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__C
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__D
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__D
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_108
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _25_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_181
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _51_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _55_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__54__B
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__B
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__B
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__51__D
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__D
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 130 592
use scs8hd_inv_8  _32_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__B
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_or4_4  _54_
timestamp 1586364061
transform 1 0 2300 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_11
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _45_
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__46__B
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__C
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__51__C
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__D
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__B
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_112
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _56_
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _36_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 1 4896
box -38 -48 682 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__58__D
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _24_
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__46__C
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_28
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _46_
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__C
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__D
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_100
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _33_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 20884 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use scs8hd_or4_4  _37_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use scs8hd_nor4_4  _58_
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 1602 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _57_
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 1602 592
use scs8hd_conb_1  _61_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_37
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_37
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__C
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__B
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__39__C
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_nor4_4  _38_
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__C
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__B
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_70
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__D
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__B
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_103
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _34_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _62_
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 20884 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use scs8hd_inv_8  _23_
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__37__C
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_11
timestamp 1586364061
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _59_
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__B
timestamp 1586364061
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__B
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _39_
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_37
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_42
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__39__D
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _35_
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_115
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_139
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _41_
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 1602 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__41__C
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__B
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _53_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__B
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__C
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__B
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _29_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_12
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__B
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__B
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__B
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _40_
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__43__D
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__40__D
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__B
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _52_
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_121
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _63_
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _42_
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _27_
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__43__C
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 20884 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__D
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_8
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _43_
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__42__C
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__D
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _30_
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _28_
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _26_
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_25
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_21
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__D
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _31_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_170
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 20884 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 590 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_conb_1  _60_
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 20884 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_20
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_78
timestamp 1586364061
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 20884 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_192
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_192
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 20884 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_211
timestamp 1586364061
transform 1 0 20516 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_54
timestamp 1586364061
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_131
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_63
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_125
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_137
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_211
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 846 21520 902 22000 6 address[0]
port 0 nsew default input
rlabel metal2 s 3238 0 3294 480 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 1096 480 1216 6 address[2]
port 2 nsew default input
rlabel metal2 s 2502 21520 2558 22000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 3272 480 3392 6 address[4]
port 4 nsew default input
rlabel metal2 s 4526 0 4582 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 4158 21520 4214 22000 6 chany_bottom_in[0]
port 6 nsew default input
rlabel metal3 s 21520 1232 22000 1352 6 chany_bottom_in[1]
port 7 nsew default input
rlabel metal3 s 21520 3680 22000 3800 6 chany_bottom_in[2]
port 8 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chany_bottom_in[3]
port 9 nsew default input
rlabel metal3 s 21520 6128 22000 6248 6 chany_bottom_in[4]
port 10 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chany_bottom_in[5]
port 11 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[6]
port 12 nsew default input
rlabel metal2 s 5906 21520 5962 22000 6 chany_bottom_in[7]
port 13 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chany_bottom_in[8]
port 14 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_out[0]
port 15 nsew default tristate
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_out[1]
port 16 nsew default tristate
rlabel metal3 s 21520 8576 22000 8696 6 chany_bottom_out[2]
port 17 nsew default tristate
rlabel metal2 s 7562 21520 7618 22000 6 chany_bottom_out[3]
port 18 nsew default tristate
rlabel metal2 s 9678 0 9734 480 6 chany_bottom_out[4]
port 19 nsew default tristate
rlabel metal3 s 21520 11024 22000 11144 6 chany_bottom_out[5]
port 20 nsew default tristate
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_out[6]
port 21 nsew default tristate
rlabel metal3 s 21520 13472 22000 13592 6 chany_bottom_out[7]
port 22 nsew default tristate
rlabel metal3 s 0 12112 480 12232 6 chany_bottom_out[8]
port 23 nsew default tristate
rlabel metal2 s 9218 21520 9274 22000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 13542 0 13598 480 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 10966 21520 11022 22000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 12622 21520 12678 22000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 21520 15920 22000 16040 6 chany_top_in[7]
port 31 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 16118 0 16174 480 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal3 s 21520 18368 22000 18488 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 14370 21520 14426 22000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 16026 21520 16082 22000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 1950 0 2006 480 6 data_in
port 42 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 43 nsew default input
rlabel metal2 s 17682 21520 17738 22000 6 left_grid_pin_1_
port 44 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 left_grid_pin_5_
port 45 nsew default tristate
rlabel metal2 s 19430 21520 19486 22000 6 left_grid_pin_9_
port 46 nsew default tristate
rlabel metal2 s 21086 21520 21142 22000 6 right_grid_pin_3_
port 47 nsew default tristate
rlabel metal3 s 21520 20816 22000 20936 6 right_grid_pin_7_
port 48 nsew default tristate
rlabel metal4 s 4611 2128 4931 19632 6 vpwr
port 49 nsew default input
rlabel metal4 s 8277 2128 8597 19632 6 vgnd
port 50 nsew default input
<< end >>
