magic
tech EFS8A
magscale 1 2
timestamp 1602042181
<< locali >>
rect 2455 13345 2490 13379
rect 16715 13345 16842 13379
rect 8159 12257 8194 12291
rect 8251 11169 8286 11203
rect 10091 10081 10126 10115
rect 4077 9503 4111 9537
rect 4077 9469 4238 9503
rect 10919 8993 11046 9027
rect 6963 7905 6998 7939
rect 13495 6817 13530 6851
rect 14013 6103 14047 6409
rect 14139 5729 14266 5763
rect 19475 4641 19510 4675
rect 16451 2601 16589 2635
rect 18475 2601 18613 2635
<< viali >>
rect 18588 22049 18622 22083
rect 19625 21981 19659 22015
rect 20177 21913 20211 21947
rect 18659 21845 18693 21879
rect 17509 21641 17543 21675
rect 19165 21641 19199 21675
rect 19533 21641 19567 21675
rect 19717 21505 19751 21539
rect 20085 21505 20119 21539
rect 17024 21437 17058 21471
rect 18680 21437 18714 21471
rect 17095 21301 17129 21335
rect 18751 21301 18785 21335
rect 8125 21097 8159 21131
rect 19625 21097 19659 21131
rect 18613 21029 18647 21063
rect 1444 20961 1478 20995
rect 5156 20961 5190 20995
rect 7941 20961 7975 20995
rect 15980 20961 16014 20995
rect 16083 20893 16117 20927
rect 17049 20893 17083 20927
rect 18889 20893 18923 20927
rect 17601 20825 17635 20859
rect 1547 20757 1581 20791
rect 5227 20757 5261 20791
rect 19993 20757 20027 20791
rect 1593 20553 1627 20587
rect 1961 20553 1995 20587
rect 5273 20553 5307 20587
rect 7941 20553 7975 20587
rect 8631 20553 8665 20587
rect 15945 20553 15979 20587
rect 17095 20553 17129 20587
rect 17785 20553 17819 20587
rect 19349 20553 19383 20587
rect 19073 20485 19107 20519
rect 2237 20417 2271 20451
rect 4537 20417 4571 20451
rect 9045 20417 9079 20451
rect 13461 20417 13495 20451
rect 17509 20417 17543 20451
rect 8560 20349 8594 20383
rect 17024 20349 17058 20383
rect 18572 20349 18606 20383
rect 2881 20281 2915 20315
rect 3985 20281 4019 20315
rect 4261 20281 4295 20315
rect 13001 20281 13035 20315
rect 13185 20281 13219 20315
rect 18659 20281 18693 20315
rect 19625 20281 19659 20315
rect 20269 20281 20303 20315
rect 19625 20009 19659 20043
rect 4721 19941 4755 19975
rect 14013 19941 14047 19975
rect 18889 19941 18923 19975
rect 19752 19873 19786 19907
rect 2973 19805 3007 19839
rect 5089 19805 5123 19839
rect 13369 19805 13403 19839
rect 18245 19805 18279 19839
rect 19855 19669 19889 19703
rect 3801 19465 3835 19499
rect 5089 19465 5123 19499
rect 13553 19465 13587 19499
rect 18245 19465 18279 19499
rect 18567 19465 18601 19499
rect 18981 19465 19015 19499
rect 19533 19465 19567 19499
rect 4077 19329 4111 19363
rect 4721 19329 4755 19363
rect 13093 19329 13127 19363
rect 19717 19329 19751 19363
rect 20637 19329 20671 19363
rect 18496 19261 18530 19295
rect 20361 19193 20395 19227
rect 2513 18921 2547 18955
rect 4169 18853 4203 18887
rect 19349 18853 19383 18887
rect 2329 18785 2363 18819
rect 4445 18717 4479 18751
rect 19625 18717 19659 18751
rect 4169 18377 4203 18411
rect 19349 18377 19383 18411
rect 3801 18309 3835 18343
rect 3065 18241 3099 18275
rect 3249 18241 3283 18275
rect 2421 18037 2455 18071
rect 3019 17833 3053 17867
rect 2948 17697 2982 17731
rect 7640 17697 7674 17731
rect 7711 17493 7745 17527
rect 2973 17289 3007 17323
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 7665 17153 7699 17187
rect 8401 17153 8435 17187
rect 5156 17085 5190 17119
rect 5549 17085 5583 17119
rect 5227 16949 5261 16983
rect 6101 16677 6135 16711
rect 6745 16677 6779 16711
rect 4480 16609 4514 16643
rect 11044 16609 11078 16643
rect 4583 16405 4617 16439
rect 4905 16405 4939 16439
rect 11115 16405 11149 16439
rect 4445 16201 4479 16235
rect 6101 16201 6135 16235
rect 11345 16201 11379 16235
rect 11713 16201 11747 16235
rect 4905 16065 4939 16099
rect 10952 15997 10986 16031
rect 5549 15929 5583 15963
rect 11023 15861 11057 15895
rect 15485 15657 15519 15691
rect 5549 15589 5583 15623
rect 6469 15589 6503 15623
rect 11529 15589 11563 15623
rect 10460 15521 10494 15555
rect 14232 15521 14266 15555
rect 15301 15521 15335 15555
rect 4905 15453 4939 15487
rect 7021 15385 7055 15419
rect 12081 15385 12115 15419
rect 10563 15317 10597 15351
rect 14335 15317 14369 15351
rect 4307 15113 4341 15147
rect 5089 15113 5123 15147
rect 9689 15113 9723 15147
rect 10425 15113 10459 15147
rect 11805 15113 11839 15147
rect 12173 15113 12207 15147
rect 17509 15113 17543 15147
rect 15163 15045 15197 15079
rect 15853 15045 15887 15079
rect 5549 14977 5583 15011
rect 6377 14977 6411 15011
rect 12541 14977 12575 15011
rect 4236 14909 4270 14943
rect 4629 14909 4663 14943
rect 6904 14909 6938 14943
rect 9832 14909 9866 14943
rect 14080 14909 14114 14943
rect 14473 14909 14507 14943
rect 14841 14909 14875 14943
rect 15092 14909 15126 14943
rect 17024 14909 17058 14943
rect 5273 14841 5307 14875
rect 9919 14841 9953 14875
rect 10885 14841 10919 14875
rect 11529 14841 11563 14875
rect 13185 14841 13219 14875
rect 6975 14773 7009 14807
rect 7389 14773 7423 14807
rect 14151 14773 14185 14807
rect 15485 14773 15519 14807
rect 17095 14773 17129 14807
rect 5273 14569 5307 14603
rect 5871 14569 5905 14603
rect 10885 14569 10919 14603
rect 6837 14501 6871 14535
rect 7481 14501 7515 14535
rect 11437 14501 11471 14535
rect 12081 14501 12115 14535
rect 13001 14501 13035 14535
rect 15485 14501 15519 14535
rect 17233 14501 17267 14535
rect 1476 14433 1510 14467
rect 4756 14433 4790 14467
rect 5800 14433 5834 14467
rect 9724 14433 9758 14467
rect 13277 14365 13311 14399
rect 17877 14365 17911 14399
rect 4859 14297 4893 14331
rect 16037 14297 16071 14331
rect 1547 14229 1581 14263
rect 9827 14229 9861 14263
rect 1593 14025 1627 14059
rect 1961 14025 1995 14059
rect 4537 14025 4571 14059
rect 5825 14025 5859 14059
rect 6653 14025 6687 14059
rect 10149 14025 10183 14059
rect 11437 14025 11471 14059
rect 14013 14025 14047 14059
rect 15485 14025 15519 14059
rect 17417 14025 17451 14059
rect 6285 13957 6319 13991
rect 9413 13957 9447 13991
rect 10977 13957 11011 13991
rect 4997 13889 5031 13923
rect 7113 13889 7147 13923
rect 10425 13889 10459 13923
rect 13001 13889 13035 13923
rect 13553 13889 13587 13923
rect 14197 13889 14231 13923
rect 1409 13821 1443 13855
rect 2329 13821 2363 13855
rect 3652 13821 3686 13855
rect 4077 13821 4111 13855
rect 3755 13753 3789 13787
rect 4721 13753 4755 13787
rect 7757 13753 7791 13787
rect 8861 13753 8895 13787
rect 12265 13753 12299 13787
rect 12633 13753 12667 13787
rect 14841 13753 14875 13787
rect 16313 13753 16347 13787
rect 16497 13753 16531 13787
rect 17141 13753 17175 13787
rect 8585 13685 8619 13719
rect 9781 13685 9815 13719
rect 4261 13481 4295 13515
rect 4721 13481 4755 13515
rect 13553 13481 13587 13515
rect 15439 13481 15473 13515
rect 16911 13481 16945 13515
rect 17969 13413 18003 13447
rect 2421 13345 2455 13379
rect 4077 13345 4111 13379
rect 13369 13345 13403 13379
rect 15368 13345 15402 13379
rect 16681 13345 16715 13379
rect 1409 13277 1443 13311
rect 5457 13277 5491 13311
rect 6101 13277 6135 13311
rect 7021 13277 7055 13311
rect 7665 13277 7699 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 11713 13277 11747 13311
rect 11989 13277 12023 13311
rect 18613 13277 18647 13311
rect 2559 13141 2593 13175
rect 4353 12937 4387 12971
rect 4997 12937 5031 12971
rect 6193 12937 6227 12971
rect 9781 12937 9815 12971
rect 10103 12937 10137 12971
rect 16865 12937 16899 12971
rect 17877 12937 17911 12971
rect 19993 12937 20027 12971
rect 3939 12869 3973 12903
rect 4629 12869 4663 12903
rect 11805 12869 11839 12903
rect 5273 12801 5307 12835
rect 6653 12801 6687 12835
rect 11391 12801 11425 12835
rect 12081 12801 12115 12835
rect 14197 12801 14231 12835
rect 18613 12801 18647 12835
rect 1444 12733 1478 12767
rect 1869 12733 1903 12767
rect 3868 12733 3902 12767
rect 9020 12733 9054 12767
rect 9413 12733 9447 12767
rect 10032 12733 10066 12767
rect 10517 12733 10551 12767
rect 11288 12733 11322 12767
rect 19809 12733 19843 12767
rect 20361 12733 20395 12767
rect 2789 12665 2823 12699
rect 5917 12665 5951 12699
rect 7113 12665 7147 12699
rect 7757 12665 7791 12699
rect 12449 12665 12483 12699
rect 13277 12665 13311 12699
rect 13553 12665 13587 12699
rect 17509 12665 17543 12699
rect 18337 12665 18371 12699
rect 1547 12597 1581 12631
rect 2513 12597 2547 12631
rect 8033 12597 8067 12631
rect 9091 12597 9125 12631
rect 13001 12597 13035 12631
rect 15393 12597 15427 12631
rect 1593 12325 1627 12359
rect 9781 12325 9815 12359
rect 12909 12325 12943 12359
rect 8125 12257 8159 12291
rect 19876 12257 19910 12291
rect 1961 12189 1995 12223
rect 4629 12189 4663 12223
rect 5089 12189 5123 12223
rect 6653 12189 6687 12223
rect 7113 12189 7147 12223
rect 10057 12189 10091 12223
rect 13553 12189 13587 12223
rect 18337 12189 18371 12223
rect 18613 12189 18647 12223
rect 8263 12053 8297 12087
rect 19947 12053 19981 12087
rect 1593 11849 1627 11883
rect 3479 11849 3513 11883
rect 5365 11849 5399 11883
rect 6653 11849 6687 11883
rect 8217 11849 8251 11883
rect 9781 11849 9815 11883
rect 14519 11849 14553 11883
rect 18567 11849 18601 11883
rect 4169 11781 4203 11815
rect 7849 11781 7883 11815
rect 18337 11781 18371 11815
rect 2145 11713 2179 11747
rect 4445 11713 4479 11747
rect 5089 11713 5123 11747
rect 13553 11713 13587 11747
rect 19809 11713 19843 11747
rect 3408 11645 3442 11679
rect 14448 11645 14482 11679
rect 14841 11645 14875 11679
rect 18496 11645 18530 11679
rect 18889 11645 18923 11679
rect 1869 11577 1903 11611
rect 7113 11577 7147 11611
rect 7297 11577 7331 11611
rect 11345 11577 11379 11611
rect 12909 11577 12943 11611
rect 19349 11577 19383 11611
rect 19533 11577 19567 11611
rect 2789 11509 2823 11543
rect 3893 11509 3927 11543
rect 12633 11509 12667 11543
rect 20545 11509 20579 11543
rect 6101 11305 6135 11339
rect 8355 11305 8389 11339
rect 12909 11305 12943 11339
rect 2421 11237 2455 11271
rect 5089 11237 5123 11271
rect 11529 11237 11563 11271
rect 13093 11237 13127 11271
rect 18429 11237 18463 11271
rect 19993 11237 20027 11271
rect 7113 11169 7147 11203
rect 8217 11169 8251 11203
rect 1777 11101 1811 11135
rect 4445 11101 4479 11135
rect 11805 11101 11839 11135
rect 13553 11101 13587 11135
rect 16681 11101 16715 11135
rect 17785 11101 17819 11135
rect 19349 11101 19383 11135
rect 7297 10965 7331 10999
rect 18705 10965 18739 10999
rect 3341 10761 3375 10795
rect 4537 10761 4571 10795
rect 5227 10761 5261 10795
rect 7113 10761 7147 10795
rect 12725 10761 12759 10795
rect 17785 10761 17819 10795
rect 13553 10693 13587 10727
rect 16083 10693 16117 10727
rect 19073 10693 19107 10727
rect 20269 10693 20303 10727
rect 2421 10625 2455 10659
rect 3617 10625 3651 10659
rect 11529 10625 11563 10659
rect 17095 10625 17129 10659
rect 18153 10625 18187 10659
rect 18429 10625 18463 10659
rect 19533 10625 19567 10659
rect 19717 10625 19751 10659
rect 5156 10557 5190 10591
rect 16012 10557 16046 10591
rect 17008 10557 17042 10591
rect 17417 10557 17451 10591
rect 2053 10489 2087 10523
rect 4261 10489 4295 10523
rect 10885 10489 10919 10523
rect 12265 10489 12299 10523
rect 13001 10489 13035 10523
rect 1685 10421 1719 10455
rect 5641 10421 5675 10455
rect 8309 10421 8343 10455
rect 10609 10421 10643 10455
rect 11805 10421 11839 10455
rect 16497 10421 16531 10455
rect 10195 10217 10229 10251
rect 14289 10217 14323 10251
rect 19809 10217 19843 10251
rect 2237 10149 2271 10183
rect 10057 10081 10091 10115
rect 11488 10081 11522 10115
rect 14105 10081 14139 10115
rect 19625 10081 19659 10115
rect 4629 10013 4663 10047
rect 4905 10013 4939 10047
rect 11575 10013 11609 10047
rect 12541 10013 12575 10047
rect 12817 10013 12851 10047
rect 17877 10013 17911 10047
rect 2789 9945 2823 9979
rect 18429 9945 18463 9979
rect 2053 9877 2087 9911
rect 2329 9673 2363 9707
rect 4721 9673 4755 9707
rect 11483 9673 11517 9707
rect 14289 9673 14323 9707
rect 17877 9673 17911 9707
rect 18199 9673 18233 9707
rect 19809 9673 19843 9707
rect 20177 9673 20211 9707
rect 5319 9605 5353 9639
rect 10057 9605 10091 9639
rect 4077 9537 4111 9571
rect 4307 9537 4341 9571
rect 4997 9537 5031 9571
rect 10425 9537 10459 9571
rect 12817 9537 12851 9571
rect 14657 9537 14691 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 2513 9469 2547 9503
rect 3065 9469 3099 9503
rect 5248 9469 5282 9503
rect 8436 9469 8470 9503
rect 8861 9469 8895 9503
rect 11412 9469 11446 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 18128 9469 18162 9503
rect 19625 9469 19659 9503
rect 8539 9401 8573 9435
rect 9229 9401 9263 9435
rect 9505 9401 9539 9435
rect 12541 9401 12575 9435
rect 13461 9401 13495 9435
rect 1593 9333 1627 9367
rect 2697 9333 2731 9367
rect 5733 9333 5767 9367
rect 11805 9333 11839 9367
rect 12173 9333 12207 9367
rect 18613 9333 18647 9367
rect 19441 9333 19475 9367
rect 1547 9129 1581 9163
rect 11115 9129 11149 9163
rect 13001 9129 13035 9163
rect 13691 9129 13725 9163
rect 19809 9129 19843 9163
rect 1476 8993 1510 9027
rect 10885 8993 10919 9027
rect 13588 8993 13622 9027
rect 19625 8993 19659 9027
rect 2513 8925 2547 8959
rect 2789 8925 2823 8959
rect 4169 8925 4203 8959
rect 4629 8925 4663 8959
rect 7113 8925 7147 8959
rect 12081 8925 12115 8959
rect 12725 8925 12759 8959
rect 7665 8857 7699 8891
rect 1593 8585 1627 8619
rect 2375 8585 2409 8619
rect 3065 8585 3099 8619
rect 4261 8585 4295 8619
rect 7849 8585 7883 8619
rect 8539 8585 8573 8619
rect 18751 8585 18785 8619
rect 3893 8517 3927 8551
rect 19809 8517 19843 8551
rect 3341 8449 3375 8483
rect 4951 8449 4985 8483
rect 7573 8449 7607 8483
rect 12909 8449 12943 8483
rect 13553 8449 13587 8483
rect 15025 8449 15059 8483
rect 2304 8381 2338 8415
rect 2697 8381 2731 8415
rect 4864 8381 4898 8415
rect 8468 8381 8502 8415
rect 18680 8381 18714 8415
rect 19073 8381 19107 8415
rect 19533 8381 19567 8415
rect 19625 8381 19659 8415
rect 6653 8313 6687 8347
rect 6929 8313 6963 8347
rect 11345 8313 11379 8347
rect 12173 8313 12207 8347
rect 12633 8313 12667 8347
rect 14381 8313 14415 8347
rect 5365 8245 5399 8279
rect 8953 8245 8987 8279
rect 10977 8245 11011 8279
rect 11805 8245 11839 8279
rect 14197 8245 14231 8279
rect 20269 8245 20303 8279
rect 3341 8041 3375 8075
rect 7067 8041 7101 8075
rect 19487 8041 19521 8075
rect 2881 7973 2915 8007
rect 5825 7905 5859 7939
rect 6929 7905 6963 7939
rect 10368 7905 10402 7939
rect 19384 7905 19418 7939
rect 2237 7837 2271 7871
rect 4353 7837 4387 7871
rect 4629 7837 4663 7871
rect 10471 7837 10505 7871
rect 11437 7837 11471 7871
rect 12081 7837 12115 7871
rect 13737 7837 13771 7871
rect 15301 7837 15335 7871
rect 14289 7769 14323 7803
rect 6009 7701 6043 7735
rect 10793 7701 10827 7735
rect 1547 7497 1581 7531
rect 2237 7497 2271 7531
rect 4445 7497 4479 7531
rect 5825 7497 5859 7531
rect 10333 7497 10367 7531
rect 11529 7497 11563 7531
rect 12955 7497 12989 7531
rect 18797 7497 18831 7531
rect 13369 7429 13403 7463
rect 3985 7361 4019 7395
rect 7021 7361 7055 7395
rect 9643 7361 9677 7395
rect 10609 7361 10643 7395
rect 11069 7361 11103 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 14565 7361 14599 7395
rect 15761 7361 15795 7395
rect 19625 7361 19659 7395
rect 1444 7293 1478 7327
rect 1869 7293 1903 7327
rect 5032 7293 5066 7327
rect 5457 7293 5491 7327
rect 9540 7293 9574 7327
rect 9965 7293 9999 7327
rect 12884 7293 12918 7327
rect 15485 7225 15519 7259
rect 18245 7225 18279 7259
rect 19073 7225 19107 7259
rect 19349 7225 19383 7259
rect 5135 7157 5169 7191
rect 15209 7157 15243 7191
rect 13599 6953 13633 6987
rect 11069 6885 11103 6919
rect 13921 6885 13955 6919
rect 5181 6817 5215 6851
rect 6285 6817 6319 6851
rect 7941 6817 7975 6851
rect 13461 6817 13495 6851
rect 17300 6817 17334 6851
rect 10425 6749 10459 6783
rect 11989 6749 12023 6783
rect 12265 6749 12299 6783
rect 15301 6749 15335 6783
rect 19257 6749 19291 6783
rect 19533 6749 19567 6783
rect 5365 6613 5399 6647
rect 6469 6613 6503 6647
rect 8125 6613 8159 6647
rect 17371 6613 17405 6647
rect 5181 6409 5215 6443
rect 6285 6409 6319 6443
rect 7941 6409 7975 6443
rect 10425 6409 10459 6443
rect 10931 6409 10965 6443
rect 12909 6409 12943 6443
rect 14013 6409 14047 6443
rect 14197 6409 14231 6443
rect 17325 6409 17359 6443
rect 17785 6409 17819 6443
rect 13185 6273 13219 6307
rect 10860 6205 10894 6239
rect 13829 6137 13863 6171
rect 14749 6273 14783 6307
rect 14933 6273 14967 6307
rect 15393 6273 15427 6307
rect 18337 6273 18371 6307
rect 16472 6205 16506 6239
rect 16957 6205 16991 6239
rect 18981 6137 19015 6171
rect 11345 6069 11379 6103
rect 11897 6069 11931 6103
rect 14013 6069 14047 6103
rect 16543 6069 16577 6103
rect 19349 6069 19383 6103
rect 11207 5865 11241 5899
rect 17049 5865 17083 5899
rect 14335 5797 14369 5831
rect 11104 5729 11138 5763
rect 12081 5729 12115 5763
rect 14105 5729 14139 5763
rect 16865 5729 16899 5763
rect 15393 5661 15427 5695
rect 19349 5661 19383 5695
rect 19625 5661 19659 5695
rect 15945 5593 15979 5627
rect 12265 5525 12299 5559
rect 11069 5321 11103 5355
rect 12081 5321 12115 5355
rect 14197 5321 14231 5355
rect 14933 5321 14967 5355
rect 16865 5321 16899 5355
rect 19349 5321 19383 5355
rect 19763 5321 19797 5355
rect 20177 5321 20211 5355
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 15761 5185 15795 5219
rect 14324 5117 14358 5151
rect 19692 5117 19726 5151
rect 12817 4981 12851 5015
rect 13737 4981 13771 5015
rect 14427 4981 14461 5015
rect 13093 4709 13127 4743
rect 15301 4641 15335 4675
rect 19441 4641 19475 4675
rect 13369 4573 13403 4607
rect 17969 4573 18003 4607
rect 18245 4573 18279 4607
rect 15485 4437 15519 4471
rect 19579 4437 19613 4471
rect 13461 4233 13495 4267
rect 15301 4233 15335 4267
rect 18245 4233 18279 4267
rect 19809 4233 19843 4267
rect 10425 4165 10459 4199
rect 13185 4097 13219 4131
rect 19165 4097 19199 4131
rect 8836 4029 8870 4063
rect 9689 3961 9723 3995
rect 9873 3961 9907 3995
rect 12541 3961 12575 3995
rect 18705 3961 18739 3995
rect 18889 3961 18923 3995
rect 8907 3893 8941 3927
rect 9321 3893 9355 3927
rect 12173 3893 12207 3927
rect 16957 3893 16991 3927
rect 8585 3689 8619 3723
rect 9781 3621 9815 3655
rect 16681 3621 16715 3655
rect 17325 3621 17359 3655
rect 18245 3621 18279 3655
rect 8401 3553 8435 3587
rect 10057 3485 10091 3519
rect 11345 3485 11379 3519
rect 11621 3485 11655 3519
rect 18521 3485 18555 3519
rect 9413 3145 9447 3179
rect 18245 3145 18279 3179
rect 8723 3077 8757 3111
rect 11713 3077 11747 3111
rect 11345 3009 11379 3043
rect 17141 3009 17175 3043
rect 17417 3009 17451 3043
rect 18797 3009 18831 3043
rect 8620 2941 8654 2975
rect 9648 2941 9682 2975
rect 9735 2873 9769 2907
rect 10425 2873 10459 2907
rect 10701 2873 10735 2907
rect 16313 2873 16347 2907
rect 16497 2873 16531 2907
rect 17877 2873 17911 2907
rect 18521 2873 18555 2907
rect 8493 2805 8527 2839
rect 9137 2805 9171 2839
rect 10149 2805 10183 2839
rect 9229 2601 9263 2635
rect 16589 2601 16623 2635
rect 18613 2601 18647 2635
rect 11989 2533 12023 2567
rect 8728 2465 8762 2499
rect 8815 2465 8849 2499
rect 9781 2465 9815 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 12909 2465 12943 2499
rect 13461 2465 13495 2499
rect 16380 2465 16414 2499
rect 18404 2465 18438 2499
rect 9965 2329 9999 2363
rect 11621 2329 11655 2363
rect 13093 2329 13127 2363
rect 16865 2261 16899 2295
rect 18889 2261 18923 2295
<< metal1 >>
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 5258 24256 5264 24268
rect 4212 24228 5264 24256
rect 4212 24216 4218 24228
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 1104 22330 21436 22352
rect 1104 22278 8497 22330
rect 8549 22278 8561 22330
rect 8613 22278 8625 22330
rect 8677 22278 8689 22330
rect 8741 22278 16012 22330
rect 16064 22278 16076 22330
rect 16128 22278 16140 22330
rect 16192 22278 16204 22330
rect 16256 22278 21436 22330
rect 1104 22256 21436 22278
rect 106 22040 112 22092
rect 164 22080 170 22092
rect 15838 22080 15844 22092
rect 164 22052 15844 22080
rect 164 22040 170 22052
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 18576 22083 18634 22089
rect 18576 22049 18588 22083
rect 18622 22080 18634 22083
rect 19150 22080 19156 22092
rect 18622 22052 19156 22080
rect 18622 22049 18634 22052
rect 18576 22043 18634 22049
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19610 22012 19616 22024
rect 19571 21984 19616 22012
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 20162 21944 20168 21956
rect 20123 21916 20168 21944
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 18647 21879 18705 21885
rect 18647 21845 18659 21879
rect 18693 21876 18705 21879
rect 19334 21876 19340 21888
rect 18693 21848 19340 21876
rect 18693 21845 18705 21848
rect 18647 21839 18705 21845
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 1104 21786 21436 21808
rect 1104 21734 4739 21786
rect 4791 21734 4803 21786
rect 4855 21734 4867 21786
rect 4919 21734 4931 21786
rect 4983 21734 12255 21786
rect 12307 21734 12319 21786
rect 12371 21734 12383 21786
rect 12435 21734 12447 21786
rect 12499 21734 19770 21786
rect 19822 21734 19834 21786
rect 19886 21734 19898 21786
rect 19950 21734 19962 21786
rect 20014 21734 21436 21786
rect 1104 21712 21436 21734
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 18506 21672 18512 21684
rect 17543 21644 18512 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17012 21471 17070 21477
rect 17012 21437 17024 21471
rect 17058 21468 17070 21471
rect 17512 21468 17540 21635
rect 18506 21632 18512 21644
rect 18564 21632 18570 21684
rect 19150 21672 19156 21684
rect 19111 21644 19156 21672
rect 19150 21632 19156 21644
rect 19208 21632 19214 21684
rect 19518 21672 19524 21684
rect 19479 21644 19524 21672
rect 19518 21632 19524 21644
rect 19576 21632 19582 21684
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19392 21508 19717 21536
rect 19392 21496 19398 21508
rect 19705 21505 19717 21508
rect 19751 21505 19763 21539
rect 20070 21536 20076 21548
rect 20031 21508 20076 21536
rect 19705 21499 19763 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 17058 21440 17540 21468
rect 18668 21471 18726 21477
rect 17058 21437 17070 21440
rect 17012 21431 17070 21437
rect 18668 21437 18680 21471
rect 18714 21468 18726 21471
rect 19518 21468 19524 21480
rect 18714 21440 19524 21468
rect 18714 21437 18726 21440
rect 18668 21431 18726 21437
rect 19518 21428 19524 21440
rect 19576 21428 19582 21480
rect 17083 21335 17141 21341
rect 17083 21301 17095 21335
rect 17129 21332 17141 21335
rect 18598 21332 18604 21344
rect 17129 21304 18604 21332
rect 17129 21301 17141 21304
rect 17083 21295 17141 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 18739 21335 18797 21341
rect 18739 21301 18751 21335
rect 18785 21332 18797 21335
rect 19426 21332 19432 21344
rect 18785 21304 19432 21332
rect 18785 21301 18797 21304
rect 18739 21295 18797 21301
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 1104 21242 21436 21264
rect 1104 21190 8497 21242
rect 8549 21190 8561 21242
rect 8613 21190 8625 21242
rect 8677 21190 8689 21242
rect 8741 21190 16012 21242
rect 16064 21190 16076 21242
rect 16128 21190 16140 21242
rect 16192 21190 16204 21242
rect 16256 21190 21436 21242
rect 1104 21168 21436 21190
rect 8110 21128 8116 21140
rect 8071 21100 8116 21128
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19613 21131 19671 21137
rect 19613 21128 19625 21131
rect 19392 21100 19625 21128
rect 19392 21088 19398 21100
rect 19613 21097 19625 21100
rect 19659 21097 19671 21131
rect 19613 21091 19671 21097
rect 18598 21060 18604 21072
rect 18559 21032 18604 21060
rect 18598 21020 18604 21032
rect 18656 21020 18662 21072
rect 1302 20952 1308 21004
rect 1360 20992 1366 21004
rect 1432 20995 1490 21001
rect 1432 20992 1444 20995
rect 1360 20964 1444 20992
rect 1360 20952 1366 20964
rect 1432 20961 1444 20964
rect 1478 20961 1490 20995
rect 1432 20955 1490 20961
rect 5144 20995 5202 21001
rect 5144 20961 5156 20995
rect 5190 20992 5202 20995
rect 5258 20992 5264 21004
rect 5190 20964 5264 20992
rect 5190 20961 5202 20964
rect 5144 20955 5202 20961
rect 5258 20952 5264 20964
rect 5316 20992 5322 21004
rect 6454 20992 6460 21004
rect 5316 20964 6460 20992
rect 5316 20952 5322 20964
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 7926 20992 7932 21004
rect 7887 20964 7932 20992
rect 7926 20952 7932 20964
rect 7984 20952 7990 21004
rect 15838 20952 15844 21004
rect 15896 20992 15902 21004
rect 15968 20995 16026 21001
rect 15968 20992 15980 20995
rect 15896 20964 15980 20992
rect 15896 20952 15902 20964
rect 15968 20961 15980 20964
rect 16014 20961 16026 20995
rect 15968 20955 16026 20961
rect 16071 20927 16129 20933
rect 16071 20893 16083 20927
rect 16117 20924 16129 20927
rect 17037 20927 17095 20933
rect 17037 20924 17049 20927
rect 16117 20896 17049 20924
rect 16117 20893 16129 20896
rect 16071 20887 16129 20893
rect 17037 20893 17049 20896
rect 17083 20924 17095 20927
rect 17770 20924 17776 20936
rect 17083 20896 17776 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 18874 20924 18880 20936
rect 18835 20896 18880 20924
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 17589 20859 17647 20865
rect 17589 20825 17601 20859
rect 17635 20856 17647 20859
rect 20254 20856 20260 20868
rect 17635 20828 20260 20856
rect 17635 20825 17647 20828
rect 17589 20819 17647 20825
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 1946 20788 1952 20800
rect 1581 20760 1952 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5215 20791 5273 20797
rect 5215 20788 5227 20791
rect 5132 20760 5227 20788
rect 5132 20748 5138 20760
rect 5215 20757 5227 20760
rect 5261 20757 5273 20791
rect 5215 20751 5273 20757
rect 17494 20748 17500 20800
rect 17552 20788 17558 20800
rect 19610 20788 19616 20800
rect 17552 20760 19616 20788
rect 17552 20748 17558 20760
rect 19610 20748 19616 20760
rect 19668 20788 19674 20800
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 19668 20760 19993 20788
rect 19668 20748 19674 20760
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 19981 20751 20039 20757
rect 1104 20698 21436 20720
rect 1104 20646 4739 20698
rect 4791 20646 4803 20698
rect 4855 20646 4867 20698
rect 4919 20646 4931 20698
rect 4983 20646 12255 20698
rect 12307 20646 12319 20698
rect 12371 20646 12383 20698
rect 12435 20646 12447 20698
rect 12499 20646 19770 20698
rect 19822 20646 19834 20698
rect 19886 20646 19898 20698
rect 19950 20646 19962 20698
rect 20014 20646 21436 20698
rect 1104 20624 21436 20646
rect 1302 20544 1308 20596
rect 1360 20584 1366 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1360 20556 1593 20584
rect 1360 20544 1366 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1581 20547 1639 20553
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 5258 20584 5264 20596
rect 5219 20556 5264 20584
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 7926 20584 7932 20596
rect 7887 20556 7932 20584
rect 7926 20544 7932 20556
rect 7984 20584 7990 20596
rect 8619 20587 8677 20593
rect 8619 20584 8631 20587
rect 7984 20556 8631 20584
rect 7984 20544 7990 20556
rect 8619 20553 8631 20556
rect 8665 20553 8677 20587
rect 8619 20547 8677 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15896 20556 15945 20584
rect 15896 20544 15902 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 17083 20587 17141 20593
rect 17083 20553 17095 20587
rect 17129 20584 17141 20587
rect 17494 20584 17500 20596
rect 17129 20556 17500 20584
rect 17129 20553 17141 20556
rect 17083 20547 17141 20553
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 17770 20584 17776 20596
rect 17731 20556 17776 20584
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 19337 20587 19395 20593
rect 19337 20584 19349 20587
rect 18656 20556 19349 20584
rect 18656 20544 18662 20556
rect 19337 20553 19349 20556
rect 19383 20553 19395 20587
rect 19337 20547 19395 20553
rect 1964 20448 1992 20544
rect 19061 20519 19119 20525
rect 19061 20485 19073 20519
rect 19107 20516 19119 20519
rect 21358 20516 21364 20528
rect 19107 20488 21364 20516
rect 19107 20485 19119 20488
rect 19061 20479 19119 20485
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 1964 20420 2237 20448
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 3936 20420 4537 20448
rect 3936 20408 3942 20420
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 9033 20451 9091 20457
rect 9033 20417 9045 20451
rect 9079 20448 9091 20451
rect 9398 20448 9404 20460
rect 9079 20420 9404 20448
rect 9079 20417 9091 20420
rect 9033 20411 9091 20417
rect 8548 20383 8606 20389
rect 8548 20349 8560 20383
rect 8594 20380 8606 20383
rect 9048 20380 9076 20411
rect 9398 20408 9404 20420
rect 9456 20448 9462 20460
rect 13449 20451 13507 20457
rect 13449 20448 13461 20451
rect 9456 20420 13461 20448
rect 9456 20408 9462 20420
rect 13449 20417 13461 20420
rect 13495 20417 13507 20451
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 13449 20411 13507 20417
rect 17027 20420 17509 20448
rect 17027 20389 17055 20420
rect 17497 20417 17509 20420
rect 17543 20448 17555 20451
rect 17586 20448 17592 20460
rect 17543 20420 17592 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 8594 20352 9076 20380
rect 17012 20383 17070 20389
rect 8594 20349 8606 20352
rect 8548 20343 8606 20349
rect 17012 20349 17024 20383
rect 17058 20349 17070 20383
rect 17012 20343 17070 20349
rect 18560 20383 18618 20389
rect 18560 20349 18572 20383
rect 18606 20380 18618 20383
rect 19076 20380 19104 20479
rect 21358 20476 21364 20488
rect 21416 20476 21422 20528
rect 18606 20352 19104 20380
rect 18606 20349 18618 20352
rect 18560 20343 18618 20349
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20312 2927 20315
rect 3973 20315 4031 20321
rect 3973 20312 3985 20315
rect 2915 20284 3985 20312
rect 2915 20281 2927 20284
rect 2869 20275 2927 20281
rect 3973 20281 3985 20284
rect 4019 20312 4031 20315
rect 4249 20315 4307 20321
rect 4249 20312 4261 20315
rect 4019 20284 4261 20312
rect 4019 20281 4031 20284
rect 3973 20275 4031 20281
rect 4249 20281 4261 20284
rect 4295 20312 4307 20315
rect 7374 20312 7380 20324
rect 4295 20284 7380 20312
rect 4295 20281 4307 20284
rect 4249 20275 4307 20281
rect 7374 20272 7380 20284
rect 7432 20272 7438 20324
rect 12989 20315 13047 20321
rect 12989 20281 13001 20315
rect 13035 20312 13047 20315
rect 13170 20312 13176 20324
rect 13035 20284 13176 20312
rect 13035 20281 13047 20284
rect 12989 20275 13047 20281
rect 13170 20272 13176 20284
rect 13228 20272 13234 20324
rect 18647 20315 18705 20321
rect 18647 20281 18659 20315
rect 18693 20312 18705 20315
rect 19610 20312 19616 20324
rect 18693 20284 19616 20312
rect 18693 20281 18705 20284
rect 18647 20275 18705 20281
rect 19610 20272 19616 20284
rect 19668 20272 19674 20324
rect 20254 20312 20260 20324
rect 20215 20284 20260 20312
rect 20254 20272 20260 20284
rect 20312 20272 20318 20324
rect 1104 20154 21436 20176
rect 1104 20102 8497 20154
rect 8549 20102 8561 20154
rect 8613 20102 8625 20154
rect 8677 20102 8689 20154
rect 8741 20102 16012 20154
rect 16064 20102 16076 20154
rect 16128 20102 16140 20154
rect 16192 20102 16204 20154
rect 16256 20102 21436 20154
rect 1104 20080 21436 20102
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19972 4767 19975
rect 5074 19972 5080 19984
rect 4755 19944 5080 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 13170 19932 13176 19984
rect 13228 19972 13234 19984
rect 14001 19975 14059 19981
rect 14001 19972 14013 19975
rect 13228 19944 14013 19972
rect 13228 19932 13234 19944
rect 14001 19941 14013 19944
rect 14047 19972 14059 19975
rect 18874 19972 18880 19984
rect 14047 19944 18880 19972
rect 14047 19941 14059 19944
rect 14001 19935 14059 19941
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 19518 19864 19524 19916
rect 19576 19904 19582 19916
rect 19740 19907 19798 19913
rect 19740 19904 19752 19907
rect 19576 19876 19752 19904
rect 19576 19864 19582 19876
rect 19740 19873 19752 19876
rect 19786 19873 19798 19907
rect 19740 19867 19798 19873
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3786 19836 3792 19848
rect 3007 19808 3792 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 5074 19836 5080 19848
rect 5035 19808 5080 19836
rect 5074 19796 5080 19808
rect 5132 19796 5138 19848
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19843 19703 19901 19709
rect 19843 19700 19855 19703
rect 19392 19672 19855 19700
rect 19392 19660 19398 19672
rect 19843 19669 19855 19672
rect 19889 19669 19901 19703
rect 19843 19663 19901 19669
rect 1104 19610 21436 19632
rect 1104 19558 4739 19610
rect 4791 19558 4803 19610
rect 4855 19558 4867 19610
rect 4919 19558 4931 19610
rect 4983 19558 12255 19610
rect 12307 19558 12319 19610
rect 12371 19558 12383 19610
rect 12435 19558 12447 19610
rect 12499 19558 19770 19610
rect 19822 19558 19834 19610
rect 19886 19558 19898 19610
rect 19950 19558 19962 19610
rect 20014 19558 21436 19610
rect 1104 19536 21436 19558
rect 3786 19496 3792 19508
rect 3747 19468 3792 19496
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 5077 19499 5135 19505
rect 5077 19465 5089 19499
rect 5123 19496 5135 19499
rect 5166 19496 5172 19508
rect 5123 19468 5172 19496
rect 5123 19465 5135 19468
rect 5077 19459 5135 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 13354 19496 13360 19508
rect 13096 19468 13360 19496
rect 3804 19360 3832 19456
rect 3970 19388 3976 19440
rect 4028 19428 4034 19440
rect 4028 19400 4752 19428
rect 4028 19388 4034 19400
rect 4724 19369 4752 19400
rect 4065 19363 4123 19369
rect 4065 19360 4077 19363
rect 3804 19332 4077 19360
rect 4065 19329 4077 19332
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19360 4767 19363
rect 5074 19360 5080 19372
rect 4755 19332 5080 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 13096 19369 13124 19468
rect 13354 19456 13360 19468
rect 13412 19496 13418 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 13412 19468 13553 19496
rect 13412 19456 13418 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 18230 19496 18236 19508
rect 18191 19468 18236 19496
rect 13541 19459 13599 19465
rect 18230 19456 18236 19468
rect 18288 19496 18294 19508
rect 18555 19499 18613 19505
rect 18555 19496 18567 19499
rect 18288 19468 18567 19496
rect 18288 19456 18294 19468
rect 18555 19465 18567 19468
rect 18601 19465 18613 19499
rect 18966 19496 18972 19508
rect 18927 19468 18972 19496
rect 18555 19459 18613 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19518 19496 19524 19508
rect 19479 19468 19524 19496
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 13081 19363 13139 19369
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19484 19332 19717 19360
rect 19484 19320 19490 19332
rect 19705 19329 19717 19332
rect 19751 19360 19763 19363
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 19751 19332 20637 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 18484 19295 18542 19301
rect 18484 19261 18496 19295
rect 18530 19292 18542 19295
rect 18966 19292 18972 19304
rect 18530 19264 18972 19292
rect 18530 19261 18542 19264
rect 18484 19255 18542 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19426 19184 19432 19236
rect 19484 19224 19490 19236
rect 20070 19224 20076 19236
rect 19484 19196 20076 19224
rect 19484 19184 19490 19196
rect 20070 19184 20076 19196
rect 20128 19224 20134 19236
rect 20349 19227 20407 19233
rect 20349 19224 20361 19227
rect 20128 19196 20361 19224
rect 20128 19184 20134 19196
rect 20349 19193 20361 19196
rect 20395 19193 20407 19227
rect 20349 19187 20407 19193
rect 1104 19066 21436 19088
rect 1104 19014 8497 19066
rect 8549 19014 8561 19066
rect 8613 19014 8625 19066
rect 8677 19014 8689 19066
rect 8741 19014 16012 19066
rect 16064 19014 16076 19066
rect 16128 19014 16140 19066
rect 16192 19014 16204 19066
rect 16256 19014 21436 19066
rect 1104 18992 21436 19014
rect 106 18912 112 18964
rect 164 18952 170 18964
rect 2501 18955 2559 18961
rect 2501 18952 2513 18955
rect 164 18924 2513 18952
rect 164 18912 170 18924
rect 2501 18921 2513 18924
rect 2547 18921 2559 18955
rect 2501 18915 2559 18921
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 4120 18924 4200 18952
rect 4120 18912 4126 18924
rect 4172 18893 4200 18924
rect 19518 18912 19524 18964
rect 19576 18952 19582 18964
rect 20346 18952 20352 18964
rect 19576 18924 20352 18952
rect 19576 18912 19582 18924
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 4157 18887 4215 18893
rect 4157 18853 4169 18887
rect 4203 18853 4215 18887
rect 19334 18884 19340 18896
rect 19295 18856 19340 18884
rect 4157 18847 4215 18853
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 2406 18816 2412 18828
rect 2363 18788 2412 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 3844 18720 4445 18748
rect 3844 18708 3850 18720
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 19610 18748 19616 18760
rect 19571 18720 19616 18748
rect 4433 18711 4491 18717
rect 19610 18708 19616 18720
rect 19668 18708 19674 18760
rect 1104 18522 21436 18544
rect 1104 18470 4739 18522
rect 4791 18470 4803 18522
rect 4855 18470 4867 18522
rect 4919 18470 4931 18522
rect 4983 18470 12255 18522
rect 12307 18470 12319 18522
rect 12371 18470 12383 18522
rect 12435 18470 12447 18522
rect 12499 18470 19770 18522
rect 19822 18470 19834 18522
rect 19886 18470 19898 18522
rect 19950 18470 19962 18522
rect 20014 18470 21436 18522
rect 1104 18448 21436 18470
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 4157 18411 4215 18417
rect 4157 18408 4169 18411
rect 4120 18380 4169 18408
rect 4120 18368 4126 18380
rect 4157 18377 4169 18380
rect 4203 18377 4215 18411
rect 19334 18408 19340 18420
rect 19295 18380 19340 18408
rect 4157 18371 4215 18377
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 3786 18340 3792 18352
rect 3747 18312 3792 18340
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18272 3111 18275
rect 3237 18275 3295 18281
rect 3237 18272 3249 18275
rect 3099 18244 3249 18272
rect 3099 18241 3111 18244
rect 3053 18235 3111 18241
rect 3237 18241 3249 18244
rect 3283 18272 3295 18275
rect 3970 18272 3976 18284
rect 3283 18244 3976 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 3970 18232 3976 18244
rect 4028 18232 4034 18284
rect 2406 18068 2412 18080
rect 2367 18040 2412 18068
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 1104 17978 21436 18000
rect 1104 17926 8497 17978
rect 8549 17926 8561 17978
rect 8613 17926 8625 17978
rect 8677 17926 8689 17978
rect 8741 17926 16012 17978
rect 16064 17926 16076 17978
rect 16128 17926 16140 17978
rect 16192 17926 16204 17978
rect 16256 17926 21436 17978
rect 1104 17904 21436 17926
rect 2406 17824 2412 17876
rect 2464 17864 2470 17876
rect 3007 17867 3065 17873
rect 3007 17864 3019 17867
rect 2464 17836 3019 17864
rect 2464 17824 2470 17836
rect 3007 17833 3019 17836
rect 3053 17833 3065 17867
rect 3007 17827 3065 17833
rect 2958 17737 2964 17740
rect 2936 17731 2964 17737
rect 2936 17728 2948 17731
rect 2871 17700 2948 17728
rect 2936 17697 2948 17700
rect 3016 17728 3022 17740
rect 3786 17728 3792 17740
rect 3016 17700 3792 17728
rect 2936 17691 2964 17697
rect 2958 17688 2964 17691
rect 3016 17688 3022 17700
rect 3786 17688 3792 17700
rect 3844 17688 3850 17740
rect 7628 17731 7686 17737
rect 7628 17697 7640 17731
rect 7674 17728 7686 17731
rect 8386 17728 8392 17740
rect 7674 17700 8392 17728
rect 7674 17697 7686 17700
rect 7628 17691 7686 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 7699 17527 7757 17533
rect 7699 17524 7711 17527
rect 7432 17496 7711 17524
rect 7432 17484 7438 17496
rect 7699 17493 7711 17496
rect 7745 17493 7757 17527
rect 7699 17487 7757 17493
rect 1104 17434 21436 17456
rect 1104 17382 4739 17434
rect 4791 17382 4803 17434
rect 4855 17382 4867 17434
rect 4919 17382 4931 17434
rect 4983 17382 12255 17434
rect 12307 17382 12319 17434
rect 12371 17382 12383 17434
rect 12435 17382 12447 17434
rect 12499 17382 19770 17434
rect 19822 17382 19834 17434
rect 19886 17382 19898 17434
rect 19950 17382 19962 17434
rect 20014 17382 21436 17434
rect 1104 17360 21436 17382
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 7374 17184 7380 17196
rect 7239 17156 7380 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 7650 17184 7656 17196
rect 7611 17156 7656 17184
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8386 17184 8392 17196
rect 8347 17156 8392 17184
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 2774 17076 2780 17128
rect 2832 17116 2838 17128
rect 4062 17116 4068 17128
rect 2832 17088 4068 17116
rect 2832 17076 2838 17088
rect 4062 17076 4068 17088
rect 4120 17116 4126 17128
rect 5144 17119 5202 17125
rect 5144 17116 5156 17119
rect 4120 17088 5156 17116
rect 4120 17076 4126 17088
rect 5144 17085 5156 17088
rect 5190 17116 5202 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5190 17088 5549 17116
rect 5190 17085 5202 17088
rect 5144 17079 5202 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 5215 16983 5273 16989
rect 5215 16949 5227 16983
rect 5261 16980 5273 16983
rect 6086 16980 6092 16992
rect 5261 16952 6092 16980
rect 5261 16949 5273 16952
rect 5215 16943 5273 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 1104 16890 21436 16912
rect 1104 16838 8497 16890
rect 8549 16838 8561 16890
rect 8613 16838 8625 16890
rect 8677 16838 8689 16890
rect 8741 16838 16012 16890
rect 16064 16838 16076 16890
rect 16128 16838 16140 16890
rect 16192 16838 16204 16890
rect 16256 16838 21436 16890
rect 1104 16816 21436 16838
rect 6086 16708 6092 16720
rect 6047 16680 6092 16708
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 6733 16711 6791 16717
rect 6733 16677 6745 16711
rect 6779 16708 6791 16711
rect 7650 16708 7656 16720
rect 6779 16680 7656 16708
rect 6779 16677 6791 16680
rect 6733 16671 6791 16677
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4430 16640 4436 16652
rect 4488 16649 4494 16652
rect 4488 16643 4526 16649
rect 4120 16612 4436 16640
rect 4120 16600 4126 16612
rect 4430 16600 4436 16612
rect 4514 16609 4526 16643
rect 4488 16603 4526 16609
rect 11032 16643 11090 16649
rect 11032 16609 11044 16643
rect 11078 16640 11090 16643
rect 11146 16640 11152 16652
rect 11078 16612 11152 16640
rect 11078 16609 11090 16612
rect 11032 16603 11090 16609
rect 4488 16600 4494 16603
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 4614 16445 4620 16448
rect 4571 16439 4620 16445
rect 4571 16436 4583 16439
rect 4527 16408 4583 16436
rect 4571 16405 4583 16408
rect 4617 16405 4620 16439
rect 4571 16399 4620 16405
rect 4614 16396 4620 16399
rect 4672 16436 4678 16448
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4672 16408 4905 16436
rect 4672 16396 4678 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 11103 16439 11161 16445
rect 11103 16405 11115 16439
rect 11149 16436 11161 16439
rect 11974 16436 11980 16448
rect 11149 16408 11980 16436
rect 11149 16405 11161 16408
rect 11103 16399 11161 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 1104 16346 21436 16368
rect 1104 16294 4739 16346
rect 4791 16294 4803 16346
rect 4855 16294 4867 16346
rect 4919 16294 4931 16346
rect 4983 16294 12255 16346
rect 12307 16294 12319 16346
rect 12371 16294 12383 16346
rect 12435 16294 12447 16346
rect 12499 16294 19770 16346
rect 19822 16294 19834 16346
rect 19886 16294 19898 16346
rect 19950 16294 19962 16346
rect 20014 16294 21436 16346
rect 1104 16272 21436 16294
rect 4430 16232 4436 16244
rect 4391 16204 4436 16232
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 6086 16232 6092 16244
rect 6047 16204 6092 16232
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11204 16204 11345 16232
rect 11204 16192 11210 16204
rect 11333 16201 11345 16204
rect 11379 16232 11391 16235
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11379 16204 11713 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 11701 16195 11759 16201
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 4672 16068 4905 16096
rect 4672 16056 4678 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 10940 16031 10998 16037
rect 10940 15997 10952 16031
rect 10986 16028 10998 16031
rect 11146 16028 11152 16040
rect 10986 16000 11152 16028
rect 10986 15997 10998 16000
rect 10940 15991 10998 15997
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 5534 15960 5540 15972
rect 5495 15932 5540 15960
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 11011 15895 11069 15901
rect 11011 15861 11023 15895
rect 11057 15892 11069 15895
rect 11238 15892 11244 15904
rect 11057 15864 11244 15892
rect 11057 15861 11069 15864
rect 11011 15855 11069 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 1104 15802 21436 15824
rect 1104 15750 8497 15802
rect 8549 15750 8561 15802
rect 8613 15750 8625 15802
rect 8677 15750 8689 15802
rect 8741 15750 16012 15802
rect 16064 15750 16076 15802
rect 16128 15750 16140 15802
rect 16192 15750 16204 15802
rect 16256 15750 21436 15802
rect 1104 15728 21436 15750
rect 15470 15688 15476 15700
rect 15431 15660 15476 15688
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 5534 15620 5540 15632
rect 5495 15592 5540 15620
rect 5534 15580 5540 15592
rect 5592 15620 5598 15632
rect 6457 15623 6515 15629
rect 6457 15620 6469 15623
rect 5592 15592 6469 15620
rect 5592 15580 5598 15592
rect 6457 15589 6469 15592
rect 6503 15589 6515 15623
rect 6457 15583 6515 15589
rect 11238 15580 11244 15632
rect 11296 15620 11302 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11296 15592 11529 15620
rect 11296 15580 11302 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 11517 15583 11575 15589
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 10448 15555 10506 15561
rect 10448 15552 10460 15555
rect 9916 15524 10460 15552
rect 9916 15512 9922 15524
rect 10448 15521 10460 15524
rect 10494 15521 10506 15555
rect 10448 15515 10506 15521
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 14220 15555 14278 15561
rect 14220 15552 14232 15555
rect 12952 15524 14232 15552
rect 12952 15512 12958 15524
rect 14220 15521 14232 15524
rect 14266 15552 14278 15555
rect 14458 15552 14464 15564
rect 14266 15524 14464 15552
rect 14266 15521 14278 15524
rect 14220 15515 14278 15521
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15484 4951 15487
rect 5074 15484 5080 15496
rect 4939 15456 5080 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 3878 15376 3884 15428
rect 3936 15416 3942 15428
rect 7009 15419 7067 15425
rect 7009 15416 7021 15419
rect 3936 15388 4154 15416
rect 3936 15376 3942 15388
rect 4126 15348 4154 15388
rect 6104 15388 7021 15416
rect 6104 15348 6132 15388
rect 7009 15385 7021 15388
rect 7055 15385 7067 15419
rect 12066 15416 12072 15428
rect 12027 15388 12072 15416
rect 7009 15379 7067 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 4126 15320 6132 15348
rect 10551 15351 10609 15357
rect 10551 15317 10563 15351
rect 10597 15348 10609 15351
rect 11422 15348 11428 15360
rect 10597 15320 11428 15348
rect 10597 15317 10609 15320
rect 10551 15311 10609 15317
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 14323 15351 14381 15357
rect 14323 15317 14335 15351
rect 14369 15348 14381 15351
rect 15470 15348 15476 15360
rect 14369 15320 15476 15348
rect 14369 15317 14381 15320
rect 14323 15311 14381 15317
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 1104 15258 21436 15280
rect 1104 15206 4739 15258
rect 4791 15206 4803 15258
rect 4855 15206 4867 15258
rect 4919 15206 4931 15258
rect 4983 15206 12255 15258
rect 12307 15206 12319 15258
rect 12371 15206 12383 15258
rect 12435 15206 12447 15258
rect 12499 15206 19770 15258
rect 19822 15206 19834 15258
rect 19886 15206 19898 15258
rect 19950 15206 19962 15258
rect 20014 15206 21436 15258
rect 1104 15184 21436 15206
rect 4295 15147 4353 15153
rect 4295 15113 4307 15147
rect 4341 15144 4353 15147
rect 5074 15144 5080 15156
rect 4341 15116 5080 15144
rect 4341 15113 4353 15116
rect 4295 15107 4353 15113
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 9858 15144 9864 15156
rect 9723 15116 9864 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 9835 15104 9864 15116
rect 9916 15144 9922 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 9916 15116 10425 15144
rect 9916 15104 9922 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11296 15116 11805 15144
rect 11296 15104 11302 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 12032 15116 12173 15144
rect 12032 15104 12038 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 12161 15107 12219 15113
rect 5534 15008 5540 15020
rect 5495 14980 5540 15008
rect 5534 14968 5540 14980
rect 5592 15008 5598 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5592 14980 6377 15008
rect 5592 14968 5598 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 4224 14943 4282 14949
rect 4224 14909 4236 14943
rect 4270 14940 4282 14943
rect 4614 14940 4620 14952
rect 4270 14912 4620 14940
rect 4270 14909 4282 14912
rect 4224 14903 4282 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5902 14900 5908 14952
rect 5960 14940 5966 14952
rect 6892 14943 6950 14949
rect 6892 14940 6904 14943
rect 5960 14912 6904 14940
rect 5960 14900 5966 14912
rect 6892 14909 6904 14912
rect 6938 14940 6950 14943
rect 7374 14940 7380 14952
rect 6938 14912 7380 14940
rect 6938 14909 6950 14912
rect 6892 14903 6950 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 9835 14949 9863 15104
rect 12176 15008 12204 15107
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 15151 15079 15209 15085
rect 15151 15045 15163 15079
rect 15197 15076 15209 15079
rect 15286 15076 15292 15088
rect 15197 15048 15292 15076
rect 15197 15045 15209 15048
rect 15151 15039 15209 15045
rect 15286 15036 15292 15048
rect 15344 15076 15350 15088
rect 15841 15079 15899 15085
rect 15841 15076 15853 15079
rect 15344 15048 15853 15076
rect 15344 15036 15350 15048
rect 15841 15045 15853 15048
rect 15887 15045 15899 15079
rect 15841 15039 15899 15045
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 12176 14980 12541 15008
rect 12529 14977 12541 14980
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 9820 14943 9878 14949
rect 9820 14909 9832 14943
rect 9866 14909 9878 14943
rect 9820 14903 9878 14909
rect 14068 14943 14126 14949
rect 14068 14909 14080 14943
rect 14114 14940 14126 14943
rect 14458 14940 14464 14952
rect 14114 14912 14464 14940
rect 14114 14909 14126 14912
rect 14068 14903 14126 14909
rect 14458 14900 14464 14912
rect 14516 14940 14522 14952
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14516 14912 14841 14940
rect 14516 14900 14522 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 15080 14943 15138 14949
rect 15080 14909 15092 14943
rect 15126 14940 15138 14943
rect 15126 14912 15424 14940
rect 15126 14909 15138 14912
rect 15080 14903 15138 14909
rect 5258 14872 5264 14884
rect 5219 14844 5264 14872
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 9907 14875 9965 14881
rect 9907 14841 9919 14875
rect 9953 14872 9965 14875
rect 10870 14872 10876 14884
rect 9953 14844 10876 14872
rect 9953 14841 9965 14844
rect 9907 14835 9965 14841
rect 10870 14832 10876 14844
rect 10928 14832 10934 14884
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14872 11575 14875
rect 12986 14872 12992 14884
rect 11563 14844 12992 14872
rect 11563 14841 11575 14844
rect 11517 14835 11575 14841
rect 12986 14832 12992 14844
rect 13044 14872 13050 14884
rect 13173 14875 13231 14881
rect 13173 14872 13185 14875
rect 13044 14844 13185 14872
rect 13044 14832 13050 14844
rect 13173 14841 13185 14844
rect 13219 14841 13231 14875
rect 13173 14835 13231 14841
rect 15396 14816 15424 14912
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 17012 14943 17070 14949
rect 17012 14940 17024 14943
rect 16908 14912 17024 14940
rect 16908 14900 16914 14912
rect 17012 14909 17024 14912
rect 17058 14940 17070 14943
rect 17494 14940 17500 14952
rect 17058 14912 17500 14940
rect 17058 14909 17070 14912
rect 17012 14903 17070 14909
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 6963 14807 7021 14813
rect 6963 14804 6975 14807
rect 6880 14776 6975 14804
rect 6880 14764 6886 14776
rect 6963 14773 6975 14776
rect 7009 14773 7021 14807
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 6963 14767 7021 14773
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 13998 14764 14004 14816
rect 14056 14804 14062 14816
rect 14139 14807 14197 14813
rect 14139 14804 14151 14807
rect 14056 14776 14151 14804
rect 14056 14764 14062 14776
rect 14139 14773 14151 14776
rect 14185 14773 14197 14807
rect 14139 14767 14197 14773
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15473 14807 15531 14813
rect 15473 14804 15485 14807
rect 15436 14776 15485 14804
rect 15436 14764 15442 14776
rect 15473 14773 15485 14776
rect 15519 14773 15531 14807
rect 15473 14767 15531 14773
rect 17083 14807 17141 14813
rect 17083 14773 17095 14807
rect 17129 14804 17141 14807
rect 17218 14804 17224 14816
rect 17129 14776 17224 14804
rect 17129 14773 17141 14776
rect 17083 14767 17141 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 1104 14714 21436 14736
rect 1104 14662 8497 14714
rect 8549 14662 8561 14714
rect 8613 14662 8625 14714
rect 8677 14662 8689 14714
rect 8741 14662 16012 14714
rect 16064 14662 16076 14714
rect 16128 14662 16140 14714
rect 16192 14662 16204 14714
rect 16256 14662 21436 14714
rect 1104 14640 21436 14662
rect 5258 14600 5264 14612
rect 5219 14572 5264 14600
rect 5258 14560 5264 14572
rect 5316 14600 5322 14612
rect 5859 14603 5917 14609
rect 5859 14600 5871 14603
rect 5316 14572 5871 14600
rect 5316 14560 5322 14572
rect 5859 14569 5871 14572
rect 5905 14569 5917 14603
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 5859 14563 5917 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 6822 14532 6828 14544
rect 6783 14504 6828 14532
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 7469 14535 7527 14541
rect 7469 14501 7481 14535
rect 7515 14532 7527 14535
rect 7650 14532 7656 14544
rect 7515 14504 7656 14532
rect 7515 14501 7527 14504
rect 7469 14495 7527 14501
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 11422 14532 11428 14544
rect 11383 14504 11428 14532
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 12066 14532 12072 14544
rect 12027 14504 12072 14532
rect 12066 14492 12072 14504
rect 12124 14492 12130 14544
rect 12986 14532 12992 14544
rect 12947 14504 12992 14532
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 15470 14532 15476 14544
rect 15431 14504 15476 14532
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 17218 14532 17224 14544
rect 17179 14504 17224 14532
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 1464 14467 1522 14473
rect 1464 14433 1476 14467
rect 1510 14464 1522 14467
rect 1946 14464 1952 14476
rect 1510 14436 1952 14464
rect 1510 14433 1522 14436
rect 1464 14427 1522 14433
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4744 14467 4802 14473
rect 4744 14464 4756 14467
rect 4672 14436 4756 14464
rect 4672 14424 4678 14436
rect 4744 14433 4756 14436
rect 4790 14433 4802 14467
rect 4744 14427 4802 14433
rect 5788 14467 5846 14473
rect 5788 14433 5800 14467
rect 5834 14464 5846 14467
rect 5902 14464 5908 14476
rect 5834 14436 5908 14464
rect 5834 14433 5846 14436
rect 5788 14427 5846 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 9712 14467 9770 14473
rect 9712 14464 9724 14467
rect 9364 14436 9724 14464
rect 9364 14424 9370 14436
rect 9712 14433 9724 14436
rect 9758 14433 9770 14467
rect 9712 14427 9770 14433
rect 13262 14396 13268 14408
rect 13223 14368 13268 14396
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14396 17923 14399
rect 17954 14396 17960 14408
rect 17911 14368 17960 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 17954 14356 17960 14368
rect 18012 14356 18018 14408
rect 4847 14331 4905 14337
rect 4847 14297 4859 14331
rect 4893 14328 4905 14331
rect 5442 14328 5448 14340
rect 4893 14300 5448 14328
rect 4893 14297 4905 14300
rect 4847 14291 4905 14297
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14328 16083 14331
rect 17126 14328 17132 14340
rect 16071 14300 17132 14328
rect 16071 14297 16083 14300
rect 16025 14291 16083 14297
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1535 14263 1593 14269
rect 1535 14260 1547 14263
rect 1452 14232 1547 14260
rect 1452 14220 1458 14232
rect 1535 14229 1547 14232
rect 1581 14229 1593 14263
rect 1535 14223 1593 14229
rect 9815 14263 9873 14269
rect 9815 14229 9827 14263
rect 9861 14260 9873 14263
rect 10134 14260 10140 14272
rect 9861 14232 10140 14260
rect 9861 14229 9873 14232
rect 9815 14223 9873 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 1104 14170 21436 14192
rect 1104 14118 4739 14170
rect 4791 14118 4803 14170
rect 4855 14118 4867 14170
rect 4919 14118 4931 14170
rect 4983 14118 12255 14170
rect 12307 14118 12319 14170
rect 12371 14118 12383 14170
rect 12435 14118 12447 14170
rect 12499 14118 19770 14170
rect 19822 14118 19834 14170
rect 19886 14118 19898 14170
rect 19950 14118 19962 14170
rect 20014 14118 21436 14170
rect 1104 14096 21436 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4614 14056 4620 14068
rect 4571 14028 4620 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 5902 14056 5908 14068
rect 5859 14028 5908 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 6822 14056 6828 14068
rect 6687 14028 6828 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 10134 14056 10140 14068
rect 10095 14028 10140 14056
rect 10134 14016 10140 14028
rect 10192 14056 10198 14068
rect 11422 14056 11428 14068
rect 10192 14028 10456 14056
rect 11383 14028 11428 14056
rect 10192 14016 10198 14028
rect 6273 13991 6331 13997
rect 6273 13957 6285 13991
rect 6319 13988 6331 13991
rect 7650 13988 7656 14000
rect 6319 13960 7656 13988
rect 6319 13957 6331 13960
rect 6273 13951 6331 13957
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4338 13920 4344 13932
rect 3936 13892 4344 13920
rect 3936 13880 3942 13892
rect 4338 13880 4344 13892
rect 4396 13920 4402 13932
rect 7116 13929 7144 13960
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 9398 13988 9404 14000
rect 9359 13960 9404 13988
rect 9398 13948 9404 13960
rect 9456 13988 9462 14000
rect 9674 13988 9680 14000
rect 9456 13960 9680 13988
rect 9456 13948 9462 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 10428 13929 10456 14028
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 13998 14016 14004 14028
rect 14056 14056 14062 14068
rect 15470 14056 15476 14068
rect 14056 14028 14228 14056
rect 15431 14028 15476 14056
rect 14056 14016 14062 14028
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 11011 13960 14044 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 4985 13923 5043 13929
rect 4985 13920 4997 13923
rect 4396 13892 4997 13920
rect 4396 13880 4402 13892
rect 4985 13889 4997 13892
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 7101 13923 7159 13929
rect 7101 13889 7113 13923
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 10413 13923 10471 13929
rect 10413 13889 10425 13923
rect 10459 13889 10471 13923
rect 12986 13920 12992 13932
rect 12947 13892 12992 13920
rect 10413 13883 10471 13889
rect 12986 13880 12992 13892
rect 13044 13920 13050 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13044 13892 13553 13920
rect 13044 13880 13050 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13852 1458 13864
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 1452 13824 2329 13852
rect 1452 13812 1458 13824
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 3640 13855 3698 13861
rect 3640 13852 3652 13855
rect 3568 13824 3652 13852
rect 3568 13812 3574 13824
rect 3640 13821 3652 13824
rect 3686 13852 3698 13855
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 3686 13824 4077 13852
rect 3686 13821 3698 13824
rect 3640 13815 3698 13821
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 3743 13787 3801 13793
rect 3743 13753 3755 13787
rect 3789 13784 3801 13787
rect 4522 13784 4528 13796
rect 3789 13756 4528 13784
rect 3789 13753 3801 13756
rect 3743 13747 3801 13753
rect 4522 13744 4528 13756
rect 4580 13744 4586 13796
rect 4706 13784 4712 13796
rect 4667 13756 4712 13784
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 7742 13784 7748 13796
rect 7703 13756 7748 13784
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 8588 13756 8861 13784
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8588 13725 8616 13756
rect 8849 13753 8861 13756
rect 8895 13753 8907 13787
rect 8849 13747 8907 13753
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 12253 13787 12311 13793
rect 9732 13756 10134 13784
rect 9732 13744 9738 13756
rect 8573 13719 8631 13725
rect 8573 13716 8585 13719
rect 8444 13688 8585 13716
rect 8444 13676 8450 13688
rect 8573 13685 8585 13688
rect 8619 13685 8631 13719
rect 8573 13679 8631 13685
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 9769 13719 9827 13725
rect 9769 13716 9781 13719
rect 9456 13688 9781 13716
rect 9456 13676 9462 13688
rect 9769 13685 9781 13688
rect 9815 13685 9827 13719
rect 10106 13716 10134 13756
rect 12253 13753 12265 13787
rect 12299 13784 12311 13787
rect 12621 13787 12679 13793
rect 12621 13784 12633 13787
rect 12299 13756 12633 13784
rect 12299 13753 12311 13756
rect 12253 13747 12311 13753
rect 12621 13753 12633 13756
rect 12667 13784 12679 13787
rect 13906 13784 13912 13796
rect 12667 13756 13912 13784
rect 12667 13753 12679 13756
rect 12621 13747 12679 13753
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 14016 13784 14044 13960
rect 14200 13929 14228 14028
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 17276 14028 17417 14056
rect 17276 14016 17282 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 17954 13920 17960 13932
rect 16264 13892 17960 13920
rect 16264 13880 16270 13892
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 14829 13787 14887 13793
rect 14829 13784 14841 13787
rect 14016 13756 14841 13784
rect 14829 13753 14841 13756
rect 14875 13784 14887 13787
rect 16206 13784 16212 13796
rect 14875 13756 16212 13784
rect 14875 13753 14887 13756
rect 14829 13747 14887 13753
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 16301 13787 16359 13793
rect 16301 13753 16313 13787
rect 16347 13784 16359 13787
rect 16482 13784 16488 13796
rect 16347 13756 16488 13784
rect 16347 13753 16359 13756
rect 16301 13747 16359 13753
rect 16482 13744 16488 13756
rect 16540 13744 16546 13796
rect 17126 13784 17132 13796
rect 17087 13756 17132 13784
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 13262 13716 13268 13728
rect 10106 13688 13268 13716
rect 9769 13679 9827 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 1104 13626 21436 13648
rect 1104 13574 8497 13626
rect 8549 13574 8561 13626
rect 8613 13574 8625 13626
rect 8677 13574 8689 13626
rect 8741 13574 16012 13626
rect 16064 13574 16076 13626
rect 16128 13574 16140 13626
rect 16192 13574 16204 13626
rect 16256 13574 21436 13626
rect 1104 13552 21436 13574
rect 4246 13512 4252 13524
rect 4207 13484 4252 13512
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 4706 13512 4712 13524
rect 4667 13484 4712 13512
rect 4706 13472 4712 13484
rect 4764 13512 4770 13524
rect 5074 13512 5080 13524
rect 4764 13484 5080 13512
rect 4764 13472 4770 13484
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13814 13512 13820 13524
rect 13587 13484 13820 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 15427 13515 15485 13521
rect 15427 13512 15439 13515
rect 13964 13484 15439 13512
rect 13964 13472 13970 13484
rect 15427 13481 15439 13484
rect 15473 13481 15485 13515
rect 15427 13475 15485 13481
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16899 13515 16957 13521
rect 16899 13512 16911 13515
rect 16540 13484 16911 13512
rect 16540 13472 16546 13484
rect 16899 13481 16911 13484
rect 16945 13481 16957 13515
rect 16899 13475 16957 13481
rect 17954 13444 17960 13456
rect 17915 13416 17960 13444
rect 17954 13404 17960 13416
rect 18012 13404 18018 13456
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13376 2467 13379
rect 2498 13376 2504 13388
rect 2455 13348 2504 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13044 13348 13369 13376
rect 13044 13336 13050 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 15356 13379 15414 13385
rect 15356 13345 15368 13379
rect 15402 13376 15414 13379
rect 15470 13376 15476 13388
rect 15402 13348 15476 13376
rect 15402 13345 15414 13348
rect 15356 13339 15414 13345
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 16850 13376 16856 13388
rect 16715 13348 16856 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 5442 13308 5448 13320
rect 5403 13280 5448 13308
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6135 13280 7021 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 7009 13277 7021 13280
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 7742 13308 7748 13320
rect 7699 13280 7748 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10045 13311 10103 13317
rect 10045 13277 10057 13311
rect 10091 13277 10103 13311
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 10045 13271 10103 13277
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 10060 13240 10088 13271
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 18598 13308 18604 13320
rect 18559 13280 18604 13308
rect 11977 13271 12035 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 8444 13212 10088 13240
rect 8444 13200 8450 13212
rect 2547 13175 2605 13181
rect 2547 13141 2559 13175
rect 2593 13172 2605 13175
rect 3326 13172 3332 13184
rect 2593 13144 3332 13172
rect 2593 13141 2605 13144
rect 2547 13135 2605 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 1104 13082 21436 13104
rect 1104 13030 4739 13082
rect 4791 13030 4803 13082
rect 4855 13030 4867 13082
rect 4919 13030 4931 13082
rect 4983 13030 12255 13082
rect 12307 13030 12319 13082
rect 12371 13030 12383 13082
rect 12435 13030 12447 13082
rect 12499 13030 19770 13082
rect 19822 13030 19834 13082
rect 19886 13030 19898 13082
rect 19950 13030 19962 13082
rect 20014 13030 21436 13082
rect 1104 13008 21436 13030
rect 4338 12968 4344 12980
rect 4299 12940 4344 12968
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4580 12940 4997 12968
rect 4580 12928 4586 12940
rect 4985 12937 4997 12940
rect 5031 12968 5043 12971
rect 5031 12940 5304 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 3927 12903 3985 12909
rect 3927 12869 3939 12903
rect 3973 12900 3985 12903
rect 4062 12900 4068 12912
rect 3973 12872 4068 12900
rect 3973 12869 3985 12872
rect 3927 12863 3985 12869
rect 4062 12860 4068 12872
rect 4120 12900 4126 12912
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4120 12872 4629 12900
rect 4120 12860 4126 12872
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 5276 12841 5304 12940
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5500 12940 6193 12968
rect 5500 12928 5506 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 9766 12968 9772 12980
rect 9727 12940 9772 12968
rect 6181 12931 6239 12937
rect 9766 12928 9772 12940
rect 9824 12968 9830 12980
rect 10091 12971 10149 12977
rect 10091 12968 10103 12971
rect 9824 12940 10103 12968
rect 9824 12928 9830 12940
rect 10091 12937 10103 12940
rect 10137 12937 10149 12971
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 10091 12931 10149 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17865 12971 17923 12977
rect 17865 12937 17877 12971
rect 17911 12968 17923 12971
rect 17954 12968 17960 12980
rect 17911 12940 17960 12968
rect 17911 12937 17923 12940
rect 17865 12931 17923 12937
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 21082 12968 21088 12980
rect 20027 12940 21088 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11291 12872 11805 12900
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7098 12832 7104 12844
rect 6687 12804 7104 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7098 12792 7104 12804
rect 7156 12832 7162 12844
rect 7558 12832 7564 12844
rect 7156 12804 7564 12832
rect 7156 12792 7162 12804
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 106 12724 112 12776
rect 164 12764 170 12776
rect 1432 12767 1490 12773
rect 1432 12764 1444 12767
rect 164 12736 1444 12764
rect 164 12724 170 12736
rect 1432 12733 1444 12736
rect 1478 12764 1490 12767
rect 1857 12767 1915 12773
rect 1857 12764 1869 12767
rect 1478 12736 1869 12764
rect 1478 12733 1490 12736
rect 1432 12727 1490 12733
rect 1857 12733 1869 12736
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 3856 12767 3914 12773
rect 3856 12733 3868 12767
rect 3902 12764 3914 12767
rect 4338 12764 4344 12776
rect 3902 12736 4344 12764
rect 3902 12733 3914 12736
rect 3856 12727 3914 12733
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 9008 12767 9066 12773
rect 9008 12733 9020 12767
rect 9054 12764 9066 12767
rect 9398 12764 9404 12776
rect 9054 12736 9404 12764
rect 9054 12733 9066 12736
rect 9008 12727 9066 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 11291 12773 11319 12872
rect 11793 12869 11805 12872
rect 11839 12900 11851 12903
rect 22094 12900 22100 12912
rect 11839 12872 22100 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 11379 12835 11437 12841
rect 11379 12801 11391 12835
rect 11425 12832 11437 12835
rect 11698 12832 11704 12844
rect 11425 12804 11704 12832
rect 11425 12801 11437 12804
rect 11379 12795 11437 12801
rect 11698 12792 11704 12804
rect 11756 12832 11762 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11756 12804 12081 12832
rect 11756 12792 11762 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 14182 12832 14188 12844
rect 14095 12804 14188 12832
rect 12069 12795 12127 12801
rect 14182 12792 14188 12804
rect 14240 12832 14246 12844
rect 15378 12832 15384 12844
rect 14240 12804 15384 12832
rect 14240 12792 14246 12804
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 10020 12767 10078 12773
rect 10020 12733 10032 12767
rect 10066 12764 10078 12767
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10066 12736 10517 12764
rect 10066 12733 10078 12736
rect 10020 12727 10078 12733
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 11276 12767 11334 12773
rect 11276 12764 11288 12767
rect 10551 12736 11288 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 11276 12733 11288 12736
rect 11322 12733 11334 12767
rect 11276 12727 11334 12733
rect 19610 12724 19616 12776
rect 19668 12764 19674 12776
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19668 12736 19809 12764
rect 19668 12724 19674 12736
rect 19797 12733 19809 12736
rect 19843 12764 19855 12767
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 19843 12736 20361 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 2777 12699 2835 12705
rect 2777 12665 2789 12699
rect 2823 12696 2835 12699
rect 5905 12699 5963 12705
rect 2823 12668 4154 12696
rect 2823 12665 2835 12668
rect 2777 12659 2835 12665
rect 4126 12640 4154 12668
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 7098 12696 7104 12708
rect 5951 12668 7104 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 7742 12696 7748 12708
rect 7655 12668 7748 12696
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8202 12696 8208 12708
rect 7800 12668 8208 12696
rect 7800 12656 7806 12668
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 12437 12699 12495 12705
rect 12437 12665 12449 12699
rect 12483 12696 12495 12699
rect 13265 12699 13323 12705
rect 13265 12696 13277 12699
rect 12483 12668 13277 12696
rect 12483 12665 12495 12668
rect 12437 12659 12495 12665
rect 13265 12665 13277 12668
rect 13311 12696 13323 12699
rect 13541 12699 13599 12705
rect 13541 12696 13553 12699
rect 13311 12668 13553 12696
rect 13311 12665 13323 12668
rect 13265 12659 13323 12665
rect 13541 12665 13553 12668
rect 13587 12665 13599 12699
rect 13541 12659 13599 12665
rect 17497 12699 17555 12705
rect 17497 12665 17509 12699
rect 17543 12696 17555 12699
rect 18325 12699 18383 12705
rect 18325 12696 18337 12699
rect 17543 12668 18337 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 18325 12665 18337 12668
rect 18371 12696 18383 12699
rect 18414 12696 18420 12708
rect 18371 12668 18420 12696
rect 18371 12665 18383 12668
rect 18325 12659 18383 12665
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 1535 12631 1593 12637
rect 1535 12597 1547 12631
rect 1581 12628 1593 12631
rect 2222 12628 2228 12640
rect 1581 12600 2228 12628
rect 1581 12597 1593 12600
rect 1535 12591 1593 12597
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 4126 12600 4160 12640
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 7116 12628 7144 12656
rect 7834 12628 7840 12640
rect 7116 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12628 7898 12640
rect 8021 12631 8079 12637
rect 8021 12628 8033 12631
rect 7892 12600 8033 12628
rect 7892 12588 7898 12600
rect 8021 12597 8033 12600
rect 8067 12597 8079 12631
rect 8021 12591 8079 12597
rect 9079 12631 9137 12637
rect 9079 12597 9091 12631
rect 9125 12628 9137 12631
rect 9306 12628 9312 12640
rect 9125 12600 9312 12628
rect 9125 12597 9137 12600
rect 9079 12591 9137 12597
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 15470 12628 15476 12640
rect 15427 12600 15476 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15470 12588 15476 12600
rect 15528 12628 15534 12640
rect 18046 12628 18052 12640
rect 15528 12600 18052 12628
rect 15528 12588 15534 12600
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 1104 12538 21436 12560
rect 1104 12486 8497 12538
rect 8549 12486 8561 12538
rect 8613 12486 8625 12538
rect 8677 12486 8689 12538
rect 8741 12486 16012 12538
rect 16064 12486 16076 12538
rect 16128 12486 16140 12538
rect 16192 12486 16204 12538
rect 16256 12486 21436 12538
rect 1104 12464 21436 12486
rect 1394 12316 1400 12368
rect 1452 12356 1458 12368
rect 1581 12359 1639 12365
rect 1581 12356 1593 12359
rect 1452 12328 1593 12356
rect 1452 12316 1458 12328
rect 1581 12325 1593 12328
rect 1627 12325 1639 12359
rect 1581 12319 1639 12325
rect 9306 12316 9312 12368
rect 9364 12356 9370 12368
rect 9766 12356 9772 12368
rect 9364 12328 9772 12356
rect 9364 12316 9370 12328
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 11882 12316 11888 12368
rect 11940 12356 11946 12368
rect 12894 12356 12900 12368
rect 11940 12328 12900 12356
rect 11940 12316 11946 12328
rect 12894 12316 12900 12328
rect 12952 12316 12958 12368
rect 8113 12291 8171 12297
rect 8113 12257 8125 12291
rect 8159 12288 8171 12291
rect 8202 12288 8208 12300
rect 8159 12260 8208 12288
rect 8159 12257 8171 12260
rect 8113 12251 8171 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 19864 12291 19922 12297
rect 19864 12257 19876 12291
rect 19910 12288 19922 12291
rect 20714 12288 20720 12300
rect 19910 12260 20720 12288
rect 19910 12257 19922 12260
rect 19864 12251 19922 12257
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 4614 12220 4620 12232
rect 4575 12192 4620 12220
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5074 12220 5080 12232
rect 5035 12192 5080 12220
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 6638 12220 6644 12232
rect 6599 12192 6644 12220
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7098 12220 7104 12232
rect 7059 12192 7104 12220
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13630 12220 13636 12232
rect 13587 12192 13636 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 18322 12220 18328 12232
rect 18283 12192 18328 12220
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 18598 12220 18604 12232
rect 18559 12192 18604 12220
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8251 12087 8309 12093
rect 8251 12084 8263 12087
rect 7156 12056 8263 12084
rect 7156 12044 7162 12056
rect 8251 12053 8263 12056
rect 8297 12053 8309 12087
rect 8251 12047 8309 12053
rect 19935 12087 19993 12093
rect 19935 12053 19947 12087
rect 19981 12084 19993 12087
rect 20070 12084 20076 12096
rect 19981 12056 20076 12084
rect 19981 12053 19993 12056
rect 19935 12047 19993 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 1104 11994 21436 12016
rect 1104 11942 4739 11994
rect 4791 11942 4803 11994
rect 4855 11942 4867 11994
rect 4919 11942 4931 11994
rect 4983 11942 12255 11994
rect 12307 11942 12319 11994
rect 12371 11942 12383 11994
rect 12435 11942 12447 11994
rect 12499 11942 19770 11994
rect 19822 11942 19834 11994
rect 19886 11942 19898 11994
rect 19950 11942 19962 11994
rect 20014 11942 21436 11994
rect 1104 11920 21436 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1452 11852 1593 11880
rect 1452 11840 1458 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 3467 11883 3525 11889
rect 3467 11849 3479 11883
rect 3513 11880 3525 11883
rect 4614 11880 4620 11892
rect 3513 11852 4620 11880
rect 3513 11849 3525 11852
rect 3467 11843 3525 11849
rect 4614 11840 4620 11852
rect 4672 11880 4678 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 4672 11852 5365 11880
rect 4672 11840 4678 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 5353 11843 5411 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9766 11880 9772 11892
rect 9727 11852 9772 11880
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 14507 11883 14565 11889
rect 14507 11880 14519 11883
rect 13044 11852 14519 11880
rect 13044 11840 13050 11852
rect 14507 11849 14519 11852
rect 14553 11849 14565 11883
rect 14507 11843 14565 11849
rect 18555 11883 18613 11889
rect 18555 11849 18567 11883
rect 18601 11880 18613 11883
rect 19610 11880 19616 11892
rect 18601 11852 19616 11880
rect 18601 11849 18613 11852
rect 18555 11843 18613 11849
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 7834 11812 7840 11824
rect 4212 11784 4257 11812
rect 7795 11784 7840 11812
rect 4212 11772 4218 11784
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 18322 11812 18328 11824
rect 18235 11784 18328 11812
rect 18322 11772 18328 11784
rect 18380 11812 18386 11824
rect 20254 11812 20260 11824
rect 18380 11784 20260 11812
rect 18380 11772 18386 11784
rect 20254 11772 20260 11784
rect 20312 11772 20318 11824
rect 1946 11704 1952 11756
rect 2004 11744 2010 11756
rect 2133 11747 2191 11753
rect 2133 11744 2145 11747
rect 2004 11716 2145 11744
rect 2004 11704 2010 11716
rect 2133 11713 2145 11716
rect 2179 11713 2191 11747
rect 4172 11744 4200 11772
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4172 11716 4445 11744
rect 2133 11707 2191 11713
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 5074 11744 5080 11756
rect 5035 11716 5080 11744
rect 4433 11707 4491 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 14182 11744 14188 11756
rect 13587 11716 14188 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19300 11716 19809 11744
rect 19300 11704 19306 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 3396 11679 3454 11685
rect 3396 11645 3408 11679
rect 3442 11676 3454 11679
rect 4062 11676 4068 11688
rect 3442 11648 4068 11676
rect 3442 11645 3454 11648
rect 3396 11639 3454 11645
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11577 1915 11611
rect 1857 11571 1915 11577
rect 1872 11540 1900 11571
rect 3896 11552 3924 11648
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 14436 11679 14494 11685
rect 14436 11676 14448 11679
rect 13786 11648 14448 11676
rect 7101 11611 7159 11617
rect 7101 11577 7113 11611
rect 7147 11608 7159 11611
rect 7282 11608 7288 11620
rect 7147 11580 7288 11608
rect 7147 11577 7159 11580
rect 7101 11571 7159 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 11333 11611 11391 11617
rect 11333 11577 11345 11611
rect 11379 11608 11391 11611
rect 12526 11608 12532 11620
rect 11379 11580 12532 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12636 11580 12909 11608
rect 2406 11540 2412 11552
rect 1872 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11540 2470 11552
rect 2777 11543 2835 11549
rect 2777 11540 2789 11543
rect 2464 11512 2789 11540
rect 2464 11500 2470 11512
rect 2777 11509 2789 11512
rect 2823 11509 2835 11543
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 2777 11503 2835 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12636 11549 12664 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 13786 11608 13814 11648
rect 14436 11645 14448 11648
rect 14482 11676 14494 11679
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14482 11648 14841 11676
rect 14482 11645 14494 11648
rect 14436 11639 14494 11645
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 18484 11679 18542 11685
rect 18484 11645 18496 11679
rect 18530 11676 18542 11679
rect 18598 11676 18604 11688
rect 18530 11648 18604 11676
rect 18530 11645 18542 11648
rect 18484 11639 18542 11645
rect 18598 11636 18604 11648
rect 18656 11676 18662 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18656 11648 18889 11676
rect 18656 11636 18662 11648
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 19334 11608 19340 11620
rect 13596 11580 13814 11608
rect 19247 11580 19340 11608
rect 13596 11568 13602 11580
rect 19334 11568 19340 11580
rect 19392 11608 19398 11620
rect 19521 11611 19579 11617
rect 19521 11608 19533 11611
rect 19392 11580 19533 11608
rect 19392 11568 19398 11580
rect 19521 11577 19533 11580
rect 19567 11608 19579 11611
rect 19610 11608 19616 11620
rect 19567 11580 19616 11608
rect 19567 11577 19579 11580
rect 19521 11571 19579 11577
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 12621 11543 12679 11549
rect 12621 11540 12633 11543
rect 11848 11512 12633 11540
rect 11848 11500 11854 11512
rect 12621 11509 12633 11512
rect 12667 11509 12679 11543
rect 12621 11503 12679 11509
rect 20533 11543 20591 11549
rect 20533 11509 20545 11543
rect 20579 11540 20591 11543
rect 20714 11540 20720 11552
rect 20579 11512 20720 11540
rect 20579 11509 20591 11512
rect 20533 11503 20591 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 21436 11472
rect 1104 11398 8497 11450
rect 8549 11398 8561 11450
rect 8613 11398 8625 11450
rect 8677 11398 8689 11450
rect 8741 11398 16012 11450
rect 16064 11398 16076 11450
rect 16128 11398 16140 11450
rect 16192 11398 16204 11450
rect 16256 11398 21436 11450
rect 1104 11376 21436 11398
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6638 11336 6644 11348
rect 6135 11308 6644 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 8343 11339 8401 11345
rect 8343 11336 8355 11339
rect 7340 11308 8355 11336
rect 7340 11296 7346 11308
rect 8343 11305 8355 11308
rect 8389 11305 8401 11339
rect 12894 11336 12900 11348
rect 12855 11308 12900 11336
rect 8343 11299 8401 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 2406 11268 2412 11280
rect 2367 11240 2412 11268
rect 2406 11228 2412 11240
rect 2464 11228 2470 11280
rect 5074 11268 5080 11280
rect 5035 11240 5080 11268
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 11517 11271 11575 11277
rect 11517 11237 11529 11271
rect 11563 11268 11575 11271
rect 11698 11268 11704 11280
rect 11563 11240 11704 11268
rect 11563 11237 11575 11240
rect 11517 11231 11575 11237
rect 11698 11228 11704 11240
rect 11756 11228 11762 11280
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 12710 11268 12716 11280
rect 12584 11240 12716 11268
rect 12584 11228 12590 11240
rect 12710 11228 12716 11240
rect 12768 11268 12774 11280
rect 13081 11271 13139 11277
rect 13081 11268 13093 11271
rect 12768 11240 13093 11268
rect 12768 11228 12774 11240
rect 13081 11237 13093 11240
rect 13127 11237 13139 11271
rect 18414 11268 18420 11280
rect 18375 11240 18420 11268
rect 13081 11231 13139 11237
rect 18414 11228 18420 11240
rect 18472 11228 18478 11280
rect 19981 11271 20039 11277
rect 19981 11237 19993 11271
rect 20027 11268 20039 11271
rect 20254 11268 20260 11280
rect 20027 11240 20260 11268
rect 20027 11237 20039 11240
rect 19981 11231 20039 11237
rect 20254 11228 20260 11240
rect 20312 11228 20318 11280
rect 7098 11200 7104 11212
rect 7059 11172 7104 11200
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 8294 11200 8300 11212
rect 8251 11172 8300 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11101 1823 11135
rect 4430 11132 4436 11144
rect 4391 11104 4436 11132
rect 1765 11095 1823 11101
rect 1670 11024 1676 11076
rect 1728 11064 1734 11076
rect 1780 11064 1808 11095
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 11790 11132 11796 11144
rect 11751 11104 11796 11132
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 13538 11132 13544 11144
rect 13499 11104 13544 11132
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 17770 11132 17776 11144
rect 16715 11104 17776 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 19334 11132 19340 11144
rect 19295 11104 19340 11132
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 1728 11036 1808 11064
rect 1728 11024 1734 11036
rect 7282 10996 7288 11008
rect 7243 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 18196 10968 18705 10996
rect 18196 10956 18202 10968
rect 18693 10965 18705 10968
rect 18739 10965 18751 10999
rect 18693 10959 18751 10965
rect 1104 10906 21436 10928
rect 1104 10854 4739 10906
rect 4791 10854 4803 10906
rect 4855 10854 4867 10906
rect 4919 10854 4931 10906
rect 4983 10854 12255 10906
rect 12307 10854 12319 10906
rect 12371 10854 12383 10906
rect 12435 10854 12447 10906
rect 12499 10854 19770 10906
rect 19822 10854 19834 10906
rect 19886 10854 19898 10906
rect 19950 10854 19962 10906
rect 20014 10854 21436 10906
rect 1104 10832 21436 10854
rect 3326 10792 3332 10804
rect 3287 10764 3332 10792
rect 3326 10752 3332 10764
rect 3384 10792 3390 10804
rect 3384 10764 3648 10792
rect 3384 10752 3390 10764
rect 2406 10656 2412 10668
rect 2367 10628 2412 10656
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 3620 10665 3648 10764
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4488 10764 4537 10792
rect 4488 10752 4494 10764
rect 4525 10761 4537 10764
rect 4571 10792 4583 10795
rect 5215 10795 5273 10801
rect 5215 10792 5227 10795
rect 4571 10764 5227 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 5215 10761 5227 10764
rect 5261 10761 5273 10795
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 5215 10755 5273 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 17770 10792 17776 10804
rect 17731 10764 17776 10792
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 13538 10724 13544 10736
rect 13499 10696 13544 10724
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 16071 10727 16129 10733
rect 16071 10693 16083 10727
rect 16117 10724 16129 10727
rect 19061 10727 19119 10733
rect 19061 10724 19073 10727
rect 16117 10696 19073 10724
rect 16117 10693 16129 10696
rect 16071 10687 16129 10693
rect 19061 10693 19073 10696
rect 19107 10724 19119 10727
rect 19334 10724 19340 10736
rect 19107 10696 19340 10724
rect 19107 10693 19119 10696
rect 19061 10687 19119 10693
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 19610 10684 19616 10736
rect 19668 10724 19674 10736
rect 20257 10727 20315 10733
rect 20257 10724 20269 10727
rect 19668 10696 20269 10724
rect 19668 10684 19674 10696
rect 20257 10693 20269 10696
rect 20303 10693 20315 10727
rect 20257 10687 20315 10693
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11790 10656 11796 10668
rect 11563 10628 11796 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 17083 10659 17141 10665
rect 17083 10625 17095 10659
rect 17129 10656 17141 10659
rect 18138 10656 18144 10668
rect 17129 10628 18144 10656
rect 17129 10625 17141 10628
rect 17083 10619 17141 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18414 10656 18420 10668
rect 18375 10628 18420 10656
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10656 19579 10659
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19567 10628 19717 10656
rect 19567 10625 19579 10628
rect 19521 10619 19579 10625
rect 19705 10625 19717 10628
rect 19751 10656 19763 10659
rect 20070 10656 20076 10668
rect 19751 10628 20076 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 5144 10591 5202 10597
rect 5144 10557 5156 10591
rect 5190 10588 5202 10591
rect 5626 10588 5632 10600
rect 5190 10560 5632 10588
rect 5190 10557 5202 10560
rect 5144 10551 5202 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 16000 10591 16058 10597
rect 16000 10557 16012 10591
rect 16046 10588 16058 10591
rect 16996 10591 17054 10597
rect 16046 10560 16528 10588
rect 16046 10557 16058 10560
rect 16000 10551 16058 10557
rect 2038 10520 2044 10532
rect 1999 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 4249 10523 4307 10529
rect 4249 10489 4261 10523
rect 4295 10520 4307 10523
rect 4890 10520 4896 10532
rect 4295 10492 4896 10520
rect 4295 10489 4307 10492
rect 4249 10483 4307 10489
rect 4890 10480 4896 10492
rect 4948 10520 4954 10532
rect 8386 10520 8392 10532
rect 4948 10492 8392 10520
rect 4948 10480 4954 10492
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 10873 10523 10931 10529
rect 10873 10489 10885 10523
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12802 10520 12808 10532
rect 12299 10492 12808 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 5626 10452 5632 10464
rect 5587 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 8294 10452 8300 10464
rect 8255 10424 8300 10452
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 10594 10452 10600 10464
rect 10555 10424 10600 10452
rect 10594 10412 10600 10424
rect 10652 10452 10658 10464
rect 10888 10452 10916 10483
rect 12802 10480 12808 10492
rect 12860 10520 12866 10532
rect 12989 10523 13047 10529
rect 12989 10520 13001 10523
rect 12860 10492 13001 10520
rect 12860 10480 12866 10492
rect 12989 10489 13001 10492
rect 13035 10489 13047 10523
rect 12989 10483 13047 10489
rect 11790 10452 11796 10464
rect 10652 10424 10916 10452
rect 11751 10424 11796 10452
rect 10652 10412 10658 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 16500 10461 16528 10560
rect 16996 10557 17008 10591
rect 17042 10588 17054 10591
rect 17402 10588 17408 10600
rect 17042 10560 17408 10588
rect 17042 10557 17054 10560
rect 16996 10551 17054 10557
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 16485 10455 16543 10461
rect 16485 10421 16497 10455
rect 16531 10452 16543 10455
rect 21818 10452 21824 10464
rect 16531 10424 21824 10452
rect 16531 10421 16543 10424
rect 16485 10415 16543 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 1104 10362 21436 10384
rect 1104 10310 8497 10362
rect 8549 10310 8561 10362
rect 8613 10310 8625 10362
rect 8677 10310 8689 10362
rect 8741 10310 16012 10362
rect 16064 10310 16076 10362
rect 16128 10310 16140 10362
rect 16192 10310 16204 10362
rect 16256 10310 21436 10362
rect 1104 10288 21436 10310
rect 10183 10251 10241 10257
rect 10183 10217 10195 10251
rect 10229 10248 10241 10251
rect 10594 10248 10600 10260
rect 10229 10220 10600 10248
rect 10229 10217 10241 10220
rect 10183 10211 10241 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 19797 10251 19855 10257
rect 19797 10217 19809 10251
rect 19843 10248 19855 10251
rect 20162 10248 20168 10260
rect 19843 10220 20168 10248
rect 19843 10217 19855 10220
rect 19797 10211 19855 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 2222 10180 2228 10192
rect 2183 10152 2228 10180
rect 2222 10140 2228 10152
rect 2280 10140 2286 10192
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 17460 10152 19656 10180
rect 17460 10140 17466 10152
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10134 10112 10140 10124
rect 10091 10084 10140 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11476 10115 11534 10121
rect 11476 10081 11488 10115
rect 11522 10112 11534 10115
rect 11698 10112 11704 10124
rect 11522 10084 11704 10112
rect 11522 10081 11534 10084
rect 11476 10075 11534 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14642 10112 14648 10124
rect 14139 10084 14648 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 19628 10121 19656 10152
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 20162 10112 20168 10124
rect 19659 10084 20168 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 20162 10072 20168 10084
rect 20220 10072 20226 10124
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4890 10044 4896 10056
rect 4851 10016 4896 10044
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 11563 10047 11621 10053
rect 11563 10013 11575 10047
rect 11609 10044 11621 10047
rect 12529 10047 12587 10053
rect 12529 10044 12541 10047
rect 11609 10016 12541 10044
rect 11609 10013 11621 10016
rect 11563 10007 11621 10013
rect 12529 10013 12541 10016
rect 12575 10044 12587 10047
rect 12618 10044 12624 10056
rect 12575 10016 12624 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 2774 9976 2780 9988
rect 2735 9948 2780 9976
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 18414 9976 18420 9988
rect 18375 9948 18420 9976
rect 18414 9936 18420 9948
rect 18472 9936 18478 9988
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 1104 9818 21436 9840
rect 1104 9766 4739 9818
rect 4791 9766 4803 9818
rect 4855 9766 4867 9818
rect 4919 9766 4931 9818
rect 4983 9766 12255 9818
rect 12307 9766 12319 9818
rect 12371 9766 12383 9818
rect 12435 9766 12447 9818
rect 12499 9766 19770 9818
rect 19822 9766 19834 9818
rect 19886 9766 19898 9818
rect 19950 9766 19962 9818
rect 20014 9766 21436 9818
rect 1104 9744 21436 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2317 9707 2375 9713
rect 2317 9704 2329 9707
rect 2280 9676 2329 9704
rect 2280 9664 2286 9676
rect 2317 9673 2329 9676
rect 2363 9673 2375 9707
rect 2317 9667 2375 9673
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 4212 9676 4721 9704
rect 4212 9664 4218 9676
rect 4709 9673 4721 9676
rect 4755 9704 4767 9707
rect 5810 9704 5816 9716
rect 4755 9676 5816 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 11471 9707 11529 9713
rect 11471 9673 11483 9707
rect 11517 9704 11529 9707
rect 11790 9704 11796 9716
rect 11517 9676 11796 9704
rect 11517 9673 11529 9676
rect 11471 9667 11529 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 14277 9707 14335 9713
rect 14277 9673 14289 9707
rect 14323 9704 14335 9707
rect 15194 9704 15200 9716
rect 14323 9676 15200 9704
rect 14323 9673 14335 9676
rect 14277 9667 14335 9673
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 17862 9704 17868 9716
rect 17823 9676 17868 9704
rect 17862 9664 17868 9676
rect 17920 9704 17926 9716
rect 18187 9707 18245 9713
rect 18187 9704 18199 9707
rect 17920 9676 18199 9704
rect 17920 9664 17926 9676
rect 18187 9673 18199 9676
rect 18233 9673 18245 9707
rect 18187 9667 18245 9673
rect 19426 9664 19432 9716
rect 19484 9704 19490 9716
rect 19797 9707 19855 9713
rect 19797 9704 19809 9707
rect 19484 9676 19809 9704
rect 19484 9664 19490 9676
rect 19797 9673 19809 9676
rect 19843 9673 19855 9707
rect 20162 9704 20168 9716
rect 20123 9676 20168 9704
rect 19797 9667 19855 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 2038 9596 2044 9648
rect 2096 9636 2102 9648
rect 5307 9639 5365 9645
rect 5307 9636 5319 9639
rect 2096 9608 5319 9636
rect 2096 9596 2102 9608
rect 5307 9605 5319 9608
rect 5353 9605 5365 9639
rect 10042 9636 10048 9648
rect 10003 9608 10048 9636
rect 5307 9599 5365 9605
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 4062 9568 4068 9580
rect 2648 9540 4068 9568
rect 2648 9528 2654 9540
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4295 9571 4353 9577
rect 4295 9537 4307 9571
rect 4341 9568 4353 9571
rect 4614 9568 4620 9580
rect 4341 9540 4620 9568
rect 4341 9537 4353 9540
rect 4295 9531 4353 9537
rect 4614 9528 4620 9540
rect 4672 9568 4678 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4672 9540 4997 9568
rect 4672 9528 4678 9540
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 10134 9568 10140 9580
rect 4985 9531 5043 9537
rect 8864 9540 10140 9568
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9500 1458 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1452 9472 1961 9500
rect 1452 9460 1458 9472
rect 1949 9469 1961 9472
rect 1995 9469 2007 9503
rect 2498 9500 2504 9512
rect 2459 9472 2504 9500
rect 1949 9463 2007 9469
rect 1964 9432 1992 9463
rect 2498 9460 2504 9472
rect 2556 9500 2562 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2556 9472 3065 9500
rect 2556 9460 2562 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 5236 9503 5294 9509
rect 5236 9469 5248 9503
rect 5282 9500 5294 9503
rect 5718 9500 5724 9512
rect 5282 9472 5724 9500
rect 5282 9469 5294 9472
rect 5236 9463 5294 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 8864 9509 8892 9540
rect 10134 9528 10140 9540
rect 10192 9568 10198 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10192 9540 10425 9568
rect 10192 9528 10198 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 10413 9531 10471 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 14458 9568 14464 9580
rect 13688 9540 14464 9568
rect 13688 9528 13694 9540
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 8424 9503 8482 9509
rect 8424 9469 8436 9503
rect 8470 9500 8482 9503
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8470 9472 8861 9500
rect 8470 9469 8482 9472
rect 8424 9463 8482 9469
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 11400 9503 11458 9509
rect 11400 9469 11412 9503
rect 11446 9500 11458 9503
rect 13998 9500 14004 9512
rect 11446 9472 12020 9500
rect 13911 9472 14004 9500
rect 11446 9469 11458 9472
rect 11400 9463 11458 9469
rect 8439 9432 8467 9463
rect 1964 9404 8467 9432
rect 8527 9435 8585 9441
rect 8527 9401 8539 9435
rect 8573 9432 8585 9435
rect 9217 9435 9275 9441
rect 9217 9432 9229 9435
rect 8573 9404 9229 9432
rect 8573 9401 8585 9404
rect 8527 9395 8585 9401
rect 9217 9401 9229 9404
rect 9263 9432 9275 9435
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 9263 9404 9505 9432
rect 9263 9401 9275 9404
rect 9217 9395 9275 9401
rect 9493 9401 9505 9404
rect 9539 9401 9551 9435
rect 9493 9395 9551 9401
rect 11992 9376 12020 9472
rect 13998 9460 14004 9472
rect 14056 9500 14062 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 14056 9472 14105 9500
rect 14056 9460 14062 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 18116 9503 18174 9509
rect 18116 9469 18128 9503
rect 18162 9500 18174 9503
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 18162 9472 18644 9500
rect 18162 9469 18174 9472
rect 18116 9463 18174 9469
rect 12526 9432 12532 9444
rect 12439 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9432 12590 9444
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 12584 9404 13461 9432
rect 12584 9392 12590 9404
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 18616 9376 18644 9472
rect 19444 9472 19625 9500
rect 19444 9376 19472 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 106 9324 112 9376
rect 164 9364 170 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 164 9336 1593 9364
rect 164 9324 170 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 2682 9364 2688 9376
rect 2643 9336 2688 9364
rect 1581 9327 1639 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 5718 9364 5724 9376
rect 3568 9336 5724 9364
rect 3568 9324 3574 9336
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 11790 9364 11796 9376
rect 11751 9336 11796 9364
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 12032 9336 12173 9364
rect 12032 9324 12038 9336
rect 12161 9333 12173 9336
rect 12207 9333 12219 9367
rect 18598 9364 18604 9376
rect 18559 9336 18604 9364
rect 12161 9327 12219 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 1104 9274 21436 9296
rect 1104 9222 8497 9274
rect 8549 9222 8561 9274
rect 8613 9222 8625 9274
rect 8677 9222 8689 9274
rect 8741 9222 16012 9274
rect 16064 9222 16076 9274
rect 16128 9222 16140 9274
rect 16192 9222 16204 9274
rect 16256 9222 21436 9274
rect 1104 9200 21436 9222
rect 1535 9163 1593 9169
rect 1535 9129 1547 9163
rect 1581 9160 1593 9163
rect 1670 9160 1676 9172
rect 1581 9132 1676 9160
rect 1581 9129 1593 9132
rect 1535 9123 1593 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 11103 9163 11161 9169
rect 11103 9129 11115 9163
rect 11149 9160 11161 9163
rect 12526 9160 12532 9172
rect 11149 9132 12532 9160
rect 11149 9129 11161 9132
rect 11103 9123 11161 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12676 9132 13001 9160
rect 12676 9120 12682 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 13679 9163 13737 9169
rect 13679 9129 13691 9163
rect 13725 9160 13737 9163
rect 13998 9160 14004 9172
rect 13725 9132 14004 9160
rect 13725 9129 13737 9132
rect 13679 9123 13737 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 19797 9163 19855 9169
rect 19797 9129 19809 9163
rect 19843 9160 19855 9163
rect 20162 9160 20168 9172
rect 19843 9132 20168 9160
rect 19843 9129 19855 9132
rect 19797 9123 19855 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 2498 9092 2504 9104
rect 1479 9064 2504 9092
rect 1479 9033 1507 9064
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 1578 9024 1584 9036
rect 1510 8996 1584 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 10962 9024 10968 9036
rect 10919 8996 10968 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 13576 9027 13634 9033
rect 13576 9024 13588 9027
rect 12912 8996 13588 9024
rect 12912 8968 12940 8996
rect 13576 8993 13588 8996
rect 13622 8993 13634 9027
rect 13576 8987 13634 8993
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 18656 8996 19625 9024
rect 18656 8984 18662 8996
rect 19613 8993 19625 8996
rect 19659 9024 19671 9027
rect 20254 9024 20260 9036
rect 19659 8996 20260 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20254 8984 20260 8996
rect 20312 8984 20318 9036
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2774 8956 2780 8968
rect 2735 8928 2780 8956
rect 2774 8916 2780 8928
rect 2832 8956 2838 8968
rect 4154 8956 4160 8968
rect 2832 8928 4160 8956
rect 2832 8916 2838 8928
rect 4154 8916 4160 8928
rect 4212 8956 4218 8968
rect 4614 8956 4620 8968
rect 4212 8928 4257 8956
rect 4575 8928 4620 8956
rect 4212 8916 4218 8928
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8956 7159 8959
rect 7834 8956 7840 8968
rect 7147 8928 7840 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 12066 8956 12072 8968
rect 12027 8928 12072 8956
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 12894 8956 12900 8968
rect 12759 8928 12900 8956
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7616 8860 7665 8888
rect 7616 8848 7622 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 17402 8888 17408 8900
rect 12032 8860 17408 8888
rect 12032 8848 12038 8860
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 1104 8730 21436 8752
rect 1104 8678 4739 8730
rect 4791 8678 4803 8730
rect 4855 8678 4867 8730
rect 4919 8678 4931 8730
rect 4983 8678 12255 8730
rect 12307 8678 12319 8730
rect 12371 8678 12383 8730
rect 12435 8678 12447 8730
rect 12499 8678 19770 8730
rect 19822 8678 19834 8730
rect 19886 8678 19898 8730
rect 19950 8678 19962 8730
rect 20014 8678 21436 8730
rect 1104 8656 21436 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2363 8619 2421 8625
rect 2363 8585 2375 8619
rect 2409 8616 2421 8619
rect 2498 8616 2504 8628
rect 2409 8588 2504 8616
rect 2409 8585 2421 8588
rect 2363 8579 2421 8585
rect 2498 8576 2504 8588
rect 2556 8616 2562 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2556 8588 3065 8616
rect 2556 8576 2562 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4212 8588 4261 8616
rect 4212 8576 4218 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 7834 8616 7840 8628
rect 7795 8588 7840 8616
rect 4249 8579 4307 8585
rect 7834 8576 7840 8588
rect 7892 8616 7898 8628
rect 8527 8619 8585 8625
rect 8527 8616 8539 8619
rect 7892 8588 8539 8616
rect 7892 8576 7898 8588
rect 8527 8585 8539 8588
rect 8573 8585 8585 8619
rect 8527 8579 8585 8585
rect 18739 8619 18797 8625
rect 18739 8585 18751 8619
rect 18785 8616 18797 8619
rect 19426 8616 19432 8628
rect 18785 8588 19432 8616
rect 18785 8585 18797 8588
rect 18739 8579 18797 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 3881 8551 3939 8557
rect 3881 8517 3893 8551
rect 3927 8548 3939 8551
rect 3970 8548 3976 8560
rect 3927 8520 3976 8548
rect 3927 8517 3939 8520
rect 3881 8511 3939 8517
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 19797 8551 19855 8557
rect 19797 8517 19809 8551
rect 19843 8548 19855 8551
rect 20162 8548 20168 8560
rect 19843 8520 20168 8548
rect 19843 8517 19855 8520
rect 19797 8511 19855 8517
rect 20162 8508 20168 8520
rect 20220 8508 20226 8560
rect 3326 8480 3332 8492
rect 3239 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8480 3390 8492
rect 4939 8483 4997 8489
rect 4939 8480 4951 8483
rect 3384 8452 4951 8480
rect 3384 8440 3390 8452
rect 4939 8449 4951 8452
rect 4985 8449 4997 8483
rect 7558 8480 7564 8492
rect 7519 8452 7564 8480
rect 4939 8443 4997 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8480 12958 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 12952 8452 13553 8480
rect 12952 8440 12958 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14516 8452 15025 8480
rect 14516 8440 14522 8452
rect 15013 8449 15025 8452
rect 15059 8480 15071 8483
rect 19242 8480 19248 8492
rect 15059 8452 19248 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 2292 8415 2350 8421
rect 2292 8381 2304 8415
rect 2338 8412 2350 8415
rect 2590 8412 2596 8424
rect 2338 8384 2596 8412
rect 2338 8381 2350 8384
rect 2292 8375 2350 8381
rect 2590 8372 2596 8384
rect 2648 8412 2654 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2648 8384 2697 8412
rect 2648 8372 2654 8384
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 4852 8415 4910 8421
rect 4852 8381 4864 8415
rect 4898 8412 4910 8415
rect 4898 8384 5396 8412
rect 4898 8381 4910 8384
rect 4852 8375 4910 8381
rect 5368 8288 5396 8384
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8456 8415 8514 8421
rect 8456 8412 8468 8415
rect 7984 8384 8468 8412
rect 7984 8372 7990 8384
rect 8456 8381 8468 8384
rect 8502 8412 8514 8415
rect 18668 8415 18726 8421
rect 8502 8384 8984 8412
rect 8502 8381 8514 8384
rect 8456 8375 8514 8381
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6914 8344 6920 8356
rect 6687 8316 6920 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 5350 8276 5356 8288
rect 5311 8248 5356 8276
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 8956 8285 8984 8384
rect 18668 8381 18680 8415
rect 18714 8412 18726 8415
rect 19058 8412 19064 8424
rect 18714 8384 19064 8412
rect 18714 8381 18726 8384
rect 18668 8375 18726 8381
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8412 19579 8415
rect 19610 8412 19616 8424
rect 19567 8384 19616 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11379 8316 12173 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 12161 8313 12173 8316
rect 12207 8344 12219 8347
rect 12621 8347 12679 8353
rect 12621 8344 12633 8347
rect 12207 8316 12633 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 12621 8313 12633 8316
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 8941 8279 8999 8285
rect 8941 8245 8953 8279
rect 8987 8276 8999 8279
rect 10962 8276 10968 8288
rect 8987 8248 10968 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11112 8248 11805 8276
rect 11112 8236 11118 8248
rect 11793 8245 11805 8248
rect 11839 8276 11851 8279
rect 12066 8276 12072 8288
rect 11839 8248 12072 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 14185 8279 14243 8285
rect 14185 8245 14197 8279
rect 14231 8276 14243 8279
rect 14274 8276 14280 8288
rect 14231 8248 14280 8276
rect 14231 8245 14243 8248
rect 14185 8239 14243 8245
rect 14274 8236 14280 8248
rect 14332 8276 14338 8288
rect 14384 8276 14412 8307
rect 20254 8276 20260 8288
rect 14332 8248 14412 8276
rect 20215 8248 20260 8276
rect 14332 8236 14338 8248
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 1104 8186 21436 8208
rect 1104 8134 8497 8186
rect 8549 8134 8561 8186
rect 8613 8134 8625 8186
rect 8677 8134 8689 8186
rect 8741 8134 16012 8186
rect 16064 8134 16076 8186
rect 16128 8134 16140 8186
rect 16192 8134 16204 8186
rect 16256 8134 21436 8186
rect 1104 8112 21436 8134
rect 3326 8072 3332 8084
rect 3287 8044 3332 8072
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 3660 8044 4154 8072
rect 3660 8032 3666 8044
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 3970 8004 3976 8016
rect 2915 7976 3976 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 4126 8004 4154 8044
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7055 8075 7113 8081
rect 7055 8072 7067 8075
rect 6972 8044 7067 8072
rect 6972 8032 6978 8044
rect 7055 8041 7067 8044
rect 7101 8041 7113 8075
rect 7055 8035 7113 8041
rect 19475 8075 19533 8081
rect 19475 8041 19487 8075
rect 19521 8072 19533 8075
rect 19610 8072 19616 8084
rect 19521 8044 19616 8072
rect 19521 8041 19533 8044
rect 19475 8035 19533 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 4126 7976 9628 8004
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6914 7936 6920 7948
rect 6875 7908 6920 7936
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 9600 7936 9628 7976
rect 10318 7936 10324 7948
rect 10376 7945 10382 7948
rect 10376 7939 10414 7945
rect 9600 7908 10324 7936
rect 10318 7896 10324 7908
rect 10402 7905 10414 7939
rect 10376 7899 10414 7905
rect 10376 7896 10382 7899
rect 19242 7896 19248 7948
rect 19300 7936 19306 7948
rect 19372 7939 19430 7945
rect 19372 7936 19384 7939
rect 19300 7908 19384 7936
rect 19300 7896 19306 7908
rect 19372 7905 19384 7908
rect 19418 7905 19430 7939
rect 19372 7899 19430 7905
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 4338 7868 4344 7880
rect 4299 7840 4344 7868
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 10459 7871 10517 7877
rect 10459 7837 10471 7871
rect 10505 7868 10517 7871
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10505 7840 11437 7868
rect 10505 7837 10517 7840
rect 10459 7831 10517 7837
rect 11425 7837 11437 7840
rect 11471 7868 11483 7871
rect 11514 7868 11520 7880
rect 11471 7840 11520 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 12066 7868 12072 7880
rect 12027 7840 12072 7868
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 13964 7840 15301 7868
rect 13964 7828 13970 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 14274 7800 14280 7812
rect 14235 7772 14280 7800
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6730 7732 6736 7744
rect 6043 7704 6736 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 10778 7732 10784 7744
rect 10739 7704 10784 7732
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 1104 7642 21436 7664
rect 1104 7590 4739 7642
rect 4791 7590 4803 7642
rect 4855 7590 4867 7642
rect 4919 7590 4931 7642
rect 4983 7590 12255 7642
rect 12307 7590 12319 7642
rect 12371 7590 12383 7642
rect 12435 7590 12447 7642
rect 12499 7590 19770 7642
rect 19822 7590 19834 7642
rect 19886 7590 19898 7642
rect 19950 7590 19962 7642
rect 20014 7590 21436 7642
rect 1104 7568 21436 7590
rect 1535 7531 1593 7537
rect 1535 7497 1547 7531
rect 1581 7528 1593 7531
rect 2222 7528 2228 7540
rect 1581 7500 2228 7528
rect 1581 7497 1593 7500
rect 1535 7491 1593 7497
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 4338 7528 4344 7540
rect 3988 7500 4344 7528
rect 3988 7401 4016 7500
rect 4338 7488 4344 7500
rect 4396 7528 4402 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4396 7500 4445 7528
rect 4396 7488 4402 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 5810 7528 5816 7540
rect 5771 7500 5816 7528
rect 4433 7491 4491 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 10318 7528 10324 7540
rect 10279 7500 10324 7528
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11514 7528 11520 7540
rect 11475 7500 11520 7528
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12943 7531 13001 7537
rect 12943 7497 12955 7531
rect 12989 7528 13001 7531
rect 13722 7528 13728 7540
rect 12989 7500 13728 7528
rect 12989 7497 13001 7500
rect 12943 7491 13001 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19242 7528 19248 7540
rect 18831 7500 19248 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 13354 7460 13360 7472
rect 13315 7432 13360 7460
rect 13354 7420 13360 7432
rect 13412 7420 13418 7472
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 6914 7392 6920 7404
rect 5224 7364 6920 7392
rect 5224 7352 5230 7364
rect 6914 7352 6920 7364
rect 6972 7392 6978 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 9631 7395 9689 7401
rect 9631 7361 9643 7395
rect 9677 7392 9689 7395
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 9677 7364 10609 7392
rect 9677 7361 9689 7364
rect 9631 7355 9689 7361
rect 10597 7361 10609 7364
rect 10643 7392 10655 7395
rect 10778 7392 10784 7404
rect 10643 7364 10784 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 1302 7284 1308 7336
rect 1360 7324 1366 7336
rect 1432 7327 1490 7333
rect 1432 7324 1444 7327
rect 1360 7296 1444 7324
rect 1360 7284 1366 7296
rect 1432 7293 1444 7296
rect 1478 7324 1490 7327
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1478 7296 1869 7324
rect 1478 7293 1490 7296
rect 1432 7287 1490 7293
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5020 7327 5078 7333
rect 5020 7324 5032 7327
rect 4672 7296 5032 7324
rect 4672 7284 4678 7296
rect 5020 7293 5032 7296
rect 5066 7324 5078 7327
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5066 7296 5457 7324
rect 5066 7293 5078 7296
rect 5020 7287 5078 7293
rect 5445 7293 5457 7296
rect 5491 7293 5503 7327
rect 7024 7324 7052 7355
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11054 7392 11060 7404
rect 11015 7364 11060 7392
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 9528 7327 9586 7333
rect 9528 7324 9540 7327
rect 7024 7296 9540 7324
rect 5445 7287 5503 7293
rect 9528 7293 9540 7296
rect 9574 7324 9586 7327
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9574 7296 9965 7324
rect 9574 7293 9586 7296
rect 9528 7287 9586 7293
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 12872 7327 12930 7333
rect 12872 7293 12884 7327
rect 12918 7324 12930 7327
rect 13372 7324 13400 7420
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 13906 7392 13912 7404
rect 13771 7364 13912 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14332 7364 14565 7392
rect 14332 7352 14338 7364
rect 14553 7361 14565 7364
rect 14599 7392 14611 7395
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 14599 7364 15761 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 19518 7392 19524 7404
rect 19116 7364 19524 7392
rect 19116 7352 19122 7364
rect 19518 7352 19524 7364
rect 19576 7392 19582 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19576 7364 19625 7392
rect 19576 7352 19582 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 12918 7296 13400 7324
rect 12918 7293 12930 7296
rect 12872 7287 12930 7293
rect 15473 7259 15531 7265
rect 15473 7256 15485 7259
rect 15212 7228 15485 7256
rect 15212 7200 15240 7228
rect 15473 7225 15485 7228
rect 15519 7225 15531 7259
rect 15473 7219 15531 7225
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7256 18291 7259
rect 19061 7259 19119 7265
rect 19061 7256 19073 7259
rect 18279 7228 19073 7256
rect 18279 7225 18291 7228
rect 18233 7219 18291 7225
rect 19061 7225 19073 7228
rect 19107 7256 19119 7259
rect 19337 7259 19395 7265
rect 19337 7256 19349 7259
rect 19107 7228 19349 7256
rect 19107 7225 19119 7228
rect 19061 7219 19119 7225
rect 19337 7225 19349 7228
rect 19383 7225 19395 7259
rect 19337 7219 19395 7225
rect 5123 7191 5181 7197
rect 5123 7157 5135 7191
rect 5169 7188 5181 7191
rect 5718 7188 5724 7200
rect 5169 7160 5724 7188
rect 5169 7157 5181 7160
rect 5123 7151 5181 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 1104 7098 21436 7120
rect 1104 7046 8497 7098
rect 8549 7046 8561 7098
rect 8613 7046 8625 7098
rect 8677 7046 8689 7098
rect 8741 7046 16012 7098
rect 16064 7046 16076 7098
rect 16128 7046 16140 7098
rect 16192 7046 16204 7098
rect 16256 7046 21436 7098
rect 1104 7024 21436 7046
rect 13587 6987 13645 6993
rect 13587 6953 13599 6987
rect 13633 6984 13645 6987
rect 15194 6984 15200 6996
rect 13633 6956 15200 6984
rect 13633 6953 13645 6956
rect 13587 6947 13645 6953
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 11054 6916 11060 6928
rect 11015 6888 11060 6916
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 13722 6876 13728 6928
rect 13780 6916 13786 6928
rect 13909 6919 13967 6925
rect 13909 6916 13921 6919
rect 13780 6888 13921 6916
rect 13780 6876 13786 6888
rect 13909 6885 13921 6888
rect 13955 6885 13967 6919
rect 13909 6879 13967 6885
rect 5166 6848 5172 6860
rect 5127 6820 5172 6848
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6270 6848 6276 6860
rect 5776 6820 6276 6848
rect 5776 6808 5782 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 7926 6848 7932 6860
rect 7887 6820 7932 6848
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 17288 6851 17346 6857
rect 17288 6817 17300 6851
rect 17334 6848 17346 6851
rect 17402 6848 17408 6860
rect 17334 6820 17408 6848
rect 17334 6817 17346 6820
rect 17288 6811 17346 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 10410 6780 10416 6792
rect 10371 6752 10416 6780
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 11992 6712 12020 6743
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 12124 6752 12265 6780
rect 12124 6740 12130 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 12253 6743 12311 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 19242 6780 19248 6792
rect 19203 6752 19248 6780
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 11940 6684 12020 6712
rect 11940 6672 11946 6684
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 6178 6644 6184 6656
rect 5399 6616 6184 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6454 6644 6460 6656
rect 6415 6616 6460 6644
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8938 6644 8944 6656
rect 8159 6616 8944 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 17359 6647 17417 6653
rect 17359 6613 17371 6647
rect 17405 6644 17417 6647
rect 17770 6644 17776 6656
rect 17405 6616 17776 6644
rect 17405 6613 17417 6616
rect 17359 6607 17417 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 1104 6554 21436 6576
rect 1104 6502 4739 6554
rect 4791 6502 4803 6554
rect 4855 6502 4867 6554
rect 4919 6502 4931 6554
rect 4983 6502 12255 6554
rect 12307 6502 12319 6554
rect 12371 6502 12383 6554
rect 12435 6502 12447 6554
rect 12499 6502 19770 6554
rect 19822 6502 19834 6554
rect 19886 6502 19898 6554
rect 19950 6502 19962 6554
rect 20014 6502 21436 6554
rect 1104 6480 21436 6502
rect 5166 6440 5172 6452
rect 5127 6412 5172 6440
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7926 6440 7932 6452
rect 7887 6412 7932 6440
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6440 10474 6452
rect 10919 6443 10977 6449
rect 10919 6440 10931 6443
rect 10468 6412 10931 6440
rect 10468 6400 10474 6412
rect 10919 6409 10931 6412
rect 10965 6409 10977 6443
rect 10919 6403 10977 6409
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12897 6443 12955 6449
rect 12897 6440 12909 6443
rect 12124 6412 12909 6440
rect 12124 6400 12130 6412
rect 12897 6409 12909 6412
rect 12943 6440 12955 6443
rect 14001 6443 14059 6449
rect 12943 6412 13216 6440
rect 12943 6409 12955 6412
rect 12897 6403 12955 6409
rect 13188 6313 13216 6412
rect 14001 6409 14013 6443
rect 14047 6440 14059 6443
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 14047 6412 14197 6440
rect 14047 6409 14059 6412
rect 14001 6403 14059 6409
rect 14185 6409 14197 6412
rect 14231 6440 14243 6443
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 14231 6412 17325 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 17313 6409 17325 6412
rect 17359 6440 17371 6443
rect 17402 6440 17408 6452
rect 17359 6412 17408 6440
rect 17359 6409 17371 6412
rect 17313 6403 17371 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17770 6400 17776 6412
rect 17828 6440 17834 6452
rect 17828 6412 18368 6440
rect 17828 6400 17834 6412
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 14783 6276 14933 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 14921 6273 14933 6276
rect 14967 6304 14979 6307
rect 15286 6304 15292 6316
rect 14967 6276 15292 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 18340 6313 18368 6412
rect 18325 6307 18383 6313
rect 15436 6276 15481 6304
rect 15436 6264 15442 6276
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 10848 6239 10906 6245
rect 10848 6205 10860 6239
rect 10894 6236 10906 6239
rect 16460 6239 16518 6245
rect 10894 6208 11376 6236
rect 10894 6205 10906 6208
rect 10848 6199 10906 6205
rect 11348 6109 11376 6208
rect 16460 6205 16472 6239
rect 16506 6236 16518 6239
rect 16942 6236 16948 6248
rect 16506 6208 16948 6236
rect 16506 6205 16518 6208
rect 16460 6199 16518 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 13817 6171 13875 6177
rect 13817 6137 13829 6171
rect 13863 6168 13875 6171
rect 14182 6168 14188 6180
rect 13863 6140 14188 6168
rect 13863 6137 13875 6140
rect 13817 6131 13875 6137
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 18969 6171 19027 6177
rect 18969 6137 18981 6171
rect 19015 6137 19027 6171
rect 18969 6131 19027 6137
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11422 6100 11428 6112
rect 11379 6072 11428 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12894 6060 12900 6112
rect 12952 6100 12958 6112
rect 13446 6100 13452 6112
rect 12952 6072 13452 6100
rect 12952 6060 12958 6072
rect 13446 6060 13452 6072
rect 13504 6100 13510 6112
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13504 6072 14013 6100
rect 13504 6060 13510 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 16531 6103 16589 6109
rect 16531 6100 16543 6103
rect 15528 6072 16543 6100
rect 15528 6060 15534 6072
rect 16531 6069 16543 6072
rect 16577 6069 16589 6103
rect 18984 6100 19012 6131
rect 19242 6100 19248 6112
rect 18984 6072 19248 6100
rect 16531 6063 16589 6069
rect 19242 6060 19248 6072
rect 19300 6100 19306 6112
rect 19337 6103 19395 6109
rect 19337 6100 19349 6103
rect 19300 6072 19349 6100
rect 19300 6060 19306 6072
rect 19337 6069 19349 6072
rect 19383 6100 19395 6103
rect 19610 6100 19616 6112
rect 19383 6072 19616 6100
rect 19383 6069 19395 6072
rect 19337 6063 19395 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 1104 6010 21436 6032
rect 1104 5958 8497 6010
rect 8549 5958 8561 6010
rect 8613 5958 8625 6010
rect 8677 5958 8689 6010
rect 8741 5958 16012 6010
rect 16064 5958 16076 6010
rect 16128 5958 16140 6010
rect 16192 5958 16204 6010
rect 16256 5958 21436 6010
rect 1104 5936 21436 5958
rect 11195 5899 11253 5905
rect 11195 5865 11207 5899
rect 11241 5896 11253 5899
rect 11882 5896 11888 5908
rect 11241 5868 11888 5896
rect 11241 5865 11253 5868
rect 11195 5859 11253 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 17034 5896 17040 5908
rect 16995 5868 17040 5896
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 14323 5831 14381 5837
rect 14323 5797 14335 5831
rect 14369 5828 14381 5831
rect 14369 5800 16896 5828
rect 14369 5797 14381 5800
rect 14323 5791 14381 5797
rect 16868 5772 16896 5800
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 11054 5760 11060 5772
rect 11112 5769 11118 5772
rect 11112 5763 11150 5769
rect 10008 5732 11060 5760
rect 10008 5720 10014 5732
rect 11054 5720 11060 5732
rect 11138 5760 11150 5763
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11138 5732 12081 5760
rect 11138 5729 11150 5732
rect 11112 5723 11150 5729
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 11112 5720 11118 5723
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 13412 5732 14105 5760
rect 13412 5720 13418 5732
rect 14093 5729 14105 5732
rect 14139 5729 14151 5763
rect 16850 5760 16856 5772
rect 16763 5732 16856 5760
rect 14093 5723 14151 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 19334 5692 19340 5704
rect 19295 5664 19340 5692
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19610 5692 19616 5704
rect 19571 5664 19616 5692
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 14240 5596 15945 5624
rect 14240 5584 14246 5596
rect 15933 5593 15945 5596
rect 15979 5593 15991 5627
rect 15933 5587 15991 5593
rect 12253 5559 12311 5565
rect 12253 5525 12265 5559
rect 12299 5556 12311 5559
rect 13262 5556 13268 5568
rect 12299 5528 13268 5556
rect 12299 5525 12311 5528
rect 12253 5519 12311 5525
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 1104 5466 21436 5488
rect 1104 5414 4739 5466
rect 4791 5414 4803 5466
rect 4855 5414 4867 5466
rect 4919 5414 4931 5466
rect 4983 5414 12255 5466
rect 12307 5414 12319 5466
rect 12371 5414 12383 5466
rect 12435 5414 12447 5466
rect 12499 5414 19770 5466
rect 19822 5414 19834 5466
rect 19886 5414 19898 5466
rect 19950 5414 19962 5466
rect 20014 5414 21436 5466
rect 1104 5392 21436 5414
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5352 11118 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11112 5324 12081 5352
rect 11112 5312 11118 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 12069 5315 12127 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15378 5352 15384 5364
rect 14967 5324 15384 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 19334 5352 19340 5364
rect 19295 5324 19340 5352
rect 19334 5312 19340 5324
rect 19392 5352 19398 5364
rect 19751 5355 19809 5361
rect 19751 5352 19763 5355
rect 19392 5324 19763 5352
rect 19392 5312 19398 5324
rect 19751 5321 19763 5324
rect 19797 5321 19809 5355
rect 20162 5352 20168 5364
rect 20123 5324 20168 5352
rect 19751 5315 19809 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 15396 5284 15424 5312
rect 15396 5256 15792 5284
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15470 5216 15476 5228
rect 15335 5188 15476 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 15764 5225 15792 5256
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14312 5151 14370 5157
rect 14312 5148 14324 5151
rect 14240 5120 14324 5148
rect 14240 5108 14246 5120
rect 14312 5117 14324 5120
rect 14358 5117 14370 5151
rect 14312 5111 14370 5117
rect 19680 5151 19738 5157
rect 19680 5117 19692 5151
rect 19726 5148 19738 5151
rect 20162 5148 20168 5160
rect 19726 5120 20168 5148
rect 19726 5117 19738 5120
rect 19680 5111 19738 5117
rect 20162 5108 20168 5120
rect 20220 5108 20226 5160
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 13412 4984 13737 5012
rect 13412 4972 13418 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 13725 4975 13783 4981
rect 14415 5015 14473 5021
rect 14415 4981 14427 5015
rect 14461 5012 14473 5015
rect 14734 5012 14740 5024
rect 14461 4984 14740 5012
rect 14461 4981 14473 4984
rect 14415 4975 14473 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 1104 4922 21436 4944
rect 1104 4870 8497 4922
rect 8549 4870 8561 4922
rect 8613 4870 8625 4922
rect 8677 4870 8689 4922
rect 8741 4870 16012 4922
rect 16064 4870 16076 4922
rect 16128 4870 16140 4922
rect 16192 4870 16204 4922
rect 16256 4870 21436 4922
rect 1104 4848 21436 4870
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 13081 4743 13139 4749
rect 13081 4740 13093 4743
rect 12860 4712 13093 4740
rect 12860 4700 12866 4712
rect 13081 4709 13093 4712
rect 13127 4709 13139 4743
rect 13081 4703 13139 4709
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15286 4672 15292 4684
rect 14792 4644 15292 4672
rect 14792 4632 14798 4644
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 19426 4672 19432 4684
rect 19387 4644 19432 4672
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 17954 4604 17960 4616
rect 17915 4576 17960 4604
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 17310 4496 17316 4548
rect 17368 4536 17374 4548
rect 18248 4536 18276 4567
rect 17368 4508 18276 4536
rect 17368 4496 17374 4508
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15562 4468 15568 4480
rect 15519 4440 15568 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 18874 4428 18880 4480
rect 18932 4468 18938 4480
rect 19567 4471 19625 4477
rect 19567 4468 19579 4471
rect 18932 4440 19579 4468
rect 18932 4428 18938 4440
rect 19567 4437 19579 4440
rect 19613 4437 19625 4471
rect 19567 4431 19625 4437
rect 1104 4378 21436 4400
rect 1104 4326 4739 4378
rect 4791 4326 4803 4378
rect 4855 4326 4867 4378
rect 4919 4326 4931 4378
rect 4983 4326 12255 4378
rect 12307 4326 12319 4378
rect 12371 4326 12383 4378
rect 12435 4326 12447 4378
rect 12499 4326 19770 4378
rect 19822 4326 19834 4378
rect 19886 4326 19898 4378
rect 19950 4326 19962 4378
rect 20014 4326 21436 4378
rect 1104 4304 21436 4326
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5626 4264 5632 4276
rect 4488 4236 5632 4264
rect 4488 4224 4494 4236
rect 5626 4224 5632 4236
rect 5684 4264 5690 4276
rect 11790 4264 11796 4276
rect 5684 4236 11796 4264
rect 5684 4224 5690 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 12860 4236 13461 4264
rect 12860 4224 12866 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 15286 4264 15292 4276
rect 15247 4236 15292 4264
rect 13449 4227 13507 4233
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 18012 4236 18245 4264
rect 18012 4224 18018 4236
rect 18233 4233 18245 4236
rect 18279 4264 18291 4267
rect 18322 4264 18328 4276
rect 18279 4236 18328 4264
rect 18279 4233 18291 4236
rect 18233 4227 18291 4233
rect 18322 4224 18328 4236
rect 18380 4264 18386 4276
rect 19150 4264 19156 4276
rect 18380 4236 19156 4264
rect 18380 4224 18386 4236
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 19797 4267 19855 4273
rect 19797 4264 19809 4267
rect 19484 4236 19809 4264
rect 19484 4224 19490 4236
rect 19797 4233 19809 4236
rect 19843 4233 19855 4267
rect 19797 4227 19855 4233
rect 10413 4199 10471 4205
rect 10413 4165 10425 4199
rect 10459 4196 10471 4199
rect 17310 4196 17316 4208
rect 10459 4168 17316 4196
rect 10459 4165 10471 4168
rect 10413 4159 10471 4165
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 10520 4128 10548 4168
rect 17310 4156 17316 4168
rect 17368 4156 17374 4208
rect 9272 4100 10548 4128
rect 13173 4131 13231 4137
rect 9272 4088 9278 4100
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13354 4128 13360 4140
rect 13219 4100 13360 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 8824 4063 8882 4069
rect 8824 4029 8836 4063
rect 8870 4060 8882 4063
rect 8870 4032 9352 4060
rect 8870 4029 8882 4032
rect 8824 4023 8882 4029
rect 8895 3927 8953 3933
rect 8895 3893 8907 3927
rect 8941 3924 8953 3927
rect 9122 3924 9128 3936
rect 8941 3896 9128 3924
rect 8941 3893 8953 3896
rect 8895 3887 8953 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9324 3933 9352 4032
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 9861 3995 9919 4001
rect 9861 3992 9873 3995
rect 9723 3964 9873 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 9861 3961 9873 3964
rect 9907 3992 9919 3995
rect 10042 3992 10048 4004
rect 9907 3964 10048 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 12529 3995 12587 4001
rect 12529 3961 12541 3995
rect 12575 3961 12587 3995
rect 12529 3955 12587 3961
rect 18693 3995 18751 4001
rect 18693 3961 18705 3995
rect 18739 3992 18751 3995
rect 18874 3992 18880 4004
rect 18739 3964 18880 3992
rect 18739 3961 18751 3964
rect 18693 3955 18751 3961
rect 9309 3927 9367 3933
rect 9309 3893 9321 3927
rect 9355 3924 9367 3927
rect 9490 3924 9496 3936
rect 9355 3896 9496 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11664 3896 12173 3924
rect 11664 3884 11670 3896
rect 12161 3893 12173 3896
rect 12207 3924 12219 3927
rect 12544 3924 12572 3955
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 12207 3896 12572 3924
rect 16945 3927 17003 3933
rect 12207 3893 12219 3896
rect 12161 3887 12219 3893
rect 16945 3893 16957 3927
rect 16991 3924 17003 3927
rect 18230 3924 18236 3936
rect 16991 3896 18236 3924
rect 16991 3893 17003 3896
rect 16945 3887 17003 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 21436 3856
rect 1104 3782 8497 3834
rect 8549 3782 8561 3834
rect 8613 3782 8625 3834
rect 8677 3782 8689 3834
rect 8741 3782 16012 3834
rect 16064 3782 16076 3834
rect 16128 3782 16140 3834
rect 16192 3782 16204 3834
rect 16256 3782 21436 3834
rect 1104 3760 21436 3782
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8444 3692 8585 3720
rect 8444 3680 8450 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 9122 3612 9128 3664
rect 9180 3652 9186 3664
rect 9769 3655 9827 3661
rect 9769 3652 9781 3655
rect 9180 3624 9781 3652
rect 9180 3612 9186 3624
rect 9769 3621 9781 3624
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 16669 3655 16727 3661
rect 16669 3621 16681 3655
rect 16715 3652 16727 3655
rect 17126 3652 17132 3664
rect 16715 3624 17132 3652
rect 16715 3621 16727 3624
rect 16669 3615 16727 3621
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 17310 3652 17316 3664
rect 17271 3624 17316 3652
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 18230 3652 18236 3664
rect 18191 3624 18236 3652
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 10042 3516 10048 3528
rect 10003 3488 10048 3516
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11606 3516 11612 3528
rect 11567 3488 11612 3516
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18380 3488 18521 3516
rect 18380 3476 18386 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 1104 3290 21436 3312
rect 1104 3238 4739 3290
rect 4791 3238 4803 3290
rect 4855 3238 4867 3290
rect 4919 3238 4931 3290
rect 4983 3238 12255 3290
rect 12307 3238 12319 3290
rect 12371 3238 12383 3290
rect 12435 3238 12447 3290
rect 12499 3238 19770 3290
rect 19822 3238 19834 3290
rect 19886 3238 19898 3290
rect 19950 3238 19962 3290
rect 20014 3238 21436 3290
rect 1104 3216 21436 3238
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9180 3148 9413 3176
rect 9180 3136 9186 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 11330 3136 11336 3188
rect 11388 3136 11394 3188
rect 18230 3176 18236 3188
rect 18191 3148 18236 3176
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 8711 3111 8769 3117
rect 8711 3077 8723 3111
rect 8757 3108 8769 3111
rect 11348 3108 11376 3136
rect 11701 3111 11759 3117
rect 11701 3108 11713 3111
rect 8757 3080 11713 3108
rect 8757 3077 8769 3080
rect 8711 3071 8769 3077
rect 11701 3077 11713 3080
rect 11747 3077 11759 3111
rect 11701 3071 11759 3077
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11606 3040 11612 3052
rect 11379 3012 11612 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3040 17190 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17184 3012 17417 3040
rect 17184 3000 17190 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18380 3012 18797 3040
rect 18380 3000 18386 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8608 2975 8666 2981
rect 8608 2972 8620 2975
rect 8444 2944 8620 2972
rect 8444 2932 8450 2944
rect 8608 2941 8620 2944
rect 8654 2941 8666 2975
rect 8608 2935 8666 2941
rect 9636 2975 9694 2981
rect 9636 2941 9648 2975
rect 9682 2941 9694 2975
rect 9636 2935 9694 2941
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 8623 2836 8651 2935
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8527 2808 9137 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 9125 2805 9137 2808
rect 9171 2836 9183 2839
rect 9490 2836 9496 2848
rect 9171 2808 9496 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9651 2836 9679 2935
rect 9723 2907 9781 2913
rect 9723 2873 9735 2907
rect 9769 2904 9781 2907
rect 10413 2907 10471 2913
rect 10413 2904 10425 2907
rect 9769 2876 10425 2904
rect 9769 2873 9781 2876
rect 9723 2867 9781 2873
rect 10413 2873 10425 2876
rect 10459 2904 10471 2907
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10459 2876 10701 2904
rect 10459 2873 10471 2876
rect 10413 2867 10471 2873
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 16301 2907 16359 2913
rect 16301 2873 16313 2907
rect 16347 2904 16359 2907
rect 16485 2907 16543 2913
rect 16485 2904 16497 2907
rect 16347 2876 16497 2904
rect 16347 2873 16359 2876
rect 16301 2867 16359 2873
rect 16485 2873 16497 2876
rect 16531 2904 16543 2907
rect 16574 2904 16580 2916
rect 16531 2876 16580 2904
rect 16531 2873 16543 2876
rect 16485 2867 16543 2873
rect 16574 2864 16580 2876
rect 16632 2864 16638 2916
rect 17865 2907 17923 2913
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 17911 2876 18521 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 18509 2873 18521 2876
rect 18555 2904 18567 2907
rect 18598 2904 18604 2916
rect 18555 2876 18604 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 10137 2839 10195 2845
rect 10137 2836 10149 2839
rect 9651 2808 10149 2836
rect 10137 2805 10149 2808
rect 10183 2836 10195 2839
rect 10502 2836 10508 2848
rect 10183 2808 10508 2836
rect 10183 2805 10195 2808
rect 10137 2799 10195 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 1104 2746 21436 2768
rect 1104 2694 8497 2746
rect 8549 2694 8561 2746
rect 8613 2694 8625 2746
rect 8677 2694 8689 2746
rect 8741 2694 16012 2746
rect 16064 2694 16076 2746
rect 16128 2694 16140 2746
rect 16192 2694 16204 2746
rect 16256 2694 21436 2746
rect 1104 2672 21436 2694
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 16574 2632 16580 2644
rect 16535 2604 16580 2632
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 18598 2632 18604 2644
rect 18559 2604 18604 2632
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 9232 2564 9260 2592
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 8747 2536 9260 2564
rect 11440 2536 11989 2564
rect 8747 2505 8775 2536
rect 8716 2499 8775 2505
rect 8716 2465 8728 2499
rect 8762 2468 8775 2499
rect 8803 2499 8861 2505
rect 8762 2465 8774 2468
rect 8716 2459 8774 2465
rect 8803 2465 8815 2499
rect 8849 2496 8861 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8849 2468 9781 2496
rect 8849 2465 8861 2468
rect 8803 2459 8861 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9815 2468 10333 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11440 2505 11468 2536
rect 11977 2533 11989 2536
rect 12023 2564 12035 2567
rect 12802 2564 12808 2576
rect 12023 2536 12808 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11388 2468 11437 2496
rect 11388 2456 11394 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 11848 2468 12909 2496
rect 11848 2456 11854 2468
rect 12897 2465 12909 2468
rect 12943 2496 12955 2499
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 12943 2468 13461 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 16368 2499 16426 2505
rect 16368 2465 16380 2499
rect 16414 2496 16426 2499
rect 18392 2499 18450 2505
rect 16414 2468 16896 2496
rect 16414 2465 16426 2468
rect 16368 2459 16426 2465
rect 5442 2320 5448 2372
rect 5500 2360 5506 2372
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 5500 2332 9965 2360
rect 5500 2320 5506 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 9953 2323 10011 2329
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 12618 2360 12624 2372
rect 11655 2332 12624 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 13081 2363 13139 2369
rect 13081 2329 13093 2363
rect 13127 2360 13139 2363
rect 14642 2360 14648 2372
rect 13127 2332 14648 2360
rect 13127 2329 13139 2332
rect 13081 2323 13139 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 16868 2301 16896 2468
rect 18392 2465 18404 2499
rect 18438 2496 18450 2499
rect 18438 2468 18920 2496
rect 18438 2465 18450 2468
rect 18392 2459 18450 2465
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 16942 2292 16948 2304
rect 16899 2264 16948 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 18892 2301 18920 2468
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 18966 2292 18972 2304
rect 18923 2264 18972 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 18966 2252 18972 2264
rect 19024 2252 19030 2304
rect 1104 2202 21436 2224
rect 1104 2150 4739 2202
rect 4791 2150 4803 2202
rect 4855 2150 4867 2202
rect 4919 2150 4931 2202
rect 4983 2150 12255 2202
rect 12307 2150 12319 2202
rect 12371 2150 12383 2202
rect 12435 2150 12447 2202
rect 12499 2150 19770 2202
rect 19822 2150 19834 2202
rect 19886 2150 19898 2202
rect 19950 2150 19962 2202
rect 20014 2150 21436 2202
rect 1104 2128 21436 2150
rect 7282 76 7288 128
rect 7340 116 7346 128
rect 7926 116 7932 128
rect 7340 88 7932 116
rect 7340 76 7346 88
rect 7926 76 7932 88
rect 7984 76 7990 128
<< via1 >>
rect 4160 24216 4212 24268
rect 5264 24216 5316 24268
rect 8497 22278 8549 22330
rect 8561 22278 8613 22330
rect 8625 22278 8677 22330
rect 8689 22278 8741 22330
rect 16012 22278 16064 22330
rect 16076 22278 16128 22330
rect 16140 22278 16192 22330
rect 16204 22278 16256 22330
rect 112 22040 164 22092
rect 15844 22040 15896 22092
rect 19156 22040 19208 22092
rect 19616 22015 19668 22024
rect 19616 21981 19625 22015
rect 19625 21981 19659 22015
rect 19659 21981 19668 22015
rect 19616 21972 19668 21981
rect 20168 21947 20220 21956
rect 20168 21913 20177 21947
rect 20177 21913 20211 21947
rect 20211 21913 20220 21947
rect 20168 21904 20220 21913
rect 19340 21836 19392 21888
rect 4739 21734 4791 21786
rect 4803 21734 4855 21786
rect 4867 21734 4919 21786
rect 4931 21734 4983 21786
rect 12255 21734 12307 21786
rect 12319 21734 12371 21786
rect 12383 21734 12435 21786
rect 12447 21734 12499 21786
rect 19770 21734 19822 21786
rect 19834 21734 19886 21786
rect 19898 21734 19950 21786
rect 19962 21734 20014 21786
rect 18512 21632 18564 21684
rect 19156 21675 19208 21684
rect 19156 21641 19165 21675
rect 19165 21641 19199 21675
rect 19199 21641 19208 21675
rect 19156 21632 19208 21641
rect 19524 21675 19576 21684
rect 19524 21641 19533 21675
rect 19533 21641 19567 21675
rect 19567 21641 19576 21675
rect 19524 21632 19576 21641
rect 19340 21496 19392 21548
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 19524 21428 19576 21480
rect 18604 21292 18656 21344
rect 19432 21292 19484 21344
rect 8497 21190 8549 21242
rect 8561 21190 8613 21242
rect 8625 21190 8677 21242
rect 8689 21190 8741 21242
rect 16012 21190 16064 21242
rect 16076 21190 16128 21242
rect 16140 21190 16192 21242
rect 16204 21190 16256 21242
rect 8116 21131 8168 21140
rect 8116 21097 8125 21131
rect 8125 21097 8159 21131
rect 8159 21097 8168 21131
rect 8116 21088 8168 21097
rect 19340 21088 19392 21140
rect 18604 21063 18656 21072
rect 18604 21029 18613 21063
rect 18613 21029 18647 21063
rect 18647 21029 18656 21063
rect 18604 21020 18656 21029
rect 1308 20952 1360 21004
rect 5264 20952 5316 21004
rect 6460 20952 6512 21004
rect 7932 20995 7984 21004
rect 7932 20961 7941 20995
rect 7941 20961 7975 20995
rect 7975 20961 7984 20995
rect 7932 20952 7984 20961
rect 15844 20952 15896 21004
rect 17776 20884 17828 20936
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 20260 20816 20312 20868
rect 1952 20748 2004 20800
rect 5080 20748 5132 20800
rect 17500 20748 17552 20800
rect 19616 20748 19668 20800
rect 4739 20646 4791 20698
rect 4803 20646 4855 20698
rect 4867 20646 4919 20698
rect 4931 20646 4983 20698
rect 12255 20646 12307 20698
rect 12319 20646 12371 20698
rect 12383 20646 12435 20698
rect 12447 20646 12499 20698
rect 19770 20646 19822 20698
rect 19834 20646 19886 20698
rect 19898 20646 19950 20698
rect 19962 20646 20014 20698
rect 1308 20544 1360 20596
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 7932 20587 7984 20596
rect 7932 20553 7941 20587
rect 7941 20553 7975 20587
rect 7975 20553 7984 20587
rect 7932 20544 7984 20553
rect 15844 20544 15896 20596
rect 17500 20544 17552 20596
rect 17776 20587 17828 20596
rect 17776 20553 17785 20587
rect 17785 20553 17819 20587
rect 17819 20553 17828 20587
rect 17776 20544 17828 20553
rect 18604 20544 18656 20596
rect 3884 20408 3936 20460
rect 9404 20408 9456 20460
rect 17592 20408 17644 20460
rect 21364 20476 21416 20528
rect 7380 20272 7432 20324
rect 13176 20315 13228 20324
rect 13176 20281 13185 20315
rect 13185 20281 13219 20315
rect 13219 20281 13228 20315
rect 13176 20272 13228 20281
rect 19616 20315 19668 20324
rect 19616 20281 19625 20315
rect 19625 20281 19659 20315
rect 19659 20281 19668 20315
rect 19616 20272 19668 20281
rect 20260 20315 20312 20324
rect 20260 20281 20269 20315
rect 20269 20281 20303 20315
rect 20303 20281 20312 20315
rect 20260 20272 20312 20281
rect 8497 20102 8549 20154
rect 8561 20102 8613 20154
rect 8625 20102 8677 20154
rect 8689 20102 8741 20154
rect 16012 20102 16064 20154
rect 16076 20102 16128 20154
rect 16140 20102 16192 20154
rect 16204 20102 16256 20154
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 5080 19932 5132 19984
rect 13176 19932 13228 19984
rect 18880 19975 18932 19984
rect 18880 19941 18889 19975
rect 18889 19941 18923 19975
rect 18923 19941 18932 19975
rect 18880 19932 18932 19941
rect 19524 19864 19576 19916
rect 3792 19796 3844 19848
rect 5080 19839 5132 19848
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 19340 19660 19392 19712
rect 4739 19558 4791 19610
rect 4803 19558 4855 19610
rect 4867 19558 4919 19610
rect 4931 19558 4983 19610
rect 12255 19558 12307 19610
rect 12319 19558 12371 19610
rect 12383 19558 12435 19610
rect 12447 19558 12499 19610
rect 19770 19558 19822 19610
rect 19834 19558 19886 19610
rect 19898 19558 19950 19610
rect 19962 19558 20014 19610
rect 3792 19499 3844 19508
rect 3792 19465 3801 19499
rect 3801 19465 3835 19499
rect 3835 19465 3844 19499
rect 3792 19456 3844 19465
rect 5172 19456 5224 19508
rect 3976 19388 4028 19440
rect 5080 19320 5132 19372
rect 13360 19456 13412 19508
rect 18236 19499 18288 19508
rect 18236 19465 18245 19499
rect 18245 19465 18279 19499
rect 18279 19465 18288 19499
rect 18236 19456 18288 19465
rect 18972 19499 19024 19508
rect 18972 19465 18981 19499
rect 18981 19465 19015 19499
rect 19015 19465 19024 19499
rect 18972 19456 19024 19465
rect 19524 19499 19576 19508
rect 19524 19465 19533 19499
rect 19533 19465 19567 19499
rect 19567 19465 19576 19499
rect 19524 19456 19576 19465
rect 19432 19320 19484 19372
rect 18972 19252 19024 19304
rect 19432 19184 19484 19236
rect 20076 19184 20128 19236
rect 8497 19014 8549 19066
rect 8561 19014 8613 19066
rect 8625 19014 8677 19066
rect 8689 19014 8741 19066
rect 16012 19014 16064 19066
rect 16076 19014 16128 19066
rect 16140 19014 16192 19066
rect 16204 19014 16256 19066
rect 112 18912 164 18964
rect 4068 18912 4120 18964
rect 19524 18912 19576 18964
rect 20352 18912 20404 18964
rect 19340 18887 19392 18896
rect 19340 18853 19349 18887
rect 19349 18853 19383 18887
rect 19383 18853 19392 18887
rect 19340 18844 19392 18853
rect 2412 18776 2464 18828
rect 3792 18708 3844 18760
rect 19616 18751 19668 18760
rect 19616 18717 19625 18751
rect 19625 18717 19659 18751
rect 19659 18717 19668 18751
rect 19616 18708 19668 18717
rect 4739 18470 4791 18522
rect 4803 18470 4855 18522
rect 4867 18470 4919 18522
rect 4931 18470 4983 18522
rect 12255 18470 12307 18522
rect 12319 18470 12371 18522
rect 12383 18470 12435 18522
rect 12447 18470 12499 18522
rect 19770 18470 19822 18522
rect 19834 18470 19886 18522
rect 19898 18470 19950 18522
rect 19962 18470 20014 18522
rect 4068 18368 4120 18420
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 3792 18343 3844 18352
rect 3792 18309 3801 18343
rect 3801 18309 3835 18343
rect 3835 18309 3844 18343
rect 3792 18300 3844 18309
rect 3976 18232 4028 18284
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 8497 17926 8549 17978
rect 8561 17926 8613 17978
rect 8625 17926 8677 17978
rect 8689 17926 8741 17978
rect 16012 17926 16064 17978
rect 16076 17926 16128 17978
rect 16140 17926 16192 17978
rect 16204 17926 16256 17978
rect 2412 17824 2464 17876
rect 2964 17731 3016 17740
rect 2964 17697 2982 17731
rect 2982 17697 3016 17731
rect 2964 17688 3016 17697
rect 3792 17688 3844 17740
rect 8392 17688 8444 17740
rect 7380 17484 7432 17536
rect 4739 17382 4791 17434
rect 4803 17382 4855 17434
rect 4867 17382 4919 17434
rect 4931 17382 4983 17434
rect 12255 17382 12307 17434
rect 12319 17382 12371 17434
rect 12383 17382 12435 17434
rect 12447 17382 12499 17434
rect 19770 17382 19822 17434
rect 19834 17382 19886 17434
rect 19898 17382 19950 17434
rect 19962 17382 20014 17434
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 7656 17187 7708 17196
rect 7656 17153 7665 17187
rect 7665 17153 7699 17187
rect 7699 17153 7708 17187
rect 7656 17144 7708 17153
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 2780 17076 2832 17128
rect 4068 17076 4120 17128
rect 6092 16940 6144 16992
rect 8497 16838 8549 16890
rect 8561 16838 8613 16890
rect 8625 16838 8677 16890
rect 8689 16838 8741 16890
rect 16012 16838 16064 16890
rect 16076 16838 16128 16890
rect 16140 16838 16192 16890
rect 16204 16838 16256 16890
rect 6092 16711 6144 16720
rect 6092 16677 6101 16711
rect 6101 16677 6135 16711
rect 6135 16677 6144 16711
rect 6092 16668 6144 16677
rect 7656 16668 7708 16720
rect 4068 16600 4120 16652
rect 4436 16643 4488 16652
rect 4436 16609 4480 16643
rect 4480 16609 4488 16643
rect 4436 16600 4488 16609
rect 11152 16600 11204 16652
rect 4620 16396 4672 16448
rect 11980 16396 12032 16448
rect 4739 16294 4791 16346
rect 4803 16294 4855 16346
rect 4867 16294 4919 16346
rect 4931 16294 4983 16346
rect 12255 16294 12307 16346
rect 12319 16294 12371 16346
rect 12383 16294 12435 16346
rect 12447 16294 12499 16346
rect 19770 16294 19822 16346
rect 19834 16294 19886 16346
rect 19898 16294 19950 16346
rect 19962 16294 20014 16346
rect 4436 16235 4488 16244
rect 4436 16201 4445 16235
rect 4445 16201 4479 16235
rect 4479 16201 4488 16235
rect 4436 16192 4488 16201
rect 6092 16235 6144 16244
rect 6092 16201 6101 16235
rect 6101 16201 6135 16235
rect 6135 16201 6144 16235
rect 6092 16192 6144 16201
rect 11152 16192 11204 16244
rect 4620 16056 4672 16108
rect 11152 15988 11204 16040
rect 5540 15963 5592 15972
rect 5540 15929 5549 15963
rect 5549 15929 5583 15963
rect 5583 15929 5592 15963
rect 5540 15920 5592 15929
rect 11244 15852 11296 15904
rect 8497 15750 8549 15802
rect 8561 15750 8613 15802
rect 8625 15750 8677 15802
rect 8689 15750 8741 15802
rect 16012 15750 16064 15802
rect 16076 15750 16128 15802
rect 16140 15750 16192 15802
rect 16204 15750 16256 15802
rect 15476 15691 15528 15700
rect 15476 15657 15485 15691
rect 15485 15657 15519 15691
rect 15519 15657 15528 15691
rect 15476 15648 15528 15657
rect 5540 15623 5592 15632
rect 5540 15589 5549 15623
rect 5549 15589 5583 15623
rect 5583 15589 5592 15623
rect 5540 15580 5592 15589
rect 11244 15580 11296 15632
rect 9864 15512 9916 15564
rect 12900 15512 12952 15564
rect 14464 15512 14516 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 5080 15444 5132 15496
rect 3884 15376 3936 15428
rect 12072 15419 12124 15428
rect 12072 15385 12081 15419
rect 12081 15385 12115 15419
rect 12115 15385 12124 15419
rect 12072 15376 12124 15385
rect 11428 15308 11480 15360
rect 15476 15308 15528 15360
rect 4739 15206 4791 15258
rect 4803 15206 4855 15258
rect 4867 15206 4919 15258
rect 4931 15206 4983 15258
rect 12255 15206 12307 15258
rect 12319 15206 12371 15258
rect 12383 15206 12435 15258
rect 12447 15206 12499 15258
rect 19770 15206 19822 15258
rect 19834 15206 19886 15258
rect 19898 15206 19950 15258
rect 19962 15206 20014 15258
rect 5080 15147 5132 15156
rect 5080 15113 5089 15147
rect 5089 15113 5123 15147
rect 5123 15113 5132 15147
rect 5080 15104 5132 15113
rect 9864 15104 9916 15156
rect 11244 15104 11296 15156
rect 11980 15104 12032 15156
rect 17500 15147 17552 15156
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 4620 14943 4672 14952
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 4620 14900 4672 14909
rect 5908 14900 5960 14952
rect 7380 14900 7432 14952
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 15292 15036 15344 15088
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 5264 14875 5316 14884
rect 5264 14841 5273 14875
rect 5273 14841 5307 14875
rect 5307 14841 5316 14875
rect 5264 14832 5316 14841
rect 10876 14875 10928 14884
rect 10876 14841 10885 14875
rect 10885 14841 10919 14875
rect 10919 14841 10928 14875
rect 10876 14832 10928 14841
rect 12992 14832 13044 14884
rect 16856 14900 16908 14952
rect 17500 14900 17552 14952
rect 6828 14764 6880 14816
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 14004 14764 14056 14816
rect 15384 14764 15436 14816
rect 17224 14764 17276 14816
rect 8497 14662 8549 14714
rect 8561 14662 8613 14714
rect 8625 14662 8677 14714
rect 8689 14662 8741 14714
rect 16012 14662 16064 14714
rect 16076 14662 16128 14714
rect 16140 14662 16192 14714
rect 16204 14662 16256 14714
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 6828 14535 6880 14544
rect 6828 14501 6837 14535
rect 6837 14501 6871 14535
rect 6871 14501 6880 14535
rect 6828 14492 6880 14501
rect 7656 14492 7708 14544
rect 11428 14535 11480 14544
rect 11428 14501 11437 14535
rect 11437 14501 11471 14535
rect 11471 14501 11480 14535
rect 11428 14492 11480 14501
rect 12072 14535 12124 14544
rect 12072 14501 12081 14535
rect 12081 14501 12115 14535
rect 12115 14501 12124 14535
rect 12072 14492 12124 14501
rect 12992 14535 13044 14544
rect 12992 14501 13001 14535
rect 13001 14501 13035 14535
rect 13035 14501 13044 14535
rect 12992 14492 13044 14501
rect 15476 14535 15528 14544
rect 15476 14501 15485 14535
rect 15485 14501 15519 14535
rect 15519 14501 15528 14535
rect 15476 14492 15528 14501
rect 17224 14535 17276 14544
rect 17224 14501 17233 14535
rect 17233 14501 17267 14535
rect 17267 14501 17276 14535
rect 17224 14492 17276 14501
rect 1952 14424 2004 14476
rect 4620 14424 4672 14476
rect 5908 14424 5960 14476
rect 9312 14424 9364 14476
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 17960 14356 18012 14408
rect 5448 14288 5500 14340
rect 17132 14288 17184 14340
rect 1400 14220 1452 14272
rect 10140 14220 10192 14272
rect 4739 14118 4791 14170
rect 4803 14118 4855 14170
rect 4867 14118 4919 14170
rect 4931 14118 4983 14170
rect 12255 14118 12307 14170
rect 12319 14118 12371 14170
rect 12383 14118 12435 14170
rect 12447 14118 12499 14170
rect 19770 14118 19822 14170
rect 19834 14118 19886 14170
rect 19898 14118 19950 14170
rect 19962 14118 20014 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 4620 14016 4672 14068
rect 5908 14016 5960 14068
rect 6828 14016 6880 14068
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 11428 14059 11480 14068
rect 10140 14016 10192 14025
rect 3884 13880 3936 13932
rect 4344 13880 4396 13932
rect 7656 13948 7708 14000
rect 9404 13991 9456 14000
rect 9404 13957 9413 13991
rect 9413 13957 9447 13991
rect 9447 13957 9456 13991
rect 9404 13948 9456 13957
rect 9680 13948 9732 14000
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 15476 14059 15528 14068
rect 14004 14016 14056 14025
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 3516 13812 3568 13864
rect 4528 13744 4580 13796
rect 4712 13787 4764 13796
rect 4712 13753 4721 13787
rect 4721 13753 4755 13787
rect 4755 13753 4764 13787
rect 4712 13744 4764 13753
rect 7748 13787 7800 13796
rect 7748 13753 7757 13787
rect 7757 13753 7791 13787
rect 7791 13753 7800 13787
rect 7748 13744 7800 13753
rect 8392 13676 8444 13728
rect 9680 13744 9732 13796
rect 9404 13676 9456 13728
rect 13912 13744 13964 13796
rect 15476 14025 15485 14059
rect 15485 14025 15519 14059
rect 15519 14025 15528 14059
rect 15476 14016 15528 14025
rect 17224 14016 17276 14068
rect 16212 13880 16264 13932
rect 17960 13880 18012 13932
rect 16212 13744 16264 13796
rect 16488 13787 16540 13796
rect 16488 13753 16497 13787
rect 16497 13753 16531 13787
rect 16531 13753 16540 13787
rect 16488 13744 16540 13753
rect 17132 13787 17184 13796
rect 17132 13753 17141 13787
rect 17141 13753 17175 13787
rect 17175 13753 17184 13787
rect 17132 13744 17184 13753
rect 13268 13676 13320 13728
rect 8497 13574 8549 13626
rect 8561 13574 8613 13626
rect 8625 13574 8677 13626
rect 8689 13574 8741 13626
rect 16012 13574 16064 13626
rect 16076 13574 16128 13626
rect 16140 13574 16192 13626
rect 16204 13574 16256 13626
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 4712 13515 4764 13524
rect 4712 13481 4721 13515
rect 4721 13481 4755 13515
rect 4755 13481 4764 13515
rect 4712 13472 4764 13481
rect 5080 13472 5132 13524
rect 13820 13472 13872 13524
rect 13912 13472 13964 13524
rect 16488 13472 16540 13524
rect 17960 13447 18012 13456
rect 17960 13413 17969 13447
rect 17969 13413 18003 13447
rect 18003 13413 18012 13447
rect 17960 13404 18012 13413
rect 2504 13336 2556 13388
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 12992 13336 13044 13388
rect 15476 13336 15528 13388
rect 16856 13336 16908 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 7104 13268 7156 13320
rect 7748 13268 7800 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 11704 13311 11756 13320
rect 8392 13200 8444 13252
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 11888 13268 11940 13320
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 3332 13132 3384 13184
rect 4739 13030 4791 13082
rect 4803 13030 4855 13082
rect 4867 13030 4919 13082
rect 4931 13030 4983 13082
rect 12255 13030 12307 13082
rect 12319 13030 12371 13082
rect 12383 13030 12435 13082
rect 12447 13030 12499 13082
rect 19770 13030 19822 13082
rect 19834 13030 19886 13082
rect 19898 13030 19950 13082
rect 19962 13030 20014 13082
rect 4344 12971 4396 12980
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 4528 12928 4580 12980
rect 4068 12860 4120 12912
rect 5448 12928 5500 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17960 12928 18012 12980
rect 21088 12928 21140 12980
rect 7104 12792 7156 12844
rect 7564 12792 7616 12844
rect 112 12724 164 12776
rect 4344 12724 4396 12776
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 22100 12860 22152 12912
rect 11704 12792 11756 12844
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 15384 12792 15436 12844
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 19616 12724 19668 12776
rect 7104 12699 7156 12708
rect 7104 12665 7113 12699
rect 7113 12665 7147 12699
rect 7147 12665 7156 12699
rect 7104 12656 7156 12665
rect 7748 12699 7800 12708
rect 7748 12665 7757 12699
rect 7757 12665 7791 12699
rect 7791 12665 7800 12699
rect 7748 12656 7800 12665
rect 8208 12656 8260 12708
rect 18420 12656 18472 12708
rect 2228 12588 2280 12640
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 4160 12588 4212 12640
rect 7840 12588 7892 12640
rect 9312 12588 9364 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 15476 12588 15528 12640
rect 18052 12588 18104 12640
rect 8497 12486 8549 12538
rect 8561 12486 8613 12538
rect 8625 12486 8677 12538
rect 8689 12486 8741 12538
rect 16012 12486 16064 12538
rect 16076 12486 16128 12538
rect 16140 12486 16192 12538
rect 16204 12486 16256 12538
rect 1400 12316 1452 12368
rect 9312 12316 9364 12368
rect 9772 12359 9824 12368
rect 9772 12325 9781 12359
rect 9781 12325 9815 12359
rect 9815 12325 9824 12359
rect 9772 12316 9824 12325
rect 11888 12316 11940 12368
rect 12900 12359 12952 12368
rect 12900 12325 12909 12359
rect 12909 12325 12943 12359
rect 12943 12325 12952 12359
rect 12900 12316 12952 12325
rect 8208 12248 8260 12300
rect 20720 12248 20772 12300
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 13636 12180 13688 12232
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 18604 12223 18656 12232
rect 18604 12189 18613 12223
rect 18613 12189 18647 12223
rect 18647 12189 18656 12223
rect 18604 12180 18656 12189
rect 7104 12044 7156 12096
rect 20076 12044 20128 12096
rect 4739 11942 4791 11994
rect 4803 11942 4855 11994
rect 4867 11942 4919 11994
rect 4931 11942 4983 11994
rect 12255 11942 12307 11994
rect 12319 11942 12371 11994
rect 12383 11942 12435 11994
rect 12447 11942 12499 11994
rect 19770 11942 19822 11994
rect 19834 11942 19886 11994
rect 19898 11942 19950 11994
rect 19962 11942 20014 11994
rect 1400 11840 1452 11892
rect 4620 11840 4672 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 9772 11883 9824 11892
rect 9772 11849 9781 11883
rect 9781 11849 9815 11883
rect 9815 11849 9824 11883
rect 9772 11840 9824 11849
rect 12992 11840 13044 11892
rect 19616 11840 19668 11892
rect 4160 11815 4212 11824
rect 4160 11781 4169 11815
rect 4169 11781 4203 11815
rect 4203 11781 4212 11815
rect 7840 11815 7892 11824
rect 4160 11772 4212 11781
rect 7840 11781 7849 11815
rect 7849 11781 7883 11815
rect 7883 11781 7892 11815
rect 7840 11772 7892 11781
rect 18328 11815 18380 11824
rect 18328 11781 18337 11815
rect 18337 11781 18371 11815
rect 18371 11781 18380 11815
rect 18328 11772 18380 11781
rect 20260 11772 20312 11824
rect 1952 11704 2004 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 14188 11704 14240 11756
rect 19248 11704 19300 11756
rect 4068 11636 4120 11688
rect 7288 11611 7340 11620
rect 7288 11577 7297 11611
rect 7297 11577 7331 11611
rect 7331 11577 7340 11611
rect 7288 11568 7340 11577
rect 12532 11568 12584 11620
rect 2412 11500 2464 11552
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 11796 11500 11848 11552
rect 13544 11568 13596 11620
rect 18604 11636 18656 11688
rect 19340 11611 19392 11620
rect 19340 11577 19349 11611
rect 19349 11577 19383 11611
rect 19383 11577 19392 11611
rect 19340 11568 19392 11577
rect 19616 11568 19668 11620
rect 20720 11500 20772 11552
rect 8497 11398 8549 11450
rect 8561 11398 8613 11450
rect 8625 11398 8677 11450
rect 8689 11398 8741 11450
rect 16012 11398 16064 11450
rect 16076 11398 16128 11450
rect 16140 11398 16192 11450
rect 16204 11398 16256 11450
rect 6644 11296 6696 11348
rect 7288 11296 7340 11348
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 2412 11271 2464 11280
rect 2412 11237 2421 11271
rect 2421 11237 2455 11271
rect 2455 11237 2464 11271
rect 2412 11228 2464 11237
rect 5080 11271 5132 11280
rect 5080 11237 5089 11271
rect 5089 11237 5123 11271
rect 5123 11237 5132 11271
rect 5080 11228 5132 11237
rect 11704 11228 11756 11280
rect 12532 11228 12584 11280
rect 12716 11228 12768 11280
rect 18420 11271 18472 11280
rect 18420 11237 18429 11271
rect 18429 11237 18463 11271
rect 18463 11237 18472 11271
rect 18420 11228 18472 11237
rect 20260 11228 20312 11280
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 8300 11160 8352 11212
rect 4436 11135 4488 11144
rect 1676 11024 1728 11076
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 19340 11135 19392 11144
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 19340 11092 19392 11101
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 18144 10956 18196 11008
rect 4739 10854 4791 10906
rect 4803 10854 4855 10906
rect 4867 10854 4919 10906
rect 4931 10854 4983 10906
rect 12255 10854 12307 10906
rect 12319 10854 12371 10906
rect 12383 10854 12435 10906
rect 12447 10854 12499 10906
rect 19770 10854 19822 10906
rect 19834 10854 19886 10906
rect 19898 10854 19950 10906
rect 19962 10854 20014 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 4436 10752 4488 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 17776 10795 17828 10804
rect 17776 10761 17785 10795
rect 17785 10761 17819 10795
rect 17819 10761 17828 10795
rect 17776 10752 17828 10761
rect 13544 10727 13596 10736
rect 13544 10693 13553 10727
rect 13553 10693 13587 10727
rect 13587 10693 13596 10727
rect 13544 10684 13596 10693
rect 19340 10684 19392 10736
rect 19616 10684 19668 10736
rect 11796 10616 11848 10668
rect 18144 10659 18196 10668
rect 18144 10625 18153 10659
rect 18153 10625 18187 10659
rect 18187 10625 18196 10659
rect 18144 10616 18196 10625
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 20076 10616 20128 10668
rect 5632 10548 5684 10600
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 4896 10480 4948 10532
rect 8392 10480 8444 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 8300 10455 8352 10464
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 12808 10480 12860 10532
rect 11796 10455 11848 10464
rect 10600 10412 10652 10421
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 17408 10591 17460 10600
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 21824 10412 21876 10464
rect 8497 10310 8549 10362
rect 8561 10310 8613 10362
rect 8625 10310 8677 10362
rect 8689 10310 8741 10362
rect 16012 10310 16064 10362
rect 16076 10310 16128 10362
rect 16140 10310 16192 10362
rect 16204 10310 16256 10362
rect 10600 10208 10652 10260
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 20168 10208 20220 10260
rect 2228 10183 2280 10192
rect 2228 10149 2237 10183
rect 2237 10149 2271 10183
rect 2271 10149 2280 10183
rect 2228 10140 2280 10149
rect 17408 10140 17460 10192
rect 10140 10072 10192 10124
rect 11704 10072 11756 10124
rect 14648 10072 14700 10124
rect 20168 10072 20220 10124
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 12624 10004 12676 10056
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 2780 9936 2832 9945
rect 18420 9979 18472 9988
rect 18420 9945 18429 9979
rect 18429 9945 18463 9979
rect 18463 9945 18472 9979
rect 18420 9936 18472 9945
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 4739 9766 4791 9818
rect 4803 9766 4855 9818
rect 4867 9766 4919 9818
rect 4931 9766 4983 9818
rect 12255 9766 12307 9818
rect 12319 9766 12371 9818
rect 12383 9766 12435 9818
rect 12447 9766 12499 9818
rect 19770 9766 19822 9818
rect 19834 9766 19886 9818
rect 19898 9766 19950 9818
rect 19962 9766 20014 9818
rect 2228 9664 2280 9716
rect 4160 9664 4212 9716
rect 5816 9664 5868 9716
rect 11796 9664 11848 9716
rect 15200 9664 15252 9716
rect 17868 9707 17920 9716
rect 17868 9673 17877 9707
rect 17877 9673 17911 9707
rect 17911 9673 17920 9707
rect 17868 9664 17920 9673
rect 19432 9664 19484 9716
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 2044 9596 2096 9648
rect 10048 9639 10100 9648
rect 10048 9605 10057 9639
rect 10057 9605 10091 9639
rect 10091 9605 10100 9639
rect 10048 9596 10100 9605
rect 2596 9528 2648 9580
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4620 9528 4672 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 2504 9460 2556 9469
rect 5724 9460 5776 9512
rect 10140 9528 10192 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13636 9528 13688 9580
rect 14464 9528 14516 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 12532 9435 12584 9444
rect 12532 9401 12541 9435
rect 12541 9401 12575 9435
rect 12575 9401 12584 9435
rect 12532 9392 12584 9401
rect 112 9324 164 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 3516 9324 3568 9376
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 11980 9324 12032 9376
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 8497 9222 8549 9274
rect 8561 9222 8613 9274
rect 8625 9222 8677 9274
rect 8689 9222 8741 9274
rect 16012 9222 16064 9274
rect 16076 9222 16128 9274
rect 16140 9222 16192 9274
rect 16204 9222 16256 9274
rect 1676 9120 1728 9172
rect 12532 9120 12584 9172
rect 12624 9120 12676 9172
rect 14004 9120 14056 9172
rect 20168 9120 20220 9172
rect 2504 9052 2556 9104
rect 1584 8984 1636 9036
rect 10968 8984 11020 9036
rect 18604 8984 18656 9036
rect 20260 8984 20312 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 4160 8959 4212 8968
rect 2780 8916 2832 8925
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4620 8959 4672 8968
rect 4160 8916 4212 8925
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 7840 8916 7892 8968
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 12900 8916 12952 8968
rect 7564 8848 7616 8900
rect 11980 8848 12032 8900
rect 17408 8848 17460 8900
rect 4739 8678 4791 8730
rect 4803 8678 4855 8730
rect 4867 8678 4919 8730
rect 4931 8678 4983 8730
rect 12255 8678 12307 8730
rect 12319 8678 12371 8730
rect 12383 8678 12435 8730
rect 12447 8678 12499 8730
rect 19770 8678 19822 8730
rect 19834 8678 19886 8730
rect 19898 8678 19950 8730
rect 19962 8678 20014 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2504 8576 2556 8628
rect 4160 8576 4212 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 19432 8576 19484 8628
rect 3976 8508 4028 8560
rect 20168 8508 20220 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 14464 8440 14516 8492
rect 19248 8440 19300 8492
rect 2596 8372 2648 8424
rect 7932 8372 7984 8424
rect 6920 8347 6972 8356
rect 6920 8313 6929 8347
rect 6929 8313 6963 8347
rect 6963 8313 6972 8347
rect 6920 8304 6972 8313
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 19064 8415 19116 8424
rect 19064 8381 19073 8415
rect 19073 8381 19107 8415
rect 19107 8381 19116 8415
rect 19064 8372 19116 8381
rect 19616 8415 19668 8424
rect 19616 8381 19625 8415
rect 19625 8381 19659 8415
rect 19659 8381 19668 8415
rect 19616 8372 19668 8381
rect 10968 8279 11020 8288
rect 10968 8245 10977 8279
rect 10977 8245 11011 8279
rect 11011 8245 11020 8279
rect 10968 8236 11020 8245
rect 11060 8236 11112 8288
rect 12072 8236 12124 8288
rect 14280 8236 14332 8288
rect 20260 8279 20312 8288
rect 20260 8245 20269 8279
rect 20269 8245 20303 8279
rect 20303 8245 20312 8279
rect 20260 8236 20312 8245
rect 8497 8134 8549 8186
rect 8561 8134 8613 8186
rect 8625 8134 8677 8186
rect 8689 8134 8741 8186
rect 16012 8134 16064 8186
rect 16076 8134 16128 8186
rect 16140 8134 16192 8186
rect 16204 8134 16256 8186
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 3608 8032 3660 8084
rect 3976 7964 4028 8016
rect 6920 8032 6972 8084
rect 19616 8032 19668 8084
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 10324 7939 10376 7948
rect 10324 7905 10368 7939
rect 10368 7905 10376 7939
rect 10324 7896 10376 7905
rect 19248 7896 19300 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 11520 7828 11572 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 13912 7828 13964 7880
rect 14280 7803 14332 7812
rect 14280 7769 14289 7803
rect 14289 7769 14323 7803
rect 14323 7769 14332 7803
rect 14280 7760 14332 7769
rect 6736 7692 6788 7744
rect 10784 7735 10836 7744
rect 10784 7701 10793 7735
rect 10793 7701 10827 7735
rect 10827 7701 10836 7735
rect 10784 7692 10836 7701
rect 4739 7590 4791 7642
rect 4803 7590 4855 7642
rect 4867 7590 4919 7642
rect 4931 7590 4983 7642
rect 12255 7590 12307 7642
rect 12319 7590 12371 7642
rect 12383 7590 12435 7642
rect 12447 7590 12499 7642
rect 19770 7590 19822 7642
rect 19834 7590 19886 7642
rect 19898 7590 19950 7642
rect 19962 7590 20014 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 4344 7488 4396 7540
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 10324 7531 10376 7540
rect 10324 7497 10333 7531
rect 10333 7497 10367 7531
rect 10367 7497 10376 7531
rect 10324 7488 10376 7497
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 13728 7488 13780 7540
rect 19248 7488 19300 7540
rect 13360 7463 13412 7472
rect 13360 7429 13369 7463
rect 13369 7429 13403 7463
rect 13403 7429 13412 7463
rect 13360 7420 13412 7429
rect 5172 7352 5224 7404
rect 6920 7352 6972 7404
rect 1308 7284 1360 7336
rect 4620 7284 4672 7336
rect 10784 7352 10836 7404
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 14280 7352 14332 7404
rect 19064 7352 19116 7404
rect 19524 7352 19576 7404
rect 5724 7148 5776 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 8497 7046 8549 7098
rect 8561 7046 8613 7098
rect 8625 7046 8677 7098
rect 8689 7046 8741 7098
rect 16012 7046 16064 7098
rect 16076 7046 16128 7098
rect 16140 7046 16192 7098
rect 16204 7046 16256 7098
rect 15200 6944 15252 6996
rect 11060 6919 11112 6928
rect 11060 6885 11069 6919
rect 11069 6885 11103 6919
rect 11103 6885 11112 6919
rect 11060 6876 11112 6885
rect 13728 6876 13780 6928
rect 5172 6851 5224 6860
rect 5172 6817 5181 6851
rect 5181 6817 5215 6851
rect 5215 6817 5224 6851
rect 5172 6808 5224 6817
rect 5724 6808 5776 6860
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 7932 6808 7984 6817
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 17408 6808 17460 6860
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 11888 6672 11940 6724
rect 12072 6740 12124 6792
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 6184 6604 6236 6656
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 8944 6604 8996 6656
rect 17776 6604 17828 6656
rect 4739 6502 4791 6554
rect 4803 6502 4855 6554
rect 4867 6502 4919 6554
rect 4931 6502 4983 6554
rect 12255 6502 12307 6554
rect 12319 6502 12371 6554
rect 12383 6502 12435 6554
rect 12447 6502 12499 6554
rect 19770 6502 19822 6554
rect 19834 6502 19886 6554
rect 19898 6502 19950 6554
rect 19962 6502 20014 6554
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 12072 6400 12124 6452
rect 17408 6400 17460 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 15292 6264 15344 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 14188 6128 14240 6180
rect 11428 6060 11480 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12900 6060 12952 6112
rect 13452 6060 13504 6112
rect 15476 6060 15528 6112
rect 19248 6060 19300 6112
rect 19616 6060 19668 6112
rect 8497 5958 8549 6010
rect 8561 5958 8613 6010
rect 8625 5958 8677 6010
rect 8689 5958 8741 6010
rect 16012 5958 16064 6010
rect 16076 5958 16128 6010
rect 16140 5958 16192 6010
rect 16204 5958 16256 6010
rect 11888 5856 11940 5908
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 9956 5720 10008 5772
rect 11060 5763 11112 5772
rect 11060 5729 11104 5763
rect 11104 5729 11112 5763
rect 11060 5720 11112 5729
rect 13360 5720 13412 5772
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 14188 5584 14240 5636
rect 13268 5516 13320 5568
rect 4739 5414 4791 5466
rect 4803 5414 4855 5466
rect 4867 5414 4919 5466
rect 4931 5414 4983 5466
rect 12255 5414 12307 5466
rect 12319 5414 12371 5466
rect 12383 5414 12435 5466
rect 12447 5414 12499 5466
rect 19770 5414 19822 5466
rect 19834 5414 19886 5466
rect 19898 5414 19950 5466
rect 19962 5414 20014 5466
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 15384 5312 15436 5364
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 19340 5312 19392 5321
rect 20168 5355 20220 5364
rect 20168 5321 20177 5355
rect 20177 5321 20211 5355
rect 20211 5321 20220 5355
rect 20168 5312 20220 5321
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 14188 5108 14240 5160
rect 20168 5108 20220 5160
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 13360 4972 13412 5024
rect 14740 4972 14792 5024
rect 8497 4870 8549 4922
rect 8561 4870 8613 4922
rect 8625 4870 8677 4922
rect 8689 4870 8741 4922
rect 16012 4870 16064 4922
rect 16076 4870 16128 4922
rect 16140 4870 16192 4922
rect 16204 4870 16256 4922
rect 12808 4700 12860 4752
rect 14740 4632 14792 4684
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 19432 4675 19484 4684
rect 19432 4641 19441 4675
rect 19441 4641 19475 4675
rect 19475 4641 19484 4675
rect 19432 4632 19484 4641
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 17316 4496 17368 4548
rect 15568 4428 15620 4480
rect 18880 4428 18932 4480
rect 4739 4326 4791 4378
rect 4803 4326 4855 4378
rect 4867 4326 4919 4378
rect 4931 4326 4983 4378
rect 12255 4326 12307 4378
rect 12319 4326 12371 4378
rect 12383 4326 12435 4378
rect 12447 4326 12499 4378
rect 19770 4326 19822 4378
rect 19834 4326 19886 4378
rect 19898 4326 19950 4378
rect 19962 4326 20014 4378
rect 4436 4224 4488 4276
rect 5632 4224 5684 4276
rect 11796 4224 11848 4276
rect 12808 4224 12860 4276
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 17960 4224 18012 4276
rect 18328 4224 18380 4276
rect 19156 4224 19208 4276
rect 19432 4224 19484 4276
rect 9220 4088 9272 4140
rect 17316 4156 17368 4208
rect 13360 4088 13412 4140
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 9128 3884 9180 3936
rect 10048 3952 10100 4004
rect 18880 3995 18932 4004
rect 9496 3884 9548 3936
rect 11612 3884 11664 3936
rect 18880 3961 18889 3995
rect 18889 3961 18923 3995
rect 18923 3961 18932 3995
rect 18880 3952 18932 3961
rect 18236 3884 18288 3936
rect 8497 3782 8549 3834
rect 8561 3782 8613 3834
rect 8625 3782 8677 3834
rect 8689 3782 8741 3834
rect 16012 3782 16064 3834
rect 16076 3782 16128 3834
rect 16140 3782 16192 3834
rect 16204 3782 16256 3834
rect 8392 3680 8444 3732
rect 9128 3612 9180 3664
rect 17132 3612 17184 3664
rect 17316 3655 17368 3664
rect 17316 3621 17325 3655
rect 17325 3621 17359 3655
rect 17359 3621 17368 3655
rect 17316 3612 17368 3621
rect 18236 3655 18288 3664
rect 18236 3621 18245 3655
rect 18245 3621 18279 3655
rect 18279 3621 18288 3655
rect 18236 3612 18288 3621
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 18328 3476 18380 3528
rect 4739 3238 4791 3290
rect 4803 3238 4855 3290
rect 4867 3238 4919 3290
rect 4931 3238 4983 3290
rect 12255 3238 12307 3290
rect 12319 3238 12371 3290
rect 12383 3238 12435 3290
rect 12447 3238 12499 3290
rect 19770 3238 19822 3290
rect 19834 3238 19886 3290
rect 19898 3238 19950 3290
rect 19962 3238 20014 3290
rect 9128 3136 9180 3188
rect 11336 3136 11388 3188
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 11612 3000 11664 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 18328 3000 18380 3052
rect 8392 2932 8444 2984
rect 9496 2796 9548 2848
rect 16580 2864 16632 2916
rect 18604 2864 18656 2916
rect 10508 2796 10560 2848
rect 8497 2694 8549 2746
rect 8561 2694 8613 2746
rect 8625 2694 8677 2746
rect 8689 2694 8741 2746
rect 16012 2694 16064 2746
rect 16076 2694 16128 2746
rect 16140 2694 16192 2746
rect 16204 2694 16256 2746
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 16580 2635 16632 2644
rect 16580 2601 16589 2635
rect 16589 2601 16623 2635
rect 16623 2601 16632 2635
rect 16580 2592 16632 2601
rect 18604 2635 18656 2644
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 18604 2592 18656 2601
rect 11336 2456 11388 2508
rect 12808 2524 12860 2576
rect 11796 2456 11848 2508
rect 5448 2320 5500 2372
rect 12624 2320 12676 2372
rect 14648 2320 14700 2372
rect 16948 2252 17000 2304
rect 18972 2252 19024 2304
rect 4739 2150 4791 2202
rect 4803 2150 4855 2202
rect 4867 2150 4919 2202
rect 4931 2150 4983 2202
rect 12255 2150 12307 2202
rect 12319 2150 12371 2202
rect 12383 2150 12435 2202
rect 12447 2150 12499 2202
rect 19770 2150 19822 2202
rect 19834 2150 19886 2202
rect 19898 2150 19950 2202
rect 19962 2150 20014 2202
rect 7288 76 7340 128
rect 7932 76 7984 128
<< metal2 >>
rect 754 24210 810 24690
rect 2226 24210 2282 24690
rect 3698 24290 3754 24690
rect 3620 24262 3754 24290
rect 1306 23488 1362 23497
rect 1306 23423 1362 23432
rect 110 22808 166 22817
rect 110 22743 166 22752
rect 124 22098 152 22743
rect 112 22092 164 22098
rect 112 22034 164 22040
rect 1320 21010 1348 23423
rect 3514 21040 3570 21049
rect 1308 21004 1360 21010
rect 3514 20975 3570 20984
rect 1308 20946 1360 20952
rect 1320 20602 1348 20946
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1964 20602 1992 20742
rect 1308 20596 1360 20602
rect 1308 20538 1360 20544
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 110 19136 166 19145
rect 110 19071 166 19080
rect 124 18970 152 19071
rect 112 18964 164 18970
rect 112 18906 164 18912
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 13870 1440 14214
rect 1596 14074 1624 19751
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2424 18086 2452 18770
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2424 17882 2452 18022
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2778 17368 2834 17377
rect 2976 17338 3004 17682
rect 2778 17303 2834 17312
rect 2964 17332 3016 17338
rect 2792 17134 2820 17303
rect 2964 17274 3016 17280
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1964 14074 1992 14418
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 110 13016 166 13025
rect 110 12951 166 12960
rect 124 12782 152 12951
rect 112 12776 164 12782
rect 112 12718 164 12724
rect 1412 12374 1440 13262
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 1412 11898 1440 12310
rect 1964 12238 1992 14010
rect 3528 13870 3556 20975
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 12646 2544 13330
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1964 11762 1992 12174
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10470 1716 11018
rect 2044 10532 2096 10538
rect 2044 10474 2096 10480
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1412 9518 1440 9823
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 112 9376 164 9382
rect 112 9318 164 9324
rect 124 5545 152 9318
rect 1688 9178 1716 10406
rect 2056 9926 2084 10474
rect 2240 10198 2268 12582
rect 2516 11937 2544 12582
rect 2502 11928 2558 11937
rect 2502 11863 2558 11872
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11286 2452 11494
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2424 10674 2452 11222
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9654 2084 9862
rect 2240 9722 2268 10134
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2516 9518 2544 11863
rect 3344 10810 3372 13126
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2516 9110 2544 9454
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 8634 1624 8978
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8634 2544 8910
rect 2608 8673 2636 9522
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2594 8664 2650 8673
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 2504 8628 2556 8634
rect 2594 8599 2650 8608
rect 2504 8570 2556 8576
rect 2608 8430 2636 8599
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7546 2268 7822
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 1308 7336 1360 7342
rect 2700 7313 2728 9318
rect 2792 8974 2820 9930
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 8090 3372 8434
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 1308 7278 1360 7284
rect 2686 7304 2742 7313
rect 110 5536 166 5545
rect 110 5471 166 5480
rect 1320 2417 1348 7278
rect 2686 7239 2742 7248
rect 1306 2408 1362 2417
rect 1306 2343 1362 2352
rect 2226 1456 2282 1465
rect 2226 1391 2282 1400
rect 478 0 534 480
rect 1398 0 1454 480
rect 2240 82 2268 1391
rect 2318 82 2374 480
rect 2240 54 2374 82
rect 2318 0 2374 54
rect 3238 82 3294 480
rect 3528 82 3556 9318
rect 3620 8090 3648 24262
rect 3698 24210 3754 24262
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 5262 24268 5318 24690
rect 6734 24290 6790 24690
rect 8206 24290 8262 24690
rect 5262 24216 5264 24268
rect 5316 24216 5318 24268
rect 5262 24210 5318 24216
rect 6472 24262 6790 24290
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3804 19514 3832 19790
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3804 18358 3832 18702
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 3804 17746 3832 18294
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3896 15434 3924 20402
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 3988 18952 4016 19382
rect 4068 18964 4120 18970
rect 3988 18924 4068 18952
rect 4068 18906 4120 18912
rect 4080 18426 4108 18906
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3896 13938 3924 15370
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 10577 3924 11494
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3988 8566 4016 18226
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16658 4108 17070
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12918 4108 13330
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4172 12730 4200 24210
rect 5276 24179 5304 24210
rect 4713 21788 5009 21808
rect 4769 21786 4793 21788
rect 4849 21786 4873 21788
rect 4929 21786 4953 21788
rect 4791 21734 4793 21786
rect 4855 21734 4867 21786
rect 4929 21734 4931 21786
rect 4769 21732 4793 21734
rect 4849 21732 4873 21734
rect 4929 21732 4953 21734
rect 4713 21712 5009 21732
rect 6472 21010 6500 24262
rect 6734 24210 6790 24262
rect 8128 24262 8262 24290
rect 8128 21146 8156 24262
rect 8206 24210 8262 24262
rect 9770 24290 9826 24690
rect 11242 24290 11298 24690
rect 9770 24262 9904 24290
rect 9770 24210 9826 24262
rect 8471 22332 8767 22352
rect 8527 22330 8551 22332
rect 8607 22330 8631 22332
rect 8687 22330 8711 22332
rect 8549 22278 8551 22330
rect 8613 22278 8625 22330
rect 8687 22278 8689 22330
rect 8527 22276 8551 22278
rect 8607 22276 8631 22278
rect 8687 22276 8711 22278
rect 8471 22256 8767 22276
rect 8471 21244 8767 21264
rect 8527 21242 8551 21244
rect 8607 21242 8631 21244
rect 8687 21242 8711 21244
rect 8549 21190 8551 21242
rect 8613 21190 8625 21242
rect 8687 21190 8689 21242
rect 8527 21188 8551 21190
rect 8607 21188 8631 21190
rect 8687 21188 8711 21190
rect 8471 21168 8767 21188
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 7932 21004 7984 21010
rect 7932 20946 7984 20952
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4713 20700 5009 20720
rect 4769 20698 4793 20700
rect 4849 20698 4873 20700
rect 4929 20698 4953 20700
rect 4791 20646 4793 20698
rect 4855 20646 4867 20698
rect 4929 20646 4931 20698
rect 4769 20644 4793 20646
rect 4849 20644 4873 20646
rect 4929 20644 4953 20646
rect 4713 20624 5009 20644
rect 5092 19990 5120 20742
rect 5276 20602 5304 20946
rect 7944 20602 7972 20946
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 7380 20324 7432 20330
rect 7380 20266 7432 20272
rect 5080 19984 5132 19990
rect 5132 19944 5212 19972
rect 5080 19926 5132 19932
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 4713 19612 5009 19632
rect 4769 19610 4793 19612
rect 4849 19610 4873 19612
rect 4929 19610 4953 19612
rect 4791 19558 4793 19610
rect 4855 19558 4867 19610
rect 4929 19558 4931 19610
rect 4769 19556 4793 19558
rect 4849 19556 4873 19558
rect 4929 19556 4953 19558
rect 4713 19536 5009 19556
rect 5092 19378 5120 19790
rect 5184 19514 5212 19944
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 7392 19281 7420 20266
rect 8471 20156 8767 20176
rect 8527 20154 8551 20156
rect 8607 20154 8631 20156
rect 8687 20154 8711 20156
rect 8549 20102 8551 20154
rect 8613 20102 8625 20154
rect 8687 20102 8689 20154
rect 8527 20100 8551 20102
rect 8607 20100 8631 20102
rect 8687 20100 8711 20102
rect 8471 20080 8767 20100
rect 7378 19272 7434 19281
rect 7378 19207 7434 19216
rect 8471 19068 8767 19088
rect 8527 19066 8551 19068
rect 8607 19066 8631 19068
rect 8687 19066 8711 19068
rect 8549 19014 8551 19066
rect 8613 19014 8625 19066
rect 8687 19014 8689 19066
rect 8527 19012 8551 19014
rect 8607 19012 8631 19014
rect 8687 19012 8711 19014
rect 8471 18992 8767 19012
rect 4713 18524 5009 18544
rect 4769 18522 4793 18524
rect 4849 18522 4873 18524
rect 4929 18522 4953 18524
rect 4791 18470 4793 18522
rect 4855 18470 4867 18522
rect 4929 18470 4931 18522
rect 4769 18468 4793 18470
rect 4849 18468 4873 18470
rect 4929 18468 4953 18470
rect 4713 18448 5009 18468
rect 8471 17980 8767 18000
rect 8527 17978 8551 17980
rect 8607 17978 8631 17980
rect 8687 17978 8711 17980
rect 8549 17926 8551 17978
rect 8613 17926 8625 17978
rect 8687 17926 8689 17978
rect 8527 17924 8551 17926
rect 8607 17924 8631 17926
rect 8687 17924 8711 17926
rect 8471 17904 8767 17924
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 4713 17436 5009 17456
rect 4769 17434 4793 17436
rect 4849 17434 4873 17436
rect 4929 17434 4953 17436
rect 4791 17382 4793 17434
rect 4855 17382 4867 17434
rect 4929 17382 4931 17434
rect 4769 17380 4793 17382
rect 4849 17380 4873 17382
rect 4929 17380 4953 17382
rect 4713 17360 5009 17380
rect 7392 17202 7420 17478
rect 8404 17202 8432 17682
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16726 6132 16934
rect 7668 16726 7696 17138
rect 8404 17105 8432 17138
rect 8390 17096 8446 17105
rect 8390 17031 8446 17040
rect 8471 16892 8767 16912
rect 8527 16890 8551 16892
rect 8607 16890 8631 16892
rect 8687 16890 8711 16892
rect 8549 16838 8551 16890
rect 8613 16838 8625 16890
rect 8687 16838 8689 16890
rect 8527 16836 8551 16838
rect 8607 16836 8631 16838
rect 8687 16836 8711 16838
rect 8471 16816 8767 16836
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4448 16250 4476 16594
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4632 16114 4660 16390
rect 4713 16348 5009 16368
rect 4769 16346 4793 16348
rect 4849 16346 4873 16348
rect 4929 16346 4953 16348
rect 4791 16294 4793 16346
rect 4855 16294 4867 16346
rect 4929 16294 4931 16346
rect 4769 16292 4793 16294
rect 4849 16292 4873 16294
rect 4929 16292 4953 16294
rect 4713 16272 5009 16292
rect 6104 16250 6132 16662
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5552 15638 5580 15914
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 4713 15260 5009 15280
rect 4769 15258 4793 15260
rect 4849 15258 4873 15260
rect 4929 15258 4953 15260
rect 4791 15206 4793 15258
rect 4855 15206 4867 15258
rect 4929 15206 4931 15258
rect 4769 15204 4793 15206
rect 4849 15204 4873 15206
rect 4929 15204 4953 15206
rect 4713 15184 5009 15204
rect 5092 15162 5120 15438
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 4618 15056 4674 15065
rect 5552 15026 5580 15574
rect 4618 14991 4674 15000
rect 5540 15020 5592 15026
rect 4632 14958 4660 14991
rect 5540 14962 5592 14968
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 5908 14952 5960 14958
rect 7380 14952 7432 14958
rect 5908 14894 5960 14900
rect 7378 14920 7380 14929
rect 7432 14920 7434 14929
rect 4632 14482 4660 14894
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5276 14618 5304 14826
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5920 14482 5948 14894
rect 7378 14855 7434 14864
rect 7392 14822 7420 14855
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 6840 14550 6868 14758
rect 7668 14550 7696 16662
rect 9310 16144 9366 16153
rect 9310 16079 9366 16088
rect 8471 15804 8767 15824
rect 8527 15802 8551 15804
rect 8607 15802 8631 15804
rect 8687 15802 8711 15804
rect 8549 15750 8551 15802
rect 8613 15750 8625 15802
rect 8687 15750 8689 15802
rect 8527 15748 8551 15750
rect 8607 15748 8631 15750
rect 8687 15748 8711 15750
rect 8471 15728 8767 15748
rect 8471 14716 8767 14736
rect 8527 14714 8551 14716
rect 8607 14714 8631 14716
rect 8687 14714 8711 14716
rect 8549 14662 8551 14714
rect 8613 14662 8625 14714
rect 8687 14662 8689 14714
rect 8527 14660 8551 14662
rect 8607 14660 8631 14662
rect 8687 14660 8711 14662
rect 8471 14640 8767 14660
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 4632 14074 4660 14418
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 4713 14172 5009 14192
rect 4769 14170 4793 14172
rect 4849 14170 4873 14172
rect 4929 14170 4953 14172
rect 4791 14118 4793 14170
rect 4855 14118 4867 14170
rect 4929 14118 4931 14170
rect 4769 14116 4793 14118
rect 4849 14116 4873 14118
rect 4929 14116 4953 14118
rect 4713 14096 5009 14116
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 4264 13530 4292 13631
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4356 12986 4384 13874
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4540 12986 4568 13738
rect 4724 13530 4752 13738
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4713 13084 5009 13104
rect 4769 13082 4793 13084
rect 4849 13082 4873 13084
rect 4929 13082 4953 13084
rect 4791 13030 4793 13082
rect 4855 13030 4867 13082
rect 4929 13030 4931 13082
rect 4769 13028 4793 13030
rect 4849 13028 4873 13030
rect 4929 13028 4953 13030
rect 4713 13008 5009 13028
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4356 12782 4384 12922
rect 4080 12702 4200 12730
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4080 11694 4108 12702
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 11830 4200 12582
rect 5092 12238 5120 13466
rect 5460 13326 5488 14282
rect 5920 14074 5948 14418
rect 6840 14074 6868 14486
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 7668 14006 7696 14486
rect 9324 14482 9352 16079
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 9324 13814 9352 14418
rect 9416 14006 9444 20402
rect 9876 15570 9904 24262
rect 11164 24262 11298 24290
rect 11164 16658 11192 24262
rect 11242 24210 11298 24262
rect 12714 24290 12770 24690
rect 14278 24290 14334 24690
rect 15750 24290 15806 24690
rect 17222 24290 17278 24690
rect 18786 24290 18842 24690
rect 12714 24262 12940 24290
rect 12714 24210 12770 24262
rect 12229 21788 12525 21808
rect 12285 21786 12309 21788
rect 12365 21786 12389 21788
rect 12445 21786 12469 21788
rect 12307 21734 12309 21786
rect 12371 21734 12383 21786
rect 12445 21734 12447 21786
rect 12285 21732 12309 21734
rect 12365 21732 12389 21734
rect 12445 21732 12469 21734
rect 12229 21712 12525 21732
rect 12229 20700 12525 20720
rect 12285 20698 12309 20700
rect 12365 20698 12389 20700
rect 12445 20698 12469 20700
rect 12307 20646 12309 20698
rect 12371 20646 12383 20698
rect 12445 20646 12447 20698
rect 12285 20644 12309 20646
rect 12365 20644 12389 20646
rect 12445 20644 12469 20646
rect 12229 20624 12525 20644
rect 12229 19612 12525 19632
rect 12285 19610 12309 19612
rect 12365 19610 12389 19612
rect 12445 19610 12469 19612
rect 12307 19558 12309 19610
rect 12371 19558 12383 19610
rect 12445 19558 12447 19610
rect 12285 19556 12309 19558
rect 12365 19556 12389 19558
rect 12445 19556 12469 19558
rect 12229 19536 12525 19556
rect 12229 18524 12525 18544
rect 12285 18522 12309 18524
rect 12365 18522 12389 18524
rect 12445 18522 12469 18524
rect 12307 18470 12309 18522
rect 12371 18470 12383 18522
rect 12445 18470 12447 18522
rect 12285 18468 12309 18470
rect 12365 18468 12389 18470
rect 12445 18468 12469 18470
rect 12229 18448 12525 18468
rect 12229 17436 12525 17456
rect 12285 17434 12309 17436
rect 12365 17434 12389 17436
rect 12445 17434 12469 17436
rect 12307 17382 12309 17434
rect 12371 17382 12383 17434
rect 12445 17382 12447 17434
rect 12285 17380 12309 17382
rect 12365 17380 12389 17382
rect 12445 17380 12469 17382
rect 12229 17360 12525 17380
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11164 16250 11192 16594
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 16046 11192 16186
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15638 11284 15846
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9876 15162 9904 15506
rect 11256 15162 11284 15574
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10888 14618 10916 14826
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 11440 14550 11468 15302
rect 11992 15162 12020 16390
rect 12229 16348 12525 16368
rect 12285 16346 12309 16348
rect 12365 16346 12389 16348
rect 12445 16346 12469 16348
rect 12307 16294 12309 16346
rect 12371 16294 12383 16346
rect 12445 16294 12447 16346
rect 12285 16292 12309 16294
rect 12365 16292 12389 16294
rect 12445 16292 12469 16294
rect 12229 16272 12525 16292
rect 12912 15570 12940 24262
rect 13924 24262 14334 24290
rect 13924 24154 13952 24262
rect 14278 24210 14334 24262
rect 15212 24262 15806 24290
rect 13832 24126 13952 24154
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13188 19990 13216 20266
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 19514 13400 19790
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12084 14550 12112 15370
rect 12229 15260 12525 15280
rect 12285 15258 12309 15260
rect 12365 15258 12389 15260
rect 12445 15258 12469 15260
rect 12307 15206 12309 15258
rect 12371 15206 12383 15258
rect 12445 15206 12447 15258
rect 12285 15204 12309 15206
rect 12365 15204 12389 15206
rect 12445 15204 12469 15206
rect 12229 15184 12525 15204
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13004 14550 13032 14826
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 14074 10180 14214
rect 11440 14074 11468 14486
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 7748 13796 7800 13802
rect 9324 13786 9444 13814
rect 9692 13802 9720 13942
rect 12084 13814 12112 14486
rect 12229 14172 12525 14192
rect 12285 14170 12309 14172
rect 12365 14170 12389 14172
rect 12445 14170 12469 14172
rect 12307 14118 12309 14170
rect 12371 14118 12383 14170
rect 12445 14118 12447 14170
rect 12285 14116 12309 14118
rect 12365 14116 12389 14118
rect 12445 14116 12469 14118
rect 12229 14096 12525 14116
rect 13004 13938 13032 14486
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 7748 13738 7800 13744
rect 7760 13326 7788 13738
rect 9416 13734 9444 13786
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 11900 13786 12112 13814
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 5460 12986 5488 13262
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 7116 12850 7144 13262
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7116 12238 7144 12650
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 4632 11898 4660 12174
rect 4713 11996 5009 12016
rect 4769 11994 4793 11996
rect 4849 11994 4873 11996
rect 4929 11994 4953 11996
rect 4791 11942 4793 11994
rect 4855 11942 4867 11994
rect 4929 11942 4931 11994
rect 4769 11940 4793 11942
rect 4849 11940 4873 11942
rect 4929 11940 4953 11942
rect 4713 11920 5009 11940
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 5092 11762 5120 12174
rect 6656 11898 6684 12174
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 5092 11286 5120 11698
rect 6656 11354 6684 11834
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 7116 11218 7144 12038
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7300 11354 7328 11562
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 10810 4476 11086
rect 4713 10908 5009 10928
rect 4769 10906 4793 10908
rect 4849 10906 4873 10908
rect 4929 10906 4953 10908
rect 4791 10854 4793 10906
rect 4855 10854 4867 10906
rect 4929 10854 4931 10906
rect 4769 10852 4793 10854
rect 4849 10852 4873 10854
rect 4929 10852 4953 10854
rect 4713 10832 5009 10852
rect 7116 10810 7144 11154
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 4896 10532 4948 10538
rect 4896 10474 4948 10480
rect 4908 10062 4936 10474
rect 5644 10470 5672 10542
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4068 9580 4120 9586
rect 4172 9568 4200 9658
rect 4632 9586 4660 9998
rect 4713 9820 5009 9840
rect 4769 9818 4793 9820
rect 4849 9818 4873 9820
rect 4929 9818 4953 9820
rect 4791 9766 4793 9818
rect 4855 9766 4867 9818
rect 4929 9766 4931 9818
rect 4769 9764 4793 9766
rect 4849 9764 4873 9766
rect 4929 9764 4953 9766
rect 4713 9744 5009 9764
rect 4120 9540 4200 9568
rect 4620 9580 4672 9586
rect 4068 9522 4120 9528
rect 4620 9522 4672 9528
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4172 8634 4200 8910
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3988 8022 4016 8502
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4632 7886 4660 8910
rect 4713 8732 5009 8752
rect 4769 8730 4793 8732
rect 4849 8730 4873 8732
rect 4929 8730 4953 8732
rect 4791 8678 4793 8730
rect 4855 8678 4867 8730
rect 4929 8678 4931 8730
rect 4769 8676 4793 8678
rect 4849 8676 4873 8678
rect 4929 8676 4953 8678
rect 4713 8656 5009 8676
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7993 5396 8230
rect 5354 7984 5410 7993
rect 5354 7919 5410 7928
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4356 7546 4384 7822
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4632 7342 4660 7822
rect 4713 7644 5009 7664
rect 4769 7642 4793 7644
rect 4849 7642 4873 7644
rect 4929 7642 4953 7644
rect 4791 7590 4793 7642
rect 4855 7590 4867 7642
rect 4929 7590 4931 7642
rect 4769 7588 4793 7590
rect 4849 7588 4873 7590
rect 4929 7588 4953 7590
rect 4713 7568 5009 7588
rect 5170 7440 5226 7449
rect 5170 7375 5172 7384
rect 5224 7375 5226 7384
rect 5172 7346 5224 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 5184 6866 5212 7346
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 4713 6556 5009 6576
rect 4769 6554 4793 6556
rect 4849 6554 4873 6556
rect 4929 6554 4953 6556
rect 4791 6502 4793 6554
rect 4855 6502 4867 6554
rect 4929 6502 4931 6554
rect 4769 6500 4793 6502
rect 4849 6500 4873 6502
rect 4929 6500 4953 6502
rect 4713 6480 5009 6500
rect 5184 6458 5212 6802
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 4713 5468 5009 5488
rect 4769 5466 4793 5468
rect 4849 5466 4873 5468
rect 4929 5466 4953 5468
rect 4791 5414 4793 5466
rect 4855 5414 4867 5466
rect 4929 5414 4931 5466
rect 4769 5412 4793 5414
rect 4849 5412 4873 5414
rect 4929 5412 4953 5414
rect 4713 5392 5009 5412
rect 4713 4380 5009 4400
rect 4769 4378 4793 4380
rect 4849 4378 4873 4380
rect 4929 4378 4953 4380
rect 4791 4326 4793 4378
rect 4855 4326 4867 4378
rect 4929 4326 4931 4378
rect 4769 4324 4793 4326
rect 4849 4324 4873 4326
rect 4929 4324 4953 4326
rect 4713 4304 5009 4324
rect 5644 4282 5672 10406
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5724 9512 5776 9518
rect 5722 9480 5724 9489
rect 5776 9480 5778 9489
rect 5722 9415 5778 9424
rect 5736 9382 5764 9415
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5828 7954 5856 9658
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8090 6960 8298
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 5828 7546 5856 7890
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 6866 5764 7142
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 3238 54 3556 82
rect 4158 82 4214 480
rect 4448 82 4476 4218
rect 4713 3292 5009 3312
rect 4769 3290 4793 3292
rect 4849 3290 4873 3292
rect 4929 3290 4953 3292
rect 4791 3238 4793 3290
rect 4855 3238 4867 3290
rect 4929 3238 4931 3290
rect 4769 3236 4793 3238
rect 4849 3236 4873 3238
rect 4929 3236 4953 3238
rect 4713 3216 5009 3236
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4713 2204 5009 2224
rect 4769 2202 4793 2204
rect 4849 2202 4873 2204
rect 4929 2202 4953 2204
rect 4791 2150 4793 2202
rect 4855 2150 4867 2202
rect 4929 2150 4931 2202
rect 4769 2148 4793 2150
rect 4849 2148 4873 2150
rect 4929 2148 4953 2150
rect 4713 2128 5009 2148
rect 4158 54 4476 82
rect 5170 82 5226 480
rect 5460 82 5488 2314
rect 5170 54 5488 82
rect 6090 82 6146 480
rect 6196 82 6224 6598
rect 6288 6458 6316 6802
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6472 5273 6500 6598
rect 6458 5264 6514 5273
rect 6458 5199 6514 5208
rect 6090 54 6224 82
rect 6748 82 6776 7686
rect 6932 7410 6960 7890
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7010 82 7066 480
rect 7300 134 7328 10950
rect 7576 8906 7604 12786
rect 7760 12714 7788 13262
rect 8404 13258 8432 13670
rect 8471 13628 8767 13648
rect 8527 13626 8551 13628
rect 8607 13626 8631 13628
rect 8687 13626 8711 13628
rect 8549 13574 8551 13626
rect 8613 13574 8625 13626
rect 8687 13574 8689 13626
rect 8527 13572 8551 13574
rect 8607 13572 8631 13574
rect 8687 13572 8711 13574
rect 8471 13552 8767 13572
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 11830 7880 12582
rect 8220 12306 8248 12650
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11898 8248 12242
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8312 10470 8340 11154
rect 8404 10538 8432 13194
rect 9416 12782 9444 13670
rect 11900 13326 11928 13786
rect 13280 13734 13308 14350
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13832 13530 13860 24126
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14476 14958 14504 15506
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 14074 14044 14758
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13924 13530 13952 13738
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 9784 12986 9812 13262
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 11716 12850 11744 13262
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 8471 12540 8767 12560
rect 8527 12538 8551 12540
rect 8607 12538 8631 12540
rect 8687 12538 8711 12540
rect 8549 12486 8551 12538
rect 8613 12486 8625 12538
rect 8687 12486 8689 12538
rect 8527 12484 8551 12486
rect 8607 12484 8631 12486
rect 8687 12484 8711 12486
rect 8471 12464 8767 12484
rect 9324 12374 9352 12582
rect 11900 12374 11928 13262
rect 12229 13084 12525 13104
rect 12285 13082 12309 13084
rect 12365 13082 12389 13084
rect 12445 13082 12469 13084
rect 12307 13030 12309 13082
rect 12371 13030 12383 13082
rect 12445 13030 12447 13082
rect 12285 13028 12309 13030
rect 12365 13028 12389 13030
rect 12445 13028 12469 13030
rect 12229 13008 12525 13028
rect 13004 12646 13032 13330
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 9784 11898 9812 12310
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 8471 11452 8767 11472
rect 8527 11450 8551 11452
rect 8607 11450 8631 11452
rect 8687 11450 8711 11452
rect 8549 11398 8551 11450
rect 8613 11398 8625 11450
rect 8687 11398 8689 11450
rect 8527 11396 8551 11398
rect 8607 11396 8631 11398
rect 8687 11396 8711 11398
rect 8471 11376 8767 11396
rect 9954 10568 10010 10577
rect 8392 10532 8444 10538
rect 9954 10503 10010 10512
rect 8392 10474 8444 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8498 7604 8842
rect 7852 8634 7880 8910
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 6866 7972 8366
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7944 6458 7972 6802
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8312 4185 8340 10406
rect 8471 10364 8767 10384
rect 8527 10362 8551 10364
rect 8607 10362 8631 10364
rect 8687 10362 8711 10364
rect 8549 10310 8551 10362
rect 8613 10310 8625 10362
rect 8687 10310 8689 10362
rect 8527 10308 8551 10310
rect 8607 10308 8631 10310
rect 8687 10308 8711 10310
rect 8471 10288 8767 10308
rect 8471 9276 8767 9296
rect 8527 9274 8551 9276
rect 8607 9274 8631 9276
rect 8687 9274 8711 9276
rect 8549 9222 8551 9274
rect 8613 9222 8625 9274
rect 8687 9222 8689 9274
rect 8527 9220 8551 9222
rect 8607 9220 8631 9222
rect 8687 9220 8711 9222
rect 8471 9200 8767 9220
rect 8471 8188 8767 8208
rect 8527 8186 8551 8188
rect 8607 8186 8631 8188
rect 8687 8186 8711 8188
rect 8549 8134 8551 8186
rect 8613 8134 8625 8186
rect 8687 8134 8689 8186
rect 8527 8132 8551 8134
rect 8607 8132 8631 8134
rect 8687 8132 8711 8134
rect 8471 8112 8767 8132
rect 8471 7100 8767 7120
rect 8527 7098 8551 7100
rect 8607 7098 8631 7100
rect 8687 7098 8711 7100
rect 8549 7046 8551 7098
rect 8613 7046 8625 7098
rect 8687 7046 8689 7098
rect 8527 7044 8551 7046
rect 8607 7044 8631 7046
rect 8687 7044 8711 7046
rect 8471 7024 8767 7044
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8471 6012 8767 6032
rect 8527 6010 8551 6012
rect 8607 6010 8631 6012
rect 8687 6010 8711 6012
rect 8549 5958 8551 6010
rect 8613 5958 8625 6010
rect 8687 5958 8689 6010
rect 8527 5956 8551 5958
rect 8607 5956 8631 5958
rect 8687 5956 8711 5958
rect 8471 5936 8767 5956
rect 8471 4924 8767 4944
rect 8527 4922 8551 4924
rect 8607 4922 8631 4924
rect 8687 4922 8711 4924
rect 8549 4870 8551 4922
rect 8613 4870 8625 4922
rect 8687 4870 8689 4922
rect 8527 4868 8551 4870
rect 8607 4868 8631 4870
rect 8687 4868 8711 4870
rect 8471 4848 8767 4868
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8390 4040 8446 4049
rect 8390 3975 8446 3984
rect 8404 3738 8432 3975
rect 8471 3836 8767 3856
rect 8527 3834 8551 3836
rect 8607 3834 8631 3836
rect 8687 3834 8711 3836
rect 8549 3782 8551 3834
rect 8613 3782 8625 3834
rect 8687 3782 8689 3834
rect 8527 3780 8551 3782
rect 8607 3780 8631 3782
rect 8687 3780 8711 3782
rect 8471 3760 8767 3780
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 2990 8432 3538
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8471 2748 8767 2768
rect 8527 2746 8551 2748
rect 8607 2746 8631 2748
rect 8687 2746 8711 2748
rect 8549 2694 8551 2746
rect 8613 2694 8625 2746
rect 8687 2694 8689 2746
rect 8527 2692 8551 2694
rect 8607 2692 8631 2694
rect 8687 2692 8711 2694
rect 8471 2672 8767 2692
rect 6748 54 7066 82
rect 7288 128 7340 134
rect 7288 70 7340 76
rect 7930 128 7986 480
rect 7930 76 7932 128
rect 7984 76 7986 128
rect 3238 0 3294 54
rect 4158 0 4214 54
rect 5170 0 5226 54
rect 6090 0 6146 54
rect 7010 0 7066 54
rect 7930 0 7986 76
rect 8850 82 8906 480
rect 8956 82 8984 6598
rect 9968 5778 9996 10503
rect 10060 9654 10088 12174
rect 12229 11996 12525 12016
rect 12285 11994 12309 11996
rect 12365 11994 12389 11996
rect 12445 11994 12469 11996
rect 12307 11942 12309 11994
rect 12371 11942 12383 11994
rect 12445 11942 12447 11994
rect 12285 11940 12309 11942
rect 12365 11940 12389 11942
rect 12445 11940 12469 11942
rect 12229 11920 12525 11940
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 10600 10464 10652 10470
rect 11716 10452 11744 11222
rect 11808 11150 11836 11494
rect 12544 11286 12572 11562
rect 12912 11354 12940 12310
rect 13004 11898 13032 12582
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10674 11836 11086
rect 12229 10908 12525 10928
rect 12285 10906 12309 10908
rect 12365 10906 12389 10908
rect 12445 10906 12469 10908
rect 12307 10854 12309 10906
rect 12371 10854 12383 10906
rect 12445 10854 12447 10906
rect 12285 10852 12309 10854
rect 12365 10852 12389 10854
rect 12445 10852 12469 10854
rect 12229 10832 12525 10852
rect 12728 10810 12756 11222
rect 13556 11150 13584 11562
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 13556 10742 13584 11086
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 11796 10464 11848 10470
rect 11716 10424 11796 10452
rect 10600 10406 10652 10412
rect 11796 10406 11848 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3670 9168 3878
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9140 3194 9168 3606
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9232 2650 9260 4082
rect 10060 4010 10088 9590
rect 10152 9586 10180 10066
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 11716 9364 11744 10066
rect 11808 9722 11836 10406
rect 12820 10062 12848 10474
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12229 9820 12525 9840
rect 12285 9818 12309 9820
rect 12365 9818 12389 9820
rect 12445 9818 12469 9820
rect 12307 9766 12309 9818
rect 12371 9766 12383 9818
rect 12445 9766 12447 9818
rect 12285 9764 12309 9766
rect 12365 9764 12389 9766
rect 12445 9764 12469 9766
rect 12229 9744 12525 9764
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 11796 9376 11848 9382
rect 11716 9336 11796 9364
rect 11796 9318 11848 9324
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8294 11008 8978
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 7546 10364 7890
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10796 7410 10824 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10980 7313 11008 8230
rect 11072 7410 11100 8230
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11532 7546 11560 7822
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10966 7304 11022 7313
rect 10966 7239 11022 7248
rect 11072 6934 11100 7346
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 6458 10456 6734
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11072 5370 11100 5714
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 2854 9536 3878
rect 10060 3534 10088 3946
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3194 11376 3470
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 8850 54 8984 82
rect 9508 82 9536 2790
rect 9862 82 9918 480
rect 9508 54 9918 82
rect 10520 82 10548 2790
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11348 1465 11376 2450
rect 11334 1456 11390 1465
rect 11334 1391 11390 1400
rect 10782 82 10838 480
rect 10520 54 10838 82
rect 11440 82 11468 6054
rect 11808 4282 11836 9318
rect 11992 8906 12020 9318
rect 12544 9178 12572 9386
rect 12636 9178 12664 9998
rect 12820 9586 12848 9998
rect 13648 9586 13676 12174
rect 14200 11762 14228 12786
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14278 10568 14334 10577
rect 14278 10503 14334 10512
rect 14292 10266 14320 10503
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14660 9586 14688 10066
rect 15212 9722 15240 24262
rect 15750 24210 15806 24262
rect 17052 24262 17278 24290
rect 15986 22332 16282 22352
rect 16042 22330 16066 22332
rect 16122 22330 16146 22332
rect 16202 22330 16226 22332
rect 16064 22278 16066 22330
rect 16128 22278 16140 22330
rect 16202 22278 16204 22330
rect 16042 22276 16066 22278
rect 16122 22276 16146 22278
rect 16202 22276 16226 22278
rect 15986 22256 16282 22276
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 21010 15884 22034
rect 15986 21244 16282 21264
rect 16042 21242 16066 21244
rect 16122 21242 16146 21244
rect 16202 21242 16226 21244
rect 16064 21190 16066 21242
rect 16128 21190 16140 21242
rect 16202 21190 16204 21242
rect 16042 21188 16066 21190
rect 16122 21188 16146 21190
rect 16202 21188 16226 21190
rect 15986 21168 16282 21188
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15856 20602 15884 20946
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15986 20156 16282 20176
rect 16042 20154 16066 20156
rect 16122 20154 16146 20156
rect 16202 20154 16226 20156
rect 16064 20102 16066 20154
rect 16128 20102 16140 20154
rect 16202 20102 16204 20154
rect 16042 20100 16066 20102
rect 16122 20100 16146 20102
rect 16202 20100 16226 20102
rect 15986 20080 16282 20100
rect 15986 19068 16282 19088
rect 16042 19066 16066 19068
rect 16122 19066 16146 19068
rect 16202 19066 16226 19068
rect 16064 19014 16066 19066
rect 16128 19014 16140 19066
rect 16202 19014 16204 19066
rect 16042 19012 16066 19014
rect 16122 19012 16146 19014
rect 16202 19012 16226 19014
rect 15986 18992 16282 19012
rect 15986 17980 16282 18000
rect 16042 17978 16066 17980
rect 16122 17978 16146 17980
rect 16202 17978 16226 17980
rect 16064 17926 16066 17978
rect 16128 17926 16140 17978
rect 16202 17926 16204 17978
rect 16042 17924 16066 17926
rect 16122 17924 16146 17926
rect 16202 17924 16226 17926
rect 15986 17904 16282 17924
rect 15986 16892 16282 16912
rect 16042 16890 16066 16892
rect 16122 16890 16146 16892
rect 16202 16890 16226 16892
rect 16064 16838 16066 16890
rect 16128 16838 16140 16890
rect 16202 16838 16204 16890
rect 16042 16836 16066 16838
rect 16122 16836 16146 16838
rect 16202 16836 16226 16838
rect 15986 16816 16282 16836
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 15488 15706 15516 16487
rect 15986 15804 16282 15824
rect 16042 15802 16066 15804
rect 16122 15802 16146 15804
rect 16202 15802 16226 15804
rect 16064 15750 16066 15802
rect 16128 15750 16140 15802
rect 16202 15750 16204 15802
rect 16042 15748 16066 15750
rect 16122 15748 16146 15750
rect 16202 15748 16226 15750
rect 15986 15728 16282 15748
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15304 15094 15332 15506
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 12850 15424 14758
rect 15488 14550 15516 15302
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 15986 14716 16282 14736
rect 16042 14714 16066 14716
rect 16122 14714 16146 14716
rect 16202 14714 16226 14716
rect 16064 14662 16066 14714
rect 16128 14662 16140 14714
rect 16202 14662 16204 14714
rect 16042 14660 16066 14662
rect 16122 14660 16146 14662
rect 16202 14660 16226 14662
rect 15986 14640 16282 14660
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15488 14074 15516 14486
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16224 13802 16252 13874
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 15986 13628 16282 13648
rect 16042 13626 16066 13628
rect 16122 13626 16146 13628
rect 16202 13626 16226 13628
rect 16064 13574 16066 13626
rect 16128 13574 16140 13626
rect 16202 13574 16204 13626
rect 16042 13572 16066 13574
rect 16122 13572 16146 13574
rect 16202 13572 16226 13574
rect 15986 13552 16282 13572
rect 16500 13530 16528 13738
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16868 13394 16896 14894
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15488 12646 15516 13330
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15986 12540 16282 12560
rect 16042 12538 16066 12540
rect 16122 12538 16146 12540
rect 16202 12538 16226 12540
rect 16064 12486 16066 12538
rect 16128 12486 16140 12538
rect 16202 12486 16204 12538
rect 16042 12484 16066 12486
rect 16122 12484 16146 12486
rect 16202 12484 16226 12486
rect 15986 12464 16282 12484
rect 15986 11452 16282 11472
rect 16042 11450 16066 11452
rect 16122 11450 16146 11452
rect 16202 11450 16226 11452
rect 16064 11398 16066 11450
rect 16128 11398 16140 11450
rect 16202 11398 16204 11450
rect 16042 11396 16066 11398
rect 16122 11396 16146 11398
rect 16202 11396 16226 11398
rect 15986 11376 16282 11396
rect 15986 10364 16282 10384
rect 16042 10362 16066 10364
rect 16122 10362 16146 10364
rect 16202 10362 16226 10364
rect 16064 10310 16066 10362
rect 16128 10310 16140 10362
rect 16202 10310 16204 10362
rect 16042 10308 16066 10310
rect 16122 10308 16146 10310
rect 16202 10308 16226 10310
rect 15986 10288 16282 10308
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14004 9512 14056 9518
rect 13358 9480 13414 9489
rect 14004 9454 14056 9460
rect 13358 9415 13414 9424
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6118 11928 6666
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5914 11928 6054
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3534 11652 3878
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11624 3058 11652 3470
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11808 2514 11836 4218
rect 11992 3641 12020 8842
rect 12084 8294 12112 8910
rect 12229 8732 12525 8752
rect 12285 8730 12309 8732
rect 12365 8730 12389 8732
rect 12445 8730 12469 8732
rect 12307 8678 12309 8730
rect 12371 8678 12383 8730
rect 12445 8678 12447 8730
rect 12285 8676 12309 8678
rect 12365 8676 12389 8678
rect 12445 8676 12469 8678
rect 12229 8656 12525 8676
rect 12912 8498 12940 8910
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12084 6798 12112 7822
rect 12229 7644 12525 7664
rect 12285 7642 12309 7644
rect 12365 7642 12389 7644
rect 12445 7642 12469 7644
rect 12307 7590 12309 7642
rect 12371 7590 12383 7642
rect 12445 7590 12447 7642
rect 12285 7588 12309 7590
rect 12365 7588 12389 7590
rect 12445 7588 12469 7590
rect 12229 7568 12525 7588
rect 13372 7478 13400 9415
rect 14016 9178 14044 9454
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14476 8498 14504 9522
rect 14660 9489 14688 9522
rect 14646 9480 14702 9489
rect 14646 9415 14702 9424
rect 15986 9276 16282 9296
rect 16042 9274 16066 9276
rect 16122 9274 16146 9276
rect 16202 9274 16226 9276
rect 16064 9222 16066 9274
rect 16128 9222 16140 9274
rect 16202 9222 16204 9274
rect 16042 9220 16066 9222
rect 16122 9220 16146 9222
rect 16202 9220 16226 9222
rect 15986 9200 16282 9220
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13740 7546 13768 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13740 6934 13768 7482
rect 13924 7410 13952 7822
rect 14292 7818 14320 8230
rect 15986 8188 16282 8208
rect 16042 8186 16066 8188
rect 16122 8186 16146 8188
rect 16202 8186 16226 8188
rect 16064 8134 16066 8186
rect 16128 8134 16140 8186
rect 16202 8134 16204 8186
rect 16042 8132 16066 8134
rect 16122 8132 16146 8134
rect 16202 8132 16226 8134
rect 15986 8112 16282 8132
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7410 14320 7754
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 7002 15240 7142
rect 15986 7100 16282 7120
rect 16042 7098 16066 7100
rect 16122 7098 16146 7100
rect 16202 7098 16226 7100
rect 16064 7046 16066 7098
rect 16128 7046 16140 7098
rect 16202 7046 16204 7098
rect 16042 7044 16066 7046
rect 16122 7044 16146 7046
rect 16202 7044 16226 7046
rect 15986 7024 16282 7044
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6458 12112 6734
rect 12229 6556 12525 6576
rect 12285 6554 12309 6556
rect 12365 6554 12389 6556
rect 12445 6554 12469 6556
rect 12307 6502 12309 6554
rect 12371 6502 12383 6554
rect 12445 6502 12447 6554
rect 12285 6500 12309 6502
rect 12365 6500 12389 6502
rect 12445 6500 12469 6502
rect 12229 6480 12525 6500
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 13464 6118 13492 6802
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6322 15332 6734
rect 16946 6352 17002 6361
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15384 6316 15436 6322
rect 16946 6287 17002 6296
rect 15384 6258 15436 6264
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 12229 5468 12525 5488
rect 12285 5466 12309 5468
rect 12365 5466 12389 5468
rect 12445 5466 12469 5468
rect 12307 5414 12309 5466
rect 12371 5414 12383 5466
rect 12445 5414 12447 5466
rect 12285 5412 12309 5414
rect 12365 5412 12389 5414
rect 12445 5412 12469 5414
rect 12229 5392 12525 5412
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4758 12848 4966
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12229 4380 12525 4400
rect 12285 4378 12309 4380
rect 12365 4378 12389 4380
rect 12445 4378 12469 4380
rect 12307 4326 12309 4378
rect 12371 4326 12383 4378
rect 12445 4326 12447 4378
rect 12285 4324 12309 4326
rect 12365 4324 12389 4326
rect 12445 4324 12469 4326
rect 12229 4304 12525 4324
rect 12820 4282 12848 4694
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12912 4154 12940 6054
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 12820 4126 12940 4154
rect 11978 3632 12034 3641
rect 11978 3567 12034 3576
rect 12229 3292 12525 3312
rect 12285 3290 12309 3292
rect 12365 3290 12389 3292
rect 12445 3290 12469 3292
rect 12307 3238 12309 3290
rect 12371 3238 12383 3290
rect 12445 3238 12447 3290
rect 12285 3236 12309 3238
rect 12365 3236 12389 3238
rect 12445 3236 12469 3238
rect 12229 3216 12525 3236
rect 12820 2582 12848 4126
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12229 2204 12525 2224
rect 12285 2202 12309 2204
rect 12365 2202 12389 2204
rect 12445 2202 12469 2204
rect 12307 2150 12309 2202
rect 12371 2150 12383 2202
rect 12445 2150 12447 2202
rect 12285 2148 12309 2150
rect 12365 2148 12389 2150
rect 12445 2148 12469 2150
rect 12229 2128 12525 2148
rect 12636 626 12664 2314
rect 12544 598 12664 626
rect 11702 82 11758 480
rect 11440 54 11758 82
rect 12544 82 12572 598
rect 12622 82 12678 480
rect 12544 54 12678 82
rect 13280 82 13308 5510
rect 13372 5030 13400 5714
rect 14200 5642 14228 6122
rect 15396 5710 15424 6258
rect 16960 6254 16988 6287
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14200 5370 14228 5578
rect 15396 5370 15424 5646
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 14200 5166 14228 5306
rect 15488 5234 15516 6054
rect 15986 6012 16282 6032
rect 16042 6010 16066 6012
rect 16122 6010 16146 6012
rect 16202 6010 16226 6012
rect 16064 5958 16066 6010
rect 16128 5958 16140 6010
rect 16202 5958 16204 6010
rect 16042 5956 16066 5958
rect 16122 5956 16146 5958
rect 16202 5956 16226 5958
rect 15986 5936 16282 5956
rect 17052 5914 17080 24262
rect 17222 24210 17278 24262
rect 18524 24262 18842 24290
rect 17590 23624 17646 23633
rect 17590 23559 17646 23568
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17512 20602 17540 20742
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17604 20466 17632 23559
rect 18524 21690 18552 24262
rect 18786 24210 18842 24262
rect 20258 24290 20314 24690
rect 21730 24290 21786 24690
rect 20258 24262 20392 24290
rect 20258 24210 20314 24262
rect 19154 22536 19210 22545
rect 19154 22471 19210 22480
rect 19168 22098 19196 22471
rect 19522 22128 19578 22137
rect 19156 22092 19208 22098
rect 19522 22063 19578 22072
rect 19156 22034 19208 22040
rect 19168 21690 19196 22034
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19352 21554 19380 21830
rect 19536 21690 19564 22063
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19524 21684 19576 21690
rect 19524 21626 19576 21632
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21078 18644 21286
rect 19352 21146 19380 21490
rect 19536 21486 19564 21626
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 20602 17816 20878
rect 18616 20602 18644 21014
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 18892 19990 18920 20878
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18970 19816 19026 19825
rect 18248 19514 18276 19790
rect 18970 19751 19026 19760
rect 18984 19514 19012 19751
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18984 19310 19012 19450
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19352 18902 19380 19654
rect 19444 19378 19472 21286
rect 19628 20806 19656 21966
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 19744 21788 20040 21808
rect 19800 21786 19824 21788
rect 19880 21786 19904 21788
rect 19960 21786 19984 21788
rect 19822 21734 19824 21786
rect 19886 21734 19898 21786
rect 19960 21734 19962 21786
rect 19800 21732 19824 21734
rect 19880 21732 19904 21734
rect 19960 21732 19984 21734
rect 19744 21712 20040 21732
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19744 20700 20040 20720
rect 19800 20698 19824 20700
rect 19880 20698 19904 20700
rect 19960 20698 19984 20700
rect 19822 20646 19824 20698
rect 19886 20646 19898 20698
rect 19960 20646 19962 20698
rect 19800 20644 19824 20646
rect 19880 20644 19904 20646
rect 19960 20644 19984 20646
rect 19744 20624 20040 20644
rect 19522 20496 19578 20505
rect 19522 20431 19578 20440
rect 19536 19922 19564 20431
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19628 20058 19656 20266
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19536 19514 19564 19858
rect 19744 19612 20040 19632
rect 19800 19610 19824 19612
rect 19880 19610 19904 19612
rect 19960 19610 19984 19612
rect 19822 19558 19824 19610
rect 19886 19558 19898 19610
rect 19960 19558 19962 19610
rect 19800 19556 19824 19558
rect 19880 19556 19904 19558
rect 19960 19556 19984 19558
rect 19744 19536 20040 19556
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19614 19272 19670 19281
rect 19432 19236 19484 19242
rect 20088 19242 20116 21490
rect 20180 19281 20208 21898
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20272 20330 20300 20810
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20166 19272 20222 19281
rect 19614 19207 19670 19216
rect 20076 19236 20128 19242
rect 19432 19178 19484 19184
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19352 18426 19380 18838
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19444 18306 19472 19178
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19352 18278 19472 18306
rect 17498 15464 17554 15473
rect 17498 15399 17554 15408
rect 17512 15162 17540 15399
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17512 14958 17540 15098
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14550 17264 14758
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17144 13802 17172 14282
rect 17236 14074 17264 14486
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17972 13938 18000 14350
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5370 16896 5714
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16302 5264 16358 5273
rect 15476 5228 15528 5234
rect 16302 5199 16358 5208
rect 15476 5170 15528 5176
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 13372 4622 13400 4966
rect 14752 4690 14780 4966
rect 15986 4924 16282 4944
rect 16042 4922 16066 4924
rect 16122 4922 16146 4924
rect 16202 4922 16226 4924
rect 16064 4870 16066 4922
rect 16128 4870 16140 4922
rect 16202 4870 16204 4922
rect 16042 4868 16066 4870
rect 16122 4868 16146 4870
rect 16202 4868 16226 4870
rect 15986 4848 16282 4868
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13372 4146 13400 4558
rect 15304 4282 15332 4626
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 13542 82 13598 480
rect 13280 54 13598 82
rect 8850 0 8906 54
rect 9862 0 9918 54
rect 10782 0 10838 54
rect 11702 0 11758 54
rect 12622 0 12678 54
rect 13542 0 13598 54
rect 14554 82 14610 480
rect 14660 82 14688 2314
rect 14554 54 14688 82
rect 15474 82 15530 480
rect 15580 82 15608 4422
rect 15986 3836 16282 3856
rect 16042 3834 16066 3836
rect 16122 3834 16146 3836
rect 16202 3834 16226 3836
rect 16064 3782 16066 3834
rect 16128 3782 16140 3834
rect 16202 3782 16204 3834
rect 16042 3780 16066 3782
rect 16122 3780 16146 3782
rect 16202 3780 16226 3782
rect 15986 3760 16282 3780
rect 15986 2748 16282 2768
rect 16042 2746 16066 2748
rect 16122 2746 16146 2748
rect 16202 2746 16226 2748
rect 16064 2694 16066 2746
rect 16128 2694 16140 2746
rect 16202 2694 16204 2746
rect 16042 2692 16066 2694
rect 16122 2692 16146 2694
rect 16202 2692 16226 2694
rect 15986 2672 16282 2692
rect 15474 54 15608 82
rect 16316 82 16344 5199
rect 17144 3670 17172 13738
rect 17972 13462 18000 13874
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17972 12986 18000 13398
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18616 12850 18644 13262
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17788 10810 17816 11086
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17420 10198 17448 10542
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17420 8906 17448 10134
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17880 9722 17908 9998
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17420 6458 17448 6802
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17328 4214 17356 4490
rect 17972 4282 18000 4558
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17316 4208 17368 4214
rect 17316 4150 17368 4156
rect 18064 4154 18092 12582
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18340 11830 18368 12174
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18432 11286 18460 12650
rect 18616 12238 18644 12786
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11694 18644 12174
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10674 18184 10950
rect 18432 10674 18460 11222
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18432 9994 18460 10610
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 9042 18644 9318
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 7993 18644 8978
rect 19260 8498 19288 11698
rect 19352 11626 19380 18278
rect 19430 17640 19486 17649
rect 19430 17575 19486 17584
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10742 19380 11086
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19444 9722 19472 17575
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 8634 19472 9318
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 18602 7984 18658 7993
rect 18602 7919 18658 7928
rect 19076 7410 19104 8366
rect 19260 7954 19288 8434
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7546 19288 7890
rect 19248 7540 19300 7546
rect 19536 7528 19564 18906
rect 19628 18766 19656 19207
rect 20166 19207 20222 19216
rect 20076 19178 20128 19184
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19744 18524 20040 18544
rect 19800 18522 19824 18524
rect 19880 18522 19904 18524
rect 19960 18522 19984 18524
rect 19822 18470 19824 18522
rect 19886 18470 19898 18522
rect 19960 18470 19962 18522
rect 19800 18468 19824 18470
rect 19880 18468 19904 18470
rect 19960 18468 19984 18470
rect 19744 18448 20040 18468
rect 19744 17436 20040 17456
rect 19800 17434 19824 17436
rect 19880 17434 19904 17436
rect 19960 17434 19984 17436
rect 19822 17382 19824 17434
rect 19886 17382 19898 17434
rect 19960 17382 19962 17434
rect 19800 17380 19824 17382
rect 19880 17380 19904 17382
rect 19960 17380 19984 17382
rect 19744 17360 20040 17380
rect 19744 16348 20040 16368
rect 19800 16346 19824 16348
rect 19880 16346 19904 16348
rect 19960 16346 19984 16348
rect 19822 16294 19824 16346
rect 19886 16294 19898 16346
rect 19960 16294 19962 16346
rect 19800 16292 19824 16294
rect 19880 16292 19904 16294
rect 19960 16292 19984 16294
rect 19744 16272 20040 16292
rect 19744 15260 20040 15280
rect 19800 15258 19824 15260
rect 19880 15258 19904 15260
rect 19960 15258 19984 15260
rect 19822 15206 19824 15258
rect 19886 15206 19898 15258
rect 19960 15206 19962 15258
rect 19800 15204 19824 15206
rect 19880 15204 19904 15206
rect 19960 15204 19984 15206
rect 19744 15184 20040 15204
rect 19744 14172 20040 14192
rect 19800 14170 19824 14172
rect 19880 14170 19904 14172
rect 19960 14170 19984 14172
rect 19822 14118 19824 14170
rect 19886 14118 19898 14170
rect 19960 14118 19962 14170
rect 19800 14116 19824 14118
rect 19880 14116 19904 14118
rect 19960 14116 19984 14118
rect 19744 14096 20040 14116
rect 19744 13084 20040 13104
rect 19800 13082 19824 13084
rect 19880 13082 19904 13084
rect 19960 13082 19984 13084
rect 19822 13030 19824 13082
rect 19886 13030 19898 13082
rect 19960 13030 19962 13082
rect 19800 13028 19824 13030
rect 19880 13028 19904 13030
rect 19960 13028 19984 13030
rect 19744 13008 20040 13028
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 11898 19656 12718
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19744 11996 20040 12016
rect 19800 11994 19824 11996
rect 19880 11994 19904 11996
rect 19960 11994 19984 11996
rect 19822 11942 19824 11994
rect 19886 11942 19898 11994
rect 19960 11942 19962 11994
rect 19800 11940 19824 11942
rect 19880 11940 19904 11942
rect 19960 11940 19984 11942
rect 19744 11920 20040 11940
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19628 10742 19656 11562
rect 19744 10908 20040 10928
rect 19800 10906 19824 10908
rect 19880 10906 19904 10908
rect 19960 10906 19984 10908
rect 19822 10854 19824 10906
rect 19886 10854 19898 10906
rect 19960 10854 19962 10906
rect 19800 10852 19824 10854
rect 19880 10852 19904 10854
rect 19960 10852 19984 10854
rect 19744 10832 20040 10852
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 20088 10674 20116 12038
rect 20272 11830 20300 20266
rect 20364 18970 20392 24262
rect 21376 24262 21786 24290
rect 21376 20534 21404 24262
rect 21730 24210 21786 24262
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 22098 19000 22154 19009
rect 20352 18964 20404 18970
rect 22098 18935 22154 18944
rect 20352 18906 20404 18912
rect 22112 17241 22140 18935
rect 22098 17232 22154 17241
rect 22098 17167 22154 17176
rect 22098 13832 22154 13841
rect 22098 13767 22154 13776
rect 21086 13152 21142 13161
rect 21086 13087 21142 13096
rect 21100 12986 21128 13087
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 22112 12918 22140 13767
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20272 11286 20300 11766
rect 20732 11558 20760 12242
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20260 11280 20312 11286
rect 20166 11248 20222 11257
rect 20260 11222 20312 11228
rect 20166 11183 20222 11192
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20180 10266 20208 11183
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 19744 9820 20040 9840
rect 19800 9818 19824 9820
rect 19880 9818 19904 9820
rect 19960 9818 19984 9820
rect 19822 9766 19824 9818
rect 19886 9766 19898 9818
rect 19960 9766 19962 9818
rect 19800 9764 19824 9766
rect 19880 9764 19904 9766
rect 19960 9764 19984 9766
rect 19744 9744 20040 9764
rect 20180 9722 20208 10066
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20166 9344 20222 9353
rect 20166 9279 20222 9288
rect 20180 9178 20208 9279
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20260 9036 20312 9042
rect 20260 8978 20312 8984
rect 19744 8732 20040 8752
rect 19800 8730 19824 8732
rect 19880 8730 19904 8732
rect 19960 8730 19984 8732
rect 19822 8678 19824 8730
rect 19886 8678 19898 8730
rect 19960 8678 19962 8730
rect 19800 8676 19824 8678
rect 19880 8676 19904 8678
rect 19960 8676 19984 8678
rect 19744 8656 20040 8676
rect 20166 8664 20222 8673
rect 20166 8599 20222 8608
rect 20180 8566 20208 8599
rect 20168 8560 20220 8566
rect 20168 8502 20220 8508
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19628 8090 19656 8366
rect 20272 8294 20300 8978
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19744 7644 20040 7664
rect 19800 7642 19824 7644
rect 19880 7642 19904 7644
rect 19960 7642 19984 7644
rect 19822 7590 19824 7642
rect 19886 7590 19898 7642
rect 19960 7590 19962 7642
rect 19800 7588 19824 7590
rect 19880 7588 19904 7590
rect 19960 7588 19984 7590
rect 19744 7568 20040 7588
rect 19248 7482 19300 7488
rect 19444 7500 19564 7528
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6118 19288 6734
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 4690 19472 7500
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 6798 19564 7346
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19744 6556 20040 6576
rect 19800 6554 19824 6556
rect 19880 6554 19904 6556
rect 19960 6554 19984 6556
rect 19822 6502 19824 6554
rect 19886 6502 19898 6554
rect 19960 6502 19962 6554
rect 19800 6500 19824 6502
rect 19880 6500 19904 6502
rect 19960 6500 19984 6502
rect 19744 6480 20040 6500
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5710 19656 6054
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 20166 5536 20222 5545
rect 19744 5468 20040 5488
rect 20166 5471 20222 5480
rect 19800 5466 19824 5468
rect 19880 5466 19904 5468
rect 19960 5466 19984 5468
rect 19822 5414 19824 5466
rect 19886 5414 19898 5466
rect 19960 5414 19962 5466
rect 19800 5412 19824 5414
rect 19880 5412 19904 5414
rect 19960 5412 19984 5414
rect 19744 5392 20040 5412
rect 20180 5370 20208 5471
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20180 5166 20208 5306
rect 20168 5160 20220 5166
rect 20272 5137 20300 8230
rect 20168 5102 20220 5108
rect 20258 5128 20314 5137
rect 20258 5063 20314 5072
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 17328 3670 17356 4150
rect 17972 4126 18092 4154
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17144 3058 17172 3606
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16592 2650 16620 2858
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16394 82 16450 480
rect 16316 54 16450 82
rect 16960 82 16988 2246
rect 17314 82 17370 480
rect 16960 54 17370 82
rect 17972 82 18000 4126
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3670 18276 3878
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18248 3194 18276 3606
rect 18340 3534 18368 4218
rect 18892 4010 18920 4422
rect 19444 4282 19472 4626
rect 19744 4380 20040 4400
rect 19800 4378 19824 4380
rect 19880 4378 19904 4380
rect 19960 4378 19984 4380
rect 19822 4326 19824 4378
rect 19886 4326 19898 4378
rect 19960 4326 19962 4378
rect 19800 4324 19824 4326
rect 19880 4324 19904 4326
rect 19960 4324 19984 4326
rect 19744 4304 20040 4324
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19168 4146 19196 4218
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 20074 4040 20130 4049
rect 18880 4004 18932 4010
rect 20074 3975 20130 3984
rect 18880 3946 18932 3952
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 3058 18368 3470
rect 19744 3292 20040 3312
rect 19800 3290 19824 3292
rect 19880 3290 19904 3292
rect 19960 3290 19984 3292
rect 19822 3238 19824 3290
rect 19886 3238 19898 3290
rect 19960 3238 19962 3290
rect 19800 3236 19824 3238
rect 19880 3236 19904 3238
rect 19960 3236 19984 3238
rect 19744 3216 20040 3236
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18616 2650 18644 2858
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18234 82 18290 480
rect 17972 54 18290 82
rect 18984 82 19012 2246
rect 19744 2204 20040 2224
rect 19800 2202 19824 2204
rect 19880 2202 19904 2204
rect 19960 2202 19984 2204
rect 19822 2150 19824 2202
rect 19886 2150 19898 2202
rect 19960 2150 19962 2202
rect 19800 2148 19824 2150
rect 19880 2148 19904 2150
rect 19960 2148 19984 2150
rect 19744 2128 20040 2148
rect 19246 82 19302 480
rect 18984 54 19302 82
rect 20088 82 20116 3975
rect 20166 82 20222 480
rect 20088 54 20222 82
rect 20732 82 20760 11494
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21086 82 21142 480
rect 20732 54 21142 82
rect 21836 82 21864 10406
rect 22006 82 22062 480
rect 21836 54 22062 82
rect 14554 0 14610 54
rect 15474 0 15530 54
rect 16394 0 16450 54
rect 17314 0 17370 54
rect 18234 0 18290 54
rect 19246 0 19302 54
rect 20166 0 20222 54
rect 21086 0 21142 54
rect 22006 0 22062 54
<< via2 >>
rect 1306 23432 1362 23488
rect 110 22752 166 22808
rect 3514 20984 3570 21040
rect 1582 19760 1638 19816
rect 110 19080 166 19136
rect 2778 17312 2834 17368
rect 110 12960 166 13016
rect 1398 9832 1454 9888
rect 2502 11872 2558 11928
rect 2594 8608 2650 8664
rect 110 5480 166 5536
rect 2686 7248 2742 7304
rect 1306 2352 1362 2408
rect 2226 1400 2282 1456
rect 3882 10512 3938 10568
rect 4713 21786 4769 21788
rect 4793 21786 4849 21788
rect 4873 21786 4929 21788
rect 4953 21786 5009 21788
rect 4713 21734 4739 21786
rect 4739 21734 4769 21786
rect 4793 21734 4803 21786
rect 4803 21734 4849 21786
rect 4873 21734 4919 21786
rect 4919 21734 4929 21786
rect 4953 21734 4983 21786
rect 4983 21734 5009 21786
rect 4713 21732 4769 21734
rect 4793 21732 4849 21734
rect 4873 21732 4929 21734
rect 4953 21732 5009 21734
rect 8471 22330 8527 22332
rect 8551 22330 8607 22332
rect 8631 22330 8687 22332
rect 8711 22330 8767 22332
rect 8471 22278 8497 22330
rect 8497 22278 8527 22330
rect 8551 22278 8561 22330
rect 8561 22278 8607 22330
rect 8631 22278 8677 22330
rect 8677 22278 8687 22330
rect 8711 22278 8741 22330
rect 8741 22278 8767 22330
rect 8471 22276 8527 22278
rect 8551 22276 8607 22278
rect 8631 22276 8687 22278
rect 8711 22276 8767 22278
rect 8471 21242 8527 21244
rect 8551 21242 8607 21244
rect 8631 21242 8687 21244
rect 8711 21242 8767 21244
rect 8471 21190 8497 21242
rect 8497 21190 8527 21242
rect 8551 21190 8561 21242
rect 8561 21190 8607 21242
rect 8631 21190 8677 21242
rect 8677 21190 8687 21242
rect 8711 21190 8741 21242
rect 8741 21190 8767 21242
rect 8471 21188 8527 21190
rect 8551 21188 8607 21190
rect 8631 21188 8687 21190
rect 8711 21188 8767 21190
rect 4713 20698 4769 20700
rect 4793 20698 4849 20700
rect 4873 20698 4929 20700
rect 4953 20698 5009 20700
rect 4713 20646 4739 20698
rect 4739 20646 4769 20698
rect 4793 20646 4803 20698
rect 4803 20646 4849 20698
rect 4873 20646 4919 20698
rect 4919 20646 4929 20698
rect 4953 20646 4983 20698
rect 4983 20646 5009 20698
rect 4713 20644 4769 20646
rect 4793 20644 4849 20646
rect 4873 20644 4929 20646
rect 4953 20644 5009 20646
rect 4713 19610 4769 19612
rect 4793 19610 4849 19612
rect 4873 19610 4929 19612
rect 4953 19610 5009 19612
rect 4713 19558 4739 19610
rect 4739 19558 4769 19610
rect 4793 19558 4803 19610
rect 4803 19558 4849 19610
rect 4873 19558 4919 19610
rect 4919 19558 4929 19610
rect 4953 19558 4983 19610
rect 4983 19558 5009 19610
rect 4713 19556 4769 19558
rect 4793 19556 4849 19558
rect 4873 19556 4929 19558
rect 4953 19556 5009 19558
rect 8471 20154 8527 20156
rect 8551 20154 8607 20156
rect 8631 20154 8687 20156
rect 8711 20154 8767 20156
rect 8471 20102 8497 20154
rect 8497 20102 8527 20154
rect 8551 20102 8561 20154
rect 8561 20102 8607 20154
rect 8631 20102 8677 20154
rect 8677 20102 8687 20154
rect 8711 20102 8741 20154
rect 8741 20102 8767 20154
rect 8471 20100 8527 20102
rect 8551 20100 8607 20102
rect 8631 20100 8687 20102
rect 8711 20100 8767 20102
rect 7378 19216 7434 19272
rect 8471 19066 8527 19068
rect 8551 19066 8607 19068
rect 8631 19066 8687 19068
rect 8711 19066 8767 19068
rect 8471 19014 8497 19066
rect 8497 19014 8527 19066
rect 8551 19014 8561 19066
rect 8561 19014 8607 19066
rect 8631 19014 8677 19066
rect 8677 19014 8687 19066
rect 8711 19014 8741 19066
rect 8741 19014 8767 19066
rect 8471 19012 8527 19014
rect 8551 19012 8607 19014
rect 8631 19012 8687 19014
rect 8711 19012 8767 19014
rect 4713 18522 4769 18524
rect 4793 18522 4849 18524
rect 4873 18522 4929 18524
rect 4953 18522 5009 18524
rect 4713 18470 4739 18522
rect 4739 18470 4769 18522
rect 4793 18470 4803 18522
rect 4803 18470 4849 18522
rect 4873 18470 4919 18522
rect 4919 18470 4929 18522
rect 4953 18470 4983 18522
rect 4983 18470 5009 18522
rect 4713 18468 4769 18470
rect 4793 18468 4849 18470
rect 4873 18468 4929 18470
rect 4953 18468 5009 18470
rect 8471 17978 8527 17980
rect 8551 17978 8607 17980
rect 8631 17978 8687 17980
rect 8711 17978 8767 17980
rect 8471 17926 8497 17978
rect 8497 17926 8527 17978
rect 8551 17926 8561 17978
rect 8561 17926 8607 17978
rect 8631 17926 8677 17978
rect 8677 17926 8687 17978
rect 8711 17926 8741 17978
rect 8741 17926 8767 17978
rect 8471 17924 8527 17926
rect 8551 17924 8607 17926
rect 8631 17924 8687 17926
rect 8711 17924 8767 17926
rect 4713 17434 4769 17436
rect 4793 17434 4849 17436
rect 4873 17434 4929 17436
rect 4953 17434 5009 17436
rect 4713 17382 4739 17434
rect 4739 17382 4769 17434
rect 4793 17382 4803 17434
rect 4803 17382 4849 17434
rect 4873 17382 4919 17434
rect 4919 17382 4929 17434
rect 4953 17382 4983 17434
rect 4983 17382 5009 17434
rect 4713 17380 4769 17382
rect 4793 17380 4849 17382
rect 4873 17380 4929 17382
rect 4953 17380 5009 17382
rect 8390 17040 8446 17096
rect 8471 16890 8527 16892
rect 8551 16890 8607 16892
rect 8631 16890 8687 16892
rect 8711 16890 8767 16892
rect 8471 16838 8497 16890
rect 8497 16838 8527 16890
rect 8551 16838 8561 16890
rect 8561 16838 8607 16890
rect 8631 16838 8677 16890
rect 8677 16838 8687 16890
rect 8711 16838 8741 16890
rect 8741 16838 8767 16890
rect 8471 16836 8527 16838
rect 8551 16836 8607 16838
rect 8631 16836 8687 16838
rect 8711 16836 8767 16838
rect 4713 16346 4769 16348
rect 4793 16346 4849 16348
rect 4873 16346 4929 16348
rect 4953 16346 5009 16348
rect 4713 16294 4739 16346
rect 4739 16294 4769 16346
rect 4793 16294 4803 16346
rect 4803 16294 4849 16346
rect 4873 16294 4919 16346
rect 4919 16294 4929 16346
rect 4953 16294 4983 16346
rect 4983 16294 5009 16346
rect 4713 16292 4769 16294
rect 4793 16292 4849 16294
rect 4873 16292 4929 16294
rect 4953 16292 5009 16294
rect 4713 15258 4769 15260
rect 4793 15258 4849 15260
rect 4873 15258 4929 15260
rect 4953 15258 5009 15260
rect 4713 15206 4739 15258
rect 4739 15206 4769 15258
rect 4793 15206 4803 15258
rect 4803 15206 4849 15258
rect 4873 15206 4919 15258
rect 4919 15206 4929 15258
rect 4953 15206 4983 15258
rect 4983 15206 5009 15258
rect 4713 15204 4769 15206
rect 4793 15204 4849 15206
rect 4873 15204 4929 15206
rect 4953 15204 5009 15206
rect 4618 15000 4674 15056
rect 7378 14900 7380 14920
rect 7380 14900 7432 14920
rect 7432 14900 7434 14920
rect 7378 14864 7434 14900
rect 9310 16088 9366 16144
rect 8471 15802 8527 15804
rect 8551 15802 8607 15804
rect 8631 15802 8687 15804
rect 8711 15802 8767 15804
rect 8471 15750 8497 15802
rect 8497 15750 8527 15802
rect 8551 15750 8561 15802
rect 8561 15750 8607 15802
rect 8631 15750 8677 15802
rect 8677 15750 8687 15802
rect 8711 15750 8741 15802
rect 8741 15750 8767 15802
rect 8471 15748 8527 15750
rect 8551 15748 8607 15750
rect 8631 15748 8687 15750
rect 8711 15748 8767 15750
rect 8471 14714 8527 14716
rect 8551 14714 8607 14716
rect 8631 14714 8687 14716
rect 8711 14714 8767 14716
rect 8471 14662 8497 14714
rect 8497 14662 8527 14714
rect 8551 14662 8561 14714
rect 8561 14662 8607 14714
rect 8631 14662 8677 14714
rect 8677 14662 8687 14714
rect 8711 14662 8741 14714
rect 8741 14662 8767 14714
rect 8471 14660 8527 14662
rect 8551 14660 8607 14662
rect 8631 14660 8687 14662
rect 8711 14660 8767 14662
rect 4713 14170 4769 14172
rect 4793 14170 4849 14172
rect 4873 14170 4929 14172
rect 4953 14170 5009 14172
rect 4713 14118 4739 14170
rect 4739 14118 4769 14170
rect 4793 14118 4803 14170
rect 4803 14118 4849 14170
rect 4873 14118 4919 14170
rect 4919 14118 4929 14170
rect 4953 14118 4983 14170
rect 4983 14118 5009 14170
rect 4713 14116 4769 14118
rect 4793 14116 4849 14118
rect 4873 14116 4929 14118
rect 4953 14116 5009 14118
rect 4250 13640 4306 13696
rect 4713 13082 4769 13084
rect 4793 13082 4849 13084
rect 4873 13082 4929 13084
rect 4953 13082 5009 13084
rect 4713 13030 4739 13082
rect 4739 13030 4769 13082
rect 4793 13030 4803 13082
rect 4803 13030 4849 13082
rect 4873 13030 4919 13082
rect 4919 13030 4929 13082
rect 4953 13030 4983 13082
rect 4983 13030 5009 13082
rect 4713 13028 4769 13030
rect 4793 13028 4849 13030
rect 4873 13028 4929 13030
rect 4953 13028 5009 13030
rect 12229 21786 12285 21788
rect 12309 21786 12365 21788
rect 12389 21786 12445 21788
rect 12469 21786 12525 21788
rect 12229 21734 12255 21786
rect 12255 21734 12285 21786
rect 12309 21734 12319 21786
rect 12319 21734 12365 21786
rect 12389 21734 12435 21786
rect 12435 21734 12445 21786
rect 12469 21734 12499 21786
rect 12499 21734 12525 21786
rect 12229 21732 12285 21734
rect 12309 21732 12365 21734
rect 12389 21732 12445 21734
rect 12469 21732 12525 21734
rect 12229 20698 12285 20700
rect 12309 20698 12365 20700
rect 12389 20698 12445 20700
rect 12469 20698 12525 20700
rect 12229 20646 12255 20698
rect 12255 20646 12285 20698
rect 12309 20646 12319 20698
rect 12319 20646 12365 20698
rect 12389 20646 12435 20698
rect 12435 20646 12445 20698
rect 12469 20646 12499 20698
rect 12499 20646 12525 20698
rect 12229 20644 12285 20646
rect 12309 20644 12365 20646
rect 12389 20644 12445 20646
rect 12469 20644 12525 20646
rect 12229 19610 12285 19612
rect 12309 19610 12365 19612
rect 12389 19610 12445 19612
rect 12469 19610 12525 19612
rect 12229 19558 12255 19610
rect 12255 19558 12285 19610
rect 12309 19558 12319 19610
rect 12319 19558 12365 19610
rect 12389 19558 12435 19610
rect 12435 19558 12445 19610
rect 12469 19558 12499 19610
rect 12499 19558 12525 19610
rect 12229 19556 12285 19558
rect 12309 19556 12365 19558
rect 12389 19556 12445 19558
rect 12469 19556 12525 19558
rect 12229 18522 12285 18524
rect 12309 18522 12365 18524
rect 12389 18522 12445 18524
rect 12469 18522 12525 18524
rect 12229 18470 12255 18522
rect 12255 18470 12285 18522
rect 12309 18470 12319 18522
rect 12319 18470 12365 18522
rect 12389 18470 12435 18522
rect 12435 18470 12445 18522
rect 12469 18470 12499 18522
rect 12499 18470 12525 18522
rect 12229 18468 12285 18470
rect 12309 18468 12365 18470
rect 12389 18468 12445 18470
rect 12469 18468 12525 18470
rect 12229 17434 12285 17436
rect 12309 17434 12365 17436
rect 12389 17434 12445 17436
rect 12469 17434 12525 17436
rect 12229 17382 12255 17434
rect 12255 17382 12285 17434
rect 12309 17382 12319 17434
rect 12319 17382 12365 17434
rect 12389 17382 12435 17434
rect 12435 17382 12445 17434
rect 12469 17382 12499 17434
rect 12499 17382 12525 17434
rect 12229 17380 12285 17382
rect 12309 17380 12365 17382
rect 12389 17380 12445 17382
rect 12469 17380 12525 17382
rect 12229 16346 12285 16348
rect 12309 16346 12365 16348
rect 12389 16346 12445 16348
rect 12469 16346 12525 16348
rect 12229 16294 12255 16346
rect 12255 16294 12285 16346
rect 12309 16294 12319 16346
rect 12319 16294 12365 16346
rect 12389 16294 12435 16346
rect 12435 16294 12445 16346
rect 12469 16294 12499 16346
rect 12499 16294 12525 16346
rect 12229 16292 12285 16294
rect 12309 16292 12365 16294
rect 12389 16292 12445 16294
rect 12469 16292 12525 16294
rect 12229 15258 12285 15260
rect 12309 15258 12365 15260
rect 12389 15258 12445 15260
rect 12469 15258 12525 15260
rect 12229 15206 12255 15258
rect 12255 15206 12285 15258
rect 12309 15206 12319 15258
rect 12319 15206 12365 15258
rect 12389 15206 12435 15258
rect 12435 15206 12445 15258
rect 12469 15206 12499 15258
rect 12499 15206 12525 15258
rect 12229 15204 12285 15206
rect 12309 15204 12365 15206
rect 12389 15204 12445 15206
rect 12469 15204 12525 15206
rect 12229 14170 12285 14172
rect 12309 14170 12365 14172
rect 12389 14170 12445 14172
rect 12469 14170 12525 14172
rect 12229 14118 12255 14170
rect 12255 14118 12285 14170
rect 12309 14118 12319 14170
rect 12319 14118 12365 14170
rect 12389 14118 12435 14170
rect 12435 14118 12445 14170
rect 12469 14118 12499 14170
rect 12499 14118 12525 14170
rect 12229 14116 12285 14118
rect 12309 14116 12365 14118
rect 12389 14116 12445 14118
rect 12469 14116 12525 14118
rect 4713 11994 4769 11996
rect 4793 11994 4849 11996
rect 4873 11994 4929 11996
rect 4953 11994 5009 11996
rect 4713 11942 4739 11994
rect 4739 11942 4769 11994
rect 4793 11942 4803 11994
rect 4803 11942 4849 11994
rect 4873 11942 4919 11994
rect 4919 11942 4929 11994
rect 4953 11942 4983 11994
rect 4983 11942 5009 11994
rect 4713 11940 4769 11942
rect 4793 11940 4849 11942
rect 4873 11940 4929 11942
rect 4953 11940 5009 11942
rect 4713 10906 4769 10908
rect 4793 10906 4849 10908
rect 4873 10906 4929 10908
rect 4953 10906 5009 10908
rect 4713 10854 4739 10906
rect 4739 10854 4769 10906
rect 4793 10854 4803 10906
rect 4803 10854 4849 10906
rect 4873 10854 4919 10906
rect 4919 10854 4929 10906
rect 4953 10854 4983 10906
rect 4983 10854 5009 10906
rect 4713 10852 4769 10854
rect 4793 10852 4849 10854
rect 4873 10852 4929 10854
rect 4953 10852 5009 10854
rect 4713 9818 4769 9820
rect 4793 9818 4849 9820
rect 4873 9818 4929 9820
rect 4953 9818 5009 9820
rect 4713 9766 4739 9818
rect 4739 9766 4769 9818
rect 4793 9766 4803 9818
rect 4803 9766 4849 9818
rect 4873 9766 4919 9818
rect 4919 9766 4929 9818
rect 4953 9766 4983 9818
rect 4983 9766 5009 9818
rect 4713 9764 4769 9766
rect 4793 9764 4849 9766
rect 4873 9764 4929 9766
rect 4953 9764 5009 9766
rect 4713 8730 4769 8732
rect 4793 8730 4849 8732
rect 4873 8730 4929 8732
rect 4953 8730 5009 8732
rect 4713 8678 4739 8730
rect 4739 8678 4769 8730
rect 4793 8678 4803 8730
rect 4803 8678 4849 8730
rect 4873 8678 4919 8730
rect 4919 8678 4929 8730
rect 4953 8678 4983 8730
rect 4983 8678 5009 8730
rect 4713 8676 4769 8678
rect 4793 8676 4849 8678
rect 4873 8676 4929 8678
rect 4953 8676 5009 8678
rect 5354 7928 5410 7984
rect 4713 7642 4769 7644
rect 4793 7642 4849 7644
rect 4873 7642 4929 7644
rect 4953 7642 5009 7644
rect 4713 7590 4739 7642
rect 4739 7590 4769 7642
rect 4793 7590 4803 7642
rect 4803 7590 4849 7642
rect 4873 7590 4919 7642
rect 4919 7590 4929 7642
rect 4953 7590 4983 7642
rect 4983 7590 5009 7642
rect 4713 7588 4769 7590
rect 4793 7588 4849 7590
rect 4873 7588 4929 7590
rect 4953 7588 5009 7590
rect 5170 7404 5226 7440
rect 5170 7384 5172 7404
rect 5172 7384 5224 7404
rect 5224 7384 5226 7404
rect 4713 6554 4769 6556
rect 4793 6554 4849 6556
rect 4873 6554 4929 6556
rect 4953 6554 5009 6556
rect 4713 6502 4739 6554
rect 4739 6502 4769 6554
rect 4793 6502 4803 6554
rect 4803 6502 4849 6554
rect 4873 6502 4919 6554
rect 4919 6502 4929 6554
rect 4953 6502 4983 6554
rect 4983 6502 5009 6554
rect 4713 6500 4769 6502
rect 4793 6500 4849 6502
rect 4873 6500 4929 6502
rect 4953 6500 5009 6502
rect 4713 5466 4769 5468
rect 4793 5466 4849 5468
rect 4873 5466 4929 5468
rect 4953 5466 5009 5468
rect 4713 5414 4739 5466
rect 4739 5414 4769 5466
rect 4793 5414 4803 5466
rect 4803 5414 4849 5466
rect 4873 5414 4919 5466
rect 4919 5414 4929 5466
rect 4953 5414 4983 5466
rect 4983 5414 5009 5466
rect 4713 5412 4769 5414
rect 4793 5412 4849 5414
rect 4873 5412 4929 5414
rect 4953 5412 5009 5414
rect 4713 4378 4769 4380
rect 4793 4378 4849 4380
rect 4873 4378 4929 4380
rect 4953 4378 5009 4380
rect 4713 4326 4739 4378
rect 4739 4326 4769 4378
rect 4793 4326 4803 4378
rect 4803 4326 4849 4378
rect 4873 4326 4919 4378
rect 4919 4326 4929 4378
rect 4953 4326 4983 4378
rect 4983 4326 5009 4378
rect 4713 4324 4769 4326
rect 4793 4324 4849 4326
rect 4873 4324 4929 4326
rect 4953 4324 5009 4326
rect 5722 9460 5724 9480
rect 5724 9460 5776 9480
rect 5776 9460 5778 9480
rect 5722 9424 5778 9460
rect 4713 3290 4769 3292
rect 4793 3290 4849 3292
rect 4873 3290 4929 3292
rect 4953 3290 5009 3292
rect 4713 3238 4739 3290
rect 4739 3238 4769 3290
rect 4793 3238 4803 3290
rect 4803 3238 4849 3290
rect 4873 3238 4919 3290
rect 4919 3238 4929 3290
rect 4953 3238 4983 3290
rect 4983 3238 5009 3290
rect 4713 3236 4769 3238
rect 4793 3236 4849 3238
rect 4873 3236 4929 3238
rect 4953 3236 5009 3238
rect 4713 2202 4769 2204
rect 4793 2202 4849 2204
rect 4873 2202 4929 2204
rect 4953 2202 5009 2204
rect 4713 2150 4739 2202
rect 4739 2150 4769 2202
rect 4793 2150 4803 2202
rect 4803 2150 4849 2202
rect 4873 2150 4919 2202
rect 4919 2150 4929 2202
rect 4953 2150 4983 2202
rect 4983 2150 5009 2202
rect 4713 2148 4769 2150
rect 4793 2148 4849 2150
rect 4873 2148 4929 2150
rect 4953 2148 5009 2150
rect 6458 5208 6514 5264
rect 8471 13626 8527 13628
rect 8551 13626 8607 13628
rect 8631 13626 8687 13628
rect 8711 13626 8767 13628
rect 8471 13574 8497 13626
rect 8497 13574 8527 13626
rect 8551 13574 8561 13626
rect 8561 13574 8607 13626
rect 8631 13574 8677 13626
rect 8677 13574 8687 13626
rect 8711 13574 8741 13626
rect 8741 13574 8767 13626
rect 8471 13572 8527 13574
rect 8551 13572 8607 13574
rect 8631 13572 8687 13574
rect 8711 13572 8767 13574
rect 8471 12538 8527 12540
rect 8551 12538 8607 12540
rect 8631 12538 8687 12540
rect 8711 12538 8767 12540
rect 8471 12486 8497 12538
rect 8497 12486 8527 12538
rect 8551 12486 8561 12538
rect 8561 12486 8607 12538
rect 8631 12486 8677 12538
rect 8677 12486 8687 12538
rect 8711 12486 8741 12538
rect 8741 12486 8767 12538
rect 8471 12484 8527 12486
rect 8551 12484 8607 12486
rect 8631 12484 8687 12486
rect 8711 12484 8767 12486
rect 12229 13082 12285 13084
rect 12309 13082 12365 13084
rect 12389 13082 12445 13084
rect 12469 13082 12525 13084
rect 12229 13030 12255 13082
rect 12255 13030 12285 13082
rect 12309 13030 12319 13082
rect 12319 13030 12365 13082
rect 12389 13030 12435 13082
rect 12435 13030 12445 13082
rect 12469 13030 12499 13082
rect 12499 13030 12525 13082
rect 12229 13028 12285 13030
rect 12309 13028 12365 13030
rect 12389 13028 12445 13030
rect 12469 13028 12525 13030
rect 8471 11450 8527 11452
rect 8551 11450 8607 11452
rect 8631 11450 8687 11452
rect 8711 11450 8767 11452
rect 8471 11398 8497 11450
rect 8497 11398 8527 11450
rect 8551 11398 8561 11450
rect 8561 11398 8607 11450
rect 8631 11398 8677 11450
rect 8677 11398 8687 11450
rect 8711 11398 8741 11450
rect 8741 11398 8767 11450
rect 8471 11396 8527 11398
rect 8551 11396 8607 11398
rect 8631 11396 8687 11398
rect 8711 11396 8767 11398
rect 9954 10512 10010 10568
rect 8471 10362 8527 10364
rect 8551 10362 8607 10364
rect 8631 10362 8687 10364
rect 8711 10362 8767 10364
rect 8471 10310 8497 10362
rect 8497 10310 8527 10362
rect 8551 10310 8561 10362
rect 8561 10310 8607 10362
rect 8631 10310 8677 10362
rect 8677 10310 8687 10362
rect 8711 10310 8741 10362
rect 8741 10310 8767 10362
rect 8471 10308 8527 10310
rect 8551 10308 8607 10310
rect 8631 10308 8687 10310
rect 8711 10308 8767 10310
rect 8471 9274 8527 9276
rect 8551 9274 8607 9276
rect 8631 9274 8687 9276
rect 8711 9274 8767 9276
rect 8471 9222 8497 9274
rect 8497 9222 8527 9274
rect 8551 9222 8561 9274
rect 8561 9222 8607 9274
rect 8631 9222 8677 9274
rect 8677 9222 8687 9274
rect 8711 9222 8741 9274
rect 8741 9222 8767 9274
rect 8471 9220 8527 9222
rect 8551 9220 8607 9222
rect 8631 9220 8687 9222
rect 8711 9220 8767 9222
rect 8471 8186 8527 8188
rect 8551 8186 8607 8188
rect 8631 8186 8687 8188
rect 8711 8186 8767 8188
rect 8471 8134 8497 8186
rect 8497 8134 8527 8186
rect 8551 8134 8561 8186
rect 8561 8134 8607 8186
rect 8631 8134 8677 8186
rect 8677 8134 8687 8186
rect 8711 8134 8741 8186
rect 8741 8134 8767 8186
rect 8471 8132 8527 8134
rect 8551 8132 8607 8134
rect 8631 8132 8687 8134
rect 8711 8132 8767 8134
rect 8471 7098 8527 7100
rect 8551 7098 8607 7100
rect 8631 7098 8687 7100
rect 8711 7098 8767 7100
rect 8471 7046 8497 7098
rect 8497 7046 8527 7098
rect 8551 7046 8561 7098
rect 8561 7046 8607 7098
rect 8631 7046 8677 7098
rect 8677 7046 8687 7098
rect 8711 7046 8741 7098
rect 8741 7046 8767 7098
rect 8471 7044 8527 7046
rect 8551 7044 8607 7046
rect 8631 7044 8687 7046
rect 8711 7044 8767 7046
rect 8471 6010 8527 6012
rect 8551 6010 8607 6012
rect 8631 6010 8687 6012
rect 8711 6010 8767 6012
rect 8471 5958 8497 6010
rect 8497 5958 8527 6010
rect 8551 5958 8561 6010
rect 8561 5958 8607 6010
rect 8631 5958 8677 6010
rect 8677 5958 8687 6010
rect 8711 5958 8741 6010
rect 8741 5958 8767 6010
rect 8471 5956 8527 5958
rect 8551 5956 8607 5958
rect 8631 5956 8687 5958
rect 8711 5956 8767 5958
rect 8471 4922 8527 4924
rect 8551 4922 8607 4924
rect 8631 4922 8687 4924
rect 8711 4922 8767 4924
rect 8471 4870 8497 4922
rect 8497 4870 8527 4922
rect 8551 4870 8561 4922
rect 8561 4870 8607 4922
rect 8631 4870 8677 4922
rect 8677 4870 8687 4922
rect 8711 4870 8741 4922
rect 8741 4870 8767 4922
rect 8471 4868 8527 4870
rect 8551 4868 8607 4870
rect 8631 4868 8687 4870
rect 8711 4868 8767 4870
rect 8298 4120 8354 4176
rect 8390 3984 8446 4040
rect 8471 3834 8527 3836
rect 8551 3834 8607 3836
rect 8631 3834 8687 3836
rect 8711 3834 8767 3836
rect 8471 3782 8497 3834
rect 8497 3782 8527 3834
rect 8551 3782 8561 3834
rect 8561 3782 8607 3834
rect 8631 3782 8677 3834
rect 8677 3782 8687 3834
rect 8711 3782 8741 3834
rect 8741 3782 8767 3834
rect 8471 3780 8527 3782
rect 8551 3780 8607 3782
rect 8631 3780 8687 3782
rect 8711 3780 8767 3782
rect 8471 2746 8527 2748
rect 8551 2746 8607 2748
rect 8631 2746 8687 2748
rect 8711 2746 8767 2748
rect 8471 2694 8497 2746
rect 8497 2694 8527 2746
rect 8551 2694 8561 2746
rect 8561 2694 8607 2746
rect 8631 2694 8677 2746
rect 8677 2694 8687 2746
rect 8711 2694 8741 2746
rect 8741 2694 8767 2746
rect 8471 2692 8527 2694
rect 8551 2692 8607 2694
rect 8631 2692 8687 2694
rect 8711 2692 8767 2694
rect 12229 11994 12285 11996
rect 12309 11994 12365 11996
rect 12389 11994 12445 11996
rect 12469 11994 12525 11996
rect 12229 11942 12255 11994
rect 12255 11942 12285 11994
rect 12309 11942 12319 11994
rect 12319 11942 12365 11994
rect 12389 11942 12435 11994
rect 12435 11942 12445 11994
rect 12469 11942 12499 11994
rect 12499 11942 12525 11994
rect 12229 11940 12285 11942
rect 12309 11940 12365 11942
rect 12389 11940 12445 11942
rect 12469 11940 12525 11942
rect 12229 10906 12285 10908
rect 12309 10906 12365 10908
rect 12389 10906 12445 10908
rect 12469 10906 12525 10908
rect 12229 10854 12255 10906
rect 12255 10854 12285 10906
rect 12309 10854 12319 10906
rect 12319 10854 12365 10906
rect 12389 10854 12435 10906
rect 12435 10854 12445 10906
rect 12469 10854 12499 10906
rect 12499 10854 12525 10906
rect 12229 10852 12285 10854
rect 12309 10852 12365 10854
rect 12389 10852 12445 10854
rect 12469 10852 12525 10854
rect 12229 9818 12285 9820
rect 12309 9818 12365 9820
rect 12389 9818 12445 9820
rect 12469 9818 12525 9820
rect 12229 9766 12255 9818
rect 12255 9766 12285 9818
rect 12309 9766 12319 9818
rect 12319 9766 12365 9818
rect 12389 9766 12435 9818
rect 12435 9766 12445 9818
rect 12469 9766 12499 9818
rect 12499 9766 12525 9818
rect 12229 9764 12285 9766
rect 12309 9764 12365 9766
rect 12389 9764 12445 9766
rect 12469 9764 12525 9766
rect 10966 7248 11022 7304
rect 11334 1400 11390 1456
rect 14278 10512 14334 10568
rect 15986 22330 16042 22332
rect 16066 22330 16122 22332
rect 16146 22330 16202 22332
rect 16226 22330 16282 22332
rect 15986 22278 16012 22330
rect 16012 22278 16042 22330
rect 16066 22278 16076 22330
rect 16076 22278 16122 22330
rect 16146 22278 16192 22330
rect 16192 22278 16202 22330
rect 16226 22278 16256 22330
rect 16256 22278 16282 22330
rect 15986 22276 16042 22278
rect 16066 22276 16122 22278
rect 16146 22276 16202 22278
rect 16226 22276 16282 22278
rect 15986 21242 16042 21244
rect 16066 21242 16122 21244
rect 16146 21242 16202 21244
rect 16226 21242 16282 21244
rect 15986 21190 16012 21242
rect 16012 21190 16042 21242
rect 16066 21190 16076 21242
rect 16076 21190 16122 21242
rect 16146 21190 16192 21242
rect 16192 21190 16202 21242
rect 16226 21190 16256 21242
rect 16256 21190 16282 21242
rect 15986 21188 16042 21190
rect 16066 21188 16122 21190
rect 16146 21188 16202 21190
rect 16226 21188 16282 21190
rect 15986 20154 16042 20156
rect 16066 20154 16122 20156
rect 16146 20154 16202 20156
rect 16226 20154 16282 20156
rect 15986 20102 16012 20154
rect 16012 20102 16042 20154
rect 16066 20102 16076 20154
rect 16076 20102 16122 20154
rect 16146 20102 16192 20154
rect 16192 20102 16202 20154
rect 16226 20102 16256 20154
rect 16256 20102 16282 20154
rect 15986 20100 16042 20102
rect 16066 20100 16122 20102
rect 16146 20100 16202 20102
rect 16226 20100 16282 20102
rect 15986 19066 16042 19068
rect 16066 19066 16122 19068
rect 16146 19066 16202 19068
rect 16226 19066 16282 19068
rect 15986 19014 16012 19066
rect 16012 19014 16042 19066
rect 16066 19014 16076 19066
rect 16076 19014 16122 19066
rect 16146 19014 16192 19066
rect 16192 19014 16202 19066
rect 16226 19014 16256 19066
rect 16256 19014 16282 19066
rect 15986 19012 16042 19014
rect 16066 19012 16122 19014
rect 16146 19012 16202 19014
rect 16226 19012 16282 19014
rect 15986 17978 16042 17980
rect 16066 17978 16122 17980
rect 16146 17978 16202 17980
rect 16226 17978 16282 17980
rect 15986 17926 16012 17978
rect 16012 17926 16042 17978
rect 16066 17926 16076 17978
rect 16076 17926 16122 17978
rect 16146 17926 16192 17978
rect 16192 17926 16202 17978
rect 16226 17926 16256 17978
rect 16256 17926 16282 17978
rect 15986 17924 16042 17926
rect 16066 17924 16122 17926
rect 16146 17924 16202 17926
rect 16226 17924 16282 17926
rect 15986 16890 16042 16892
rect 16066 16890 16122 16892
rect 16146 16890 16202 16892
rect 16226 16890 16282 16892
rect 15986 16838 16012 16890
rect 16012 16838 16042 16890
rect 16066 16838 16076 16890
rect 16076 16838 16122 16890
rect 16146 16838 16192 16890
rect 16192 16838 16202 16890
rect 16226 16838 16256 16890
rect 16256 16838 16282 16890
rect 15986 16836 16042 16838
rect 16066 16836 16122 16838
rect 16146 16836 16202 16838
rect 16226 16836 16282 16838
rect 15474 16496 15530 16552
rect 15986 15802 16042 15804
rect 16066 15802 16122 15804
rect 16146 15802 16202 15804
rect 16226 15802 16282 15804
rect 15986 15750 16012 15802
rect 16012 15750 16042 15802
rect 16066 15750 16076 15802
rect 16076 15750 16122 15802
rect 16146 15750 16192 15802
rect 16192 15750 16202 15802
rect 16226 15750 16256 15802
rect 16256 15750 16282 15802
rect 15986 15748 16042 15750
rect 16066 15748 16122 15750
rect 16146 15748 16202 15750
rect 16226 15748 16282 15750
rect 15986 14714 16042 14716
rect 16066 14714 16122 14716
rect 16146 14714 16202 14716
rect 16226 14714 16282 14716
rect 15986 14662 16012 14714
rect 16012 14662 16042 14714
rect 16066 14662 16076 14714
rect 16076 14662 16122 14714
rect 16146 14662 16192 14714
rect 16192 14662 16202 14714
rect 16226 14662 16256 14714
rect 16256 14662 16282 14714
rect 15986 14660 16042 14662
rect 16066 14660 16122 14662
rect 16146 14660 16202 14662
rect 16226 14660 16282 14662
rect 15986 13626 16042 13628
rect 16066 13626 16122 13628
rect 16146 13626 16202 13628
rect 16226 13626 16282 13628
rect 15986 13574 16012 13626
rect 16012 13574 16042 13626
rect 16066 13574 16076 13626
rect 16076 13574 16122 13626
rect 16146 13574 16192 13626
rect 16192 13574 16202 13626
rect 16226 13574 16256 13626
rect 16256 13574 16282 13626
rect 15986 13572 16042 13574
rect 16066 13572 16122 13574
rect 16146 13572 16202 13574
rect 16226 13572 16282 13574
rect 15986 12538 16042 12540
rect 16066 12538 16122 12540
rect 16146 12538 16202 12540
rect 16226 12538 16282 12540
rect 15986 12486 16012 12538
rect 16012 12486 16042 12538
rect 16066 12486 16076 12538
rect 16076 12486 16122 12538
rect 16146 12486 16192 12538
rect 16192 12486 16202 12538
rect 16226 12486 16256 12538
rect 16256 12486 16282 12538
rect 15986 12484 16042 12486
rect 16066 12484 16122 12486
rect 16146 12484 16202 12486
rect 16226 12484 16282 12486
rect 15986 11450 16042 11452
rect 16066 11450 16122 11452
rect 16146 11450 16202 11452
rect 16226 11450 16282 11452
rect 15986 11398 16012 11450
rect 16012 11398 16042 11450
rect 16066 11398 16076 11450
rect 16076 11398 16122 11450
rect 16146 11398 16192 11450
rect 16192 11398 16202 11450
rect 16226 11398 16256 11450
rect 16256 11398 16282 11450
rect 15986 11396 16042 11398
rect 16066 11396 16122 11398
rect 16146 11396 16202 11398
rect 16226 11396 16282 11398
rect 15986 10362 16042 10364
rect 16066 10362 16122 10364
rect 16146 10362 16202 10364
rect 16226 10362 16282 10364
rect 15986 10310 16012 10362
rect 16012 10310 16042 10362
rect 16066 10310 16076 10362
rect 16076 10310 16122 10362
rect 16146 10310 16192 10362
rect 16192 10310 16202 10362
rect 16226 10310 16256 10362
rect 16256 10310 16282 10362
rect 15986 10308 16042 10310
rect 16066 10308 16122 10310
rect 16146 10308 16202 10310
rect 16226 10308 16282 10310
rect 13358 9424 13414 9480
rect 12229 8730 12285 8732
rect 12309 8730 12365 8732
rect 12389 8730 12445 8732
rect 12469 8730 12525 8732
rect 12229 8678 12255 8730
rect 12255 8678 12285 8730
rect 12309 8678 12319 8730
rect 12319 8678 12365 8730
rect 12389 8678 12435 8730
rect 12435 8678 12445 8730
rect 12469 8678 12499 8730
rect 12499 8678 12525 8730
rect 12229 8676 12285 8678
rect 12309 8676 12365 8678
rect 12389 8676 12445 8678
rect 12469 8676 12525 8678
rect 12229 7642 12285 7644
rect 12309 7642 12365 7644
rect 12389 7642 12445 7644
rect 12469 7642 12525 7644
rect 12229 7590 12255 7642
rect 12255 7590 12285 7642
rect 12309 7590 12319 7642
rect 12319 7590 12365 7642
rect 12389 7590 12435 7642
rect 12435 7590 12445 7642
rect 12469 7590 12499 7642
rect 12499 7590 12525 7642
rect 12229 7588 12285 7590
rect 12309 7588 12365 7590
rect 12389 7588 12445 7590
rect 12469 7588 12525 7590
rect 14646 9424 14702 9480
rect 15986 9274 16042 9276
rect 16066 9274 16122 9276
rect 16146 9274 16202 9276
rect 16226 9274 16282 9276
rect 15986 9222 16012 9274
rect 16012 9222 16042 9274
rect 16066 9222 16076 9274
rect 16076 9222 16122 9274
rect 16146 9222 16192 9274
rect 16192 9222 16202 9274
rect 16226 9222 16256 9274
rect 16256 9222 16282 9274
rect 15986 9220 16042 9222
rect 16066 9220 16122 9222
rect 16146 9220 16202 9222
rect 16226 9220 16282 9222
rect 15986 8186 16042 8188
rect 16066 8186 16122 8188
rect 16146 8186 16202 8188
rect 16226 8186 16282 8188
rect 15986 8134 16012 8186
rect 16012 8134 16042 8186
rect 16066 8134 16076 8186
rect 16076 8134 16122 8186
rect 16146 8134 16192 8186
rect 16192 8134 16202 8186
rect 16226 8134 16256 8186
rect 16256 8134 16282 8186
rect 15986 8132 16042 8134
rect 16066 8132 16122 8134
rect 16146 8132 16202 8134
rect 16226 8132 16282 8134
rect 15986 7098 16042 7100
rect 16066 7098 16122 7100
rect 16146 7098 16202 7100
rect 16226 7098 16282 7100
rect 15986 7046 16012 7098
rect 16012 7046 16042 7098
rect 16066 7046 16076 7098
rect 16076 7046 16122 7098
rect 16146 7046 16192 7098
rect 16192 7046 16202 7098
rect 16226 7046 16256 7098
rect 16256 7046 16282 7098
rect 15986 7044 16042 7046
rect 16066 7044 16122 7046
rect 16146 7044 16202 7046
rect 16226 7044 16282 7046
rect 12229 6554 12285 6556
rect 12309 6554 12365 6556
rect 12389 6554 12445 6556
rect 12469 6554 12525 6556
rect 12229 6502 12255 6554
rect 12255 6502 12285 6554
rect 12309 6502 12319 6554
rect 12319 6502 12365 6554
rect 12389 6502 12435 6554
rect 12435 6502 12445 6554
rect 12469 6502 12499 6554
rect 12499 6502 12525 6554
rect 12229 6500 12285 6502
rect 12309 6500 12365 6502
rect 12389 6500 12445 6502
rect 12469 6500 12525 6502
rect 16946 6296 17002 6352
rect 12229 5466 12285 5468
rect 12309 5466 12365 5468
rect 12389 5466 12445 5468
rect 12469 5466 12525 5468
rect 12229 5414 12255 5466
rect 12255 5414 12285 5466
rect 12309 5414 12319 5466
rect 12319 5414 12365 5466
rect 12389 5414 12435 5466
rect 12435 5414 12445 5466
rect 12469 5414 12499 5466
rect 12499 5414 12525 5466
rect 12229 5412 12285 5414
rect 12309 5412 12365 5414
rect 12389 5412 12445 5414
rect 12469 5412 12525 5414
rect 12229 4378 12285 4380
rect 12309 4378 12365 4380
rect 12389 4378 12445 4380
rect 12469 4378 12525 4380
rect 12229 4326 12255 4378
rect 12255 4326 12285 4378
rect 12309 4326 12319 4378
rect 12319 4326 12365 4378
rect 12389 4326 12435 4378
rect 12435 4326 12445 4378
rect 12469 4326 12499 4378
rect 12499 4326 12525 4378
rect 12229 4324 12285 4326
rect 12309 4324 12365 4326
rect 12389 4324 12445 4326
rect 12469 4324 12525 4326
rect 11978 3576 12034 3632
rect 12229 3290 12285 3292
rect 12309 3290 12365 3292
rect 12389 3290 12445 3292
rect 12469 3290 12525 3292
rect 12229 3238 12255 3290
rect 12255 3238 12285 3290
rect 12309 3238 12319 3290
rect 12319 3238 12365 3290
rect 12389 3238 12435 3290
rect 12435 3238 12445 3290
rect 12469 3238 12499 3290
rect 12499 3238 12525 3290
rect 12229 3236 12285 3238
rect 12309 3236 12365 3238
rect 12389 3236 12445 3238
rect 12469 3236 12525 3238
rect 12229 2202 12285 2204
rect 12309 2202 12365 2204
rect 12389 2202 12445 2204
rect 12469 2202 12525 2204
rect 12229 2150 12255 2202
rect 12255 2150 12285 2202
rect 12309 2150 12319 2202
rect 12319 2150 12365 2202
rect 12389 2150 12435 2202
rect 12435 2150 12445 2202
rect 12469 2150 12499 2202
rect 12499 2150 12525 2202
rect 12229 2148 12285 2150
rect 12309 2148 12365 2150
rect 12389 2148 12445 2150
rect 12469 2148 12525 2150
rect 15986 6010 16042 6012
rect 16066 6010 16122 6012
rect 16146 6010 16202 6012
rect 16226 6010 16282 6012
rect 15986 5958 16012 6010
rect 16012 5958 16042 6010
rect 16066 5958 16076 6010
rect 16076 5958 16122 6010
rect 16146 5958 16192 6010
rect 16192 5958 16202 6010
rect 16226 5958 16256 6010
rect 16256 5958 16282 6010
rect 15986 5956 16042 5958
rect 16066 5956 16122 5958
rect 16146 5956 16202 5958
rect 16226 5956 16282 5958
rect 17590 23568 17646 23624
rect 19154 22480 19210 22536
rect 19522 22072 19578 22128
rect 18970 19760 19026 19816
rect 19744 21786 19800 21788
rect 19824 21786 19880 21788
rect 19904 21786 19960 21788
rect 19984 21786 20040 21788
rect 19744 21734 19770 21786
rect 19770 21734 19800 21786
rect 19824 21734 19834 21786
rect 19834 21734 19880 21786
rect 19904 21734 19950 21786
rect 19950 21734 19960 21786
rect 19984 21734 20014 21786
rect 20014 21734 20040 21786
rect 19744 21732 19800 21734
rect 19824 21732 19880 21734
rect 19904 21732 19960 21734
rect 19984 21732 20040 21734
rect 19744 20698 19800 20700
rect 19824 20698 19880 20700
rect 19904 20698 19960 20700
rect 19984 20698 20040 20700
rect 19744 20646 19770 20698
rect 19770 20646 19800 20698
rect 19824 20646 19834 20698
rect 19834 20646 19880 20698
rect 19904 20646 19950 20698
rect 19950 20646 19960 20698
rect 19984 20646 20014 20698
rect 20014 20646 20040 20698
rect 19744 20644 19800 20646
rect 19824 20644 19880 20646
rect 19904 20644 19960 20646
rect 19984 20644 20040 20646
rect 19522 20440 19578 20496
rect 19744 19610 19800 19612
rect 19824 19610 19880 19612
rect 19904 19610 19960 19612
rect 19984 19610 20040 19612
rect 19744 19558 19770 19610
rect 19770 19558 19800 19610
rect 19824 19558 19834 19610
rect 19834 19558 19880 19610
rect 19904 19558 19950 19610
rect 19950 19558 19960 19610
rect 19984 19558 20014 19610
rect 20014 19558 20040 19610
rect 19744 19556 19800 19558
rect 19824 19556 19880 19558
rect 19904 19556 19960 19558
rect 19984 19556 20040 19558
rect 19614 19216 19670 19272
rect 17498 15408 17554 15464
rect 16302 5208 16358 5264
rect 15986 4922 16042 4924
rect 16066 4922 16122 4924
rect 16146 4922 16202 4924
rect 16226 4922 16282 4924
rect 15986 4870 16012 4922
rect 16012 4870 16042 4922
rect 16066 4870 16076 4922
rect 16076 4870 16122 4922
rect 16146 4870 16192 4922
rect 16192 4870 16202 4922
rect 16226 4870 16256 4922
rect 16256 4870 16282 4922
rect 15986 4868 16042 4870
rect 16066 4868 16122 4870
rect 16146 4868 16202 4870
rect 16226 4868 16282 4870
rect 15986 3834 16042 3836
rect 16066 3834 16122 3836
rect 16146 3834 16202 3836
rect 16226 3834 16282 3836
rect 15986 3782 16012 3834
rect 16012 3782 16042 3834
rect 16066 3782 16076 3834
rect 16076 3782 16122 3834
rect 16146 3782 16192 3834
rect 16192 3782 16202 3834
rect 16226 3782 16256 3834
rect 16256 3782 16282 3834
rect 15986 3780 16042 3782
rect 16066 3780 16122 3782
rect 16146 3780 16202 3782
rect 16226 3780 16282 3782
rect 15986 2746 16042 2748
rect 16066 2746 16122 2748
rect 16146 2746 16202 2748
rect 16226 2746 16282 2748
rect 15986 2694 16012 2746
rect 16012 2694 16042 2746
rect 16066 2694 16076 2746
rect 16076 2694 16122 2746
rect 16146 2694 16192 2746
rect 16192 2694 16202 2746
rect 16226 2694 16256 2746
rect 16256 2694 16282 2746
rect 15986 2692 16042 2694
rect 16066 2692 16122 2694
rect 16146 2692 16202 2694
rect 16226 2692 16282 2694
rect 19430 17584 19486 17640
rect 18602 7928 18658 7984
rect 20166 19216 20222 19272
rect 19744 18522 19800 18524
rect 19824 18522 19880 18524
rect 19904 18522 19960 18524
rect 19984 18522 20040 18524
rect 19744 18470 19770 18522
rect 19770 18470 19800 18522
rect 19824 18470 19834 18522
rect 19834 18470 19880 18522
rect 19904 18470 19950 18522
rect 19950 18470 19960 18522
rect 19984 18470 20014 18522
rect 20014 18470 20040 18522
rect 19744 18468 19800 18470
rect 19824 18468 19880 18470
rect 19904 18468 19960 18470
rect 19984 18468 20040 18470
rect 19744 17434 19800 17436
rect 19824 17434 19880 17436
rect 19904 17434 19960 17436
rect 19984 17434 20040 17436
rect 19744 17382 19770 17434
rect 19770 17382 19800 17434
rect 19824 17382 19834 17434
rect 19834 17382 19880 17434
rect 19904 17382 19950 17434
rect 19950 17382 19960 17434
rect 19984 17382 20014 17434
rect 20014 17382 20040 17434
rect 19744 17380 19800 17382
rect 19824 17380 19880 17382
rect 19904 17380 19960 17382
rect 19984 17380 20040 17382
rect 19744 16346 19800 16348
rect 19824 16346 19880 16348
rect 19904 16346 19960 16348
rect 19984 16346 20040 16348
rect 19744 16294 19770 16346
rect 19770 16294 19800 16346
rect 19824 16294 19834 16346
rect 19834 16294 19880 16346
rect 19904 16294 19950 16346
rect 19950 16294 19960 16346
rect 19984 16294 20014 16346
rect 20014 16294 20040 16346
rect 19744 16292 19800 16294
rect 19824 16292 19880 16294
rect 19904 16292 19960 16294
rect 19984 16292 20040 16294
rect 19744 15258 19800 15260
rect 19824 15258 19880 15260
rect 19904 15258 19960 15260
rect 19984 15258 20040 15260
rect 19744 15206 19770 15258
rect 19770 15206 19800 15258
rect 19824 15206 19834 15258
rect 19834 15206 19880 15258
rect 19904 15206 19950 15258
rect 19950 15206 19960 15258
rect 19984 15206 20014 15258
rect 20014 15206 20040 15258
rect 19744 15204 19800 15206
rect 19824 15204 19880 15206
rect 19904 15204 19960 15206
rect 19984 15204 20040 15206
rect 19744 14170 19800 14172
rect 19824 14170 19880 14172
rect 19904 14170 19960 14172
rect 19984 14170 20040 14172
rect 19744 14118 19770 14170
rect 19770 14118 19800 14170
rect 19824 14118 19834 14170
rect 19834 14118 19880 14170
rect 19904 14118 19950 14170
rect 19950 14118 19960 14170
rect 19984 14118 20014 14170
rect 20014 14118 20040 14170
rect 19744 14116 19800 14118
rect 19824 14116 19880 14118
rect 19904 14116 19960 14118
rect 19984 14116 20040 14118
rect 19744 13082 19800 13084
rect 19824 13082 19880 13084
rect 19904 13082 19960 13084
rect 19984 13082 20040 13084
rect 19744 13030 19770 13082
rect 19770 13030 19800 13082
rect 19824 13030 19834 13082
rect 19834 13030 19880 13082
rect 19904 13030 19950 13082
rect 19950 13030 19960 13082
rect 19984 13030 20014 13082
rect 20014 13030 20040 13082
rect 19744 13028 19800 13030
rect 19824 13028 19880 13030
rect 19904 13028 19960 13030
rect 19984 13028 20040 13030
rect 19744 11994 19800 11996
rect 19824 11994 19880 11996
rect 19904 11994 19960 11996
rect 19984 11994 20040 11996
rect 19744 11942 19770 11994
rect 19770 11942 19800 11994
rect 19824 11942 19834 11994
rect 19834 11942 19880 11994
rect 19904 11942 19950 11994
rect 19950 11942 19960 11994
rect 19984 11942 20014 11994
rect 20014 11942 20040 11994
rect 19744 11940 19800 11942
rect 19824 11940 19880 11942
rect 19904 11940 19960 11942
rect 19984 11940 20040 11942
rect 19744 10906 19800 10908
rect 19824 10906 19880 10908
rect 19904 10906 19960 10908
rect 19984 10906 20040 10908
rect 19744 10854 19770 10906
rect 19770 10854 19800 10906
rect 19824 10854 19834 10906
rect 19834 10854 19880 10906
rect 19904 10854 19950 10906
rect 19950 10854 19960 10906
rect 19984 10854 20014 10906
rect 20014 10854 20040 10906
rect 19744 10852 19800 10854
rect 19824 10852 19880 10854
rect 19904 10852 19960 10854
rect 19984 10852 20040 10854
rect 22098 18944 22154 19000
rect 22098 17176 22154 17232
rect 22098 13776 22154 13832
rect 21086 13096 21142 13152
rect 20166 11192 20222 11248
rect 19744 9818 19800 9820
rect 19824 9818 19880 9820
rect 19904 9818 19960 9820
rect 19984 9818 20040 9820
rect 19744 9766 19770 9818
rect 19770 9766 19800 9818
rect 19824 9766 19834 9818
rect 19834 9766 19880 9818
rect 19904 9766 19950 9818
rect 19950 9766 19960 9818
rect 19984 9766 20014 9818
rect 20014 9766 20040 9818
rect 19744 9764 19800 9766
rect 19824 9764 19880 9766
rect 19904 9764 19960 9766
rect 19984 9764 20040 9766
rect 20166 9288 20222 9344
rect 19744 8730 19800 8732
rect 19824 8730 19880 8732
rect 19904 8730 19960 8732
rect 19984 8730 20040 8732
rect 19744 8678 19770 8730
rect 19770 8678 19800 8730
rect 19824 8678 19834 8730
rect 19834 8678 19880 8730
rect 19904 8678 19950 8730
rect 19950 8678 19960 8730
rect 19984 8678 20014 8730
rect 20014 8678 20040 8730
rect 19744 8676 19800 8678
rect 19824 8676 19880 8678
rect 19904 8676 19960 8678
rect 19984 8676 20040 8678
rect 20166 8608 20222 8664
rect 19744 7642 19800 7644
rect 19824 7642 19880 7644
rect 19904 7642 19960 7644
rect 19984 7642 20040 7644
rect 19744 7590 19770 7642
rect 19770 7590 19800 7642
rect 19824 7590 19834 7642
rect 19834 7590 19880 7642
rect 19904 7590 19950 7642
rect 19950 7590 19960 7642
rect 19984 7590 20014 7642
rect 20014 7590 20040 7642
rect 19744 7588 19800 7590
rect 19824 7588 19880 7590
rect 19904 7588 19960 7590
rect 19984 7588 20040 7590
rect 19744 6554 19800 6556
rect 19824 6554 19880 6556
rect 19904 6554 19960 6556
rect 19984 6554 20040 6556
rect 19744 6502 19770 6554
rect 19770 6502 19800 6554
rect 19824 6502 19834 6554
rect 19834 6502 19880 6554
rect 19904 6502 19950 6554
rect 19950 6502 19960 6554
rect 19984 6502 20014 6554
rect 20014 6502 20040 6554
rect 19744 6500 19800 6502
rect 19824 6500 19880 6502
rect 19904 6500 19960 6502
rect 19984 6500 20040 6502
rect 20166 5480 20222 5536
rect 19744 5466 19800 5468
rect 19824 5466 19880 5468
rect 19904 5466 19960 5468
rect 19984 5466 20040 5468
rect 19744 5414 19770 5466
rect 19770 5414 19800 5466
rect 19824 5414 19834 5466
rect 19834 5414 19880 5466
rect 19904 5414 19950 5466
rect 19950 5414 19960 5466
rect 19984 5414 20014 5466
rect 20014 5414 20040 5466
rect 19744 5412 19800 5414
rect 19824 5412 19880 5414
rect 19904 5412 19960 5414
rect 19984 5412 20040 5414
rect 20258 5072 20314 5128
rect 19744 4378 19800 4380
rect 19824 4378 19880 4380
rect 19904 4378 19960 4380
rect 19984 4378 20040 4380
rect 19744 4326 19770 4378
rect 19770 4326 19800 4378
rect 19824 4326 19834 4378
rect 19834 4326 19880 4378
rect 19904 4326 19950 4378
rect 19950 4326 19960 4378
rect 19984 4326 20014 4378
rect 20014 4326 20040 4378
rect 19744 4324 19800 4326
rect 19824 4324 19880 4326
rect 19904 4324 19960 4326
rect 19984 4324 20040 4326
rect 20074 3984 20130 4040
rect 19744 3290 19800 3292
rect 19824 3290 19880 3292
rect 19904 3290 19960 3292
rect 19984 3290 20040 3292
rect 19744 3238 19770 3290
rect 19770 3238 19800 3290
rect 19824 3238 19834 3290
rect 19834 3238 19880 3290
rect 19904 3238 19950 3290
rect 19950 3238 19960 3290
rect 19984 3238 20014 3290
rect 20014 3238 20040 3290
rect 19744 3236 19800 3238
rect 19824 3236 19880 3238
rect 19904 3236 19960 3238
rect 19984 3236 20040 3238
rect 19744 2202 19800 2204
rect 19824 2202 19880 2204
rect 19904 2202 19960 2204
rect 19984 2202 20040 2204
rect 19744 2150 19770 2202
rect 19770 2150 19800 2202
rect 19824 2150 19834 2202
rect 19834 2150 19880 2202
rect 19904 2150 19950 2202
rect 19950 2150 19960 2202
rect 19984 2150 20014 2202
rect 20014 2150 20040 2202
rect 19744 2148 19800 2150
rect 19824 2148 19880 2150
rect 19904 2148 19960 2150
rect 19984 2148 20040 2150
<< metal3 >>
rect 22066 24080 22546 24200
rect 0 23944 480 24064
rect 62 23490 122 23944
rect 17585 23626 17651 23629
rect 22142 23626 22202 24080
rect 17585 23624 22202 23626
rect 17585 23568 17590 23624
rect 17646 23568 22202 23624
rect 17585 23566 22202 23568
rect 17585 23563 17651 23566
rect 1301 23490 1367 23493
rect 62 23488 1367 23490
rect 62 23432 1306 23488
rect 1362 23432 1367 23488
rect 62 23430 1367 23432
rect 1301 23427 1367 23430
rect 22066 22992 22546 23112
rect 0 22808 480 22840
rect 0 22752 110 22808
rect 166 22752 480 22808
rect 0 22720 480 22752
rect 19149 22538 19215 22541
rect 22142 22538 22202 22992
rect 19149 22536 22202 22538
rect 19149 22480 19154 22536
rect 19210 22480 22202 22536
rect 19149 22478 22202 22480
rect 19149 22475 19215 22478
rect 8459 22336 8779 22337
rect 8459 22272 8467 22336
rect 8531 22272 8547 22336
rect 8611 22272 8627 22336
rect 8691 22272 8707 22336
rect 8771 22272 8779 22336
rect 8459 22271 8779 22272
rect 15974 22336 16294 22337
rect 15974 22272 15982 22336
rect 16046 22272 16062 22336
rect 16126 22272 16142 22336
rect 16206 22272 16222 22336
rect 16286 22272 16294 22336
rect 15974 22271 16294 22272
rect 19517 22130 19583 22133
rect 22066 22130 22546 22160
rect 19517 22128 22546 22130
rect 19517 22072 19522 22128
rect 19578 22072 22546 22128
rect 19517 22070 22546 22072
rect 19517 22067 19583 22070
rect 22066 22040 22546 22070
rect 4701 21792 5021 21793
rect 4701 21728 4709 21792
rect 4773 21728 4789 21792
rect 4853 21728 4869 21792
rect 4933 21728 4949 21792
rect 5013 21728 5021 21792
rect 4701 21727 5021 21728
rect 12217 21792 12537 21793
rect 12217 21728 12225 21792
rect 12289 21728 12305 21792
rect 12369 21728 12385 21792
rect 12449 21728 12465 21792
rect 12529 21728 12537 21792
rect 12217 21727 12537 21728
rect 19732 21792 20052 21793
rect 19732 21728 19740 21792
rect 19804 21728 19820 21792
rect 19884 21728 19900 21792
rect 19964 21728 19980 21792
rect 20044 21728 20052 21792
rect 19732 21727 20052 21728
rect 0 21496 480 21616
rect 62 21042 122 21496
rect 8459 21248 8779 21249
rect 8459 21184 8467 21248
rect 8531 21184 8547 21248
rect 8611 21184 8627 21248
rect 8691 21184 8707 21248
rect 8771 21184 8779 21248
rect 8459 21183 8779 21184
rect 15974 21248 16294 21249
rect 15974 21184 15982 21248
rect 16046 21184 16062 21248
rect 16126 21184 16142 21248
rect 16206 21184 16222 21248
rect 16286 21184 16294 21248
rect 15974 21183 16294 21184
rect 3509 21042 3575 21045
rect 62 21040 3575 21042
rect 62 20984 3514 21040
rect 3570 20984 3575 21040
rect 62 20982 3575 20984
rect 3509 20979 3575 20982
rect 22066 20952 22546 21072
rect 4701 20704 5021 20705
rect 4701 20640 4709 20704
rect 4773 20640 4789 20704
rect 4853 20640 4869 20704
rect 4933 20640 4949 20704
rect 5013 20640 5021 20704
rect 4701 20639 5021 20640
rect 12217 20704 12537 20705
rect 12217 20640 12225 20704
rect 12289 20640 12305 20704
rect 12369 20640 12385 20704
rect 12449 20640 12465 20704
rect 12529 20640 12537 20704
rect 12217 20639 12537 20640
rect 19732 20704 20052 20705
rect 19732 20640 19740 20704
rect 19804 20640 19820 20704
rect 19884 20640 19900 20704
rect 19964 20640 19980 20704
rect 20044 20640 20052 20704
rect 19732 20639 20052 20640
rect 19517 20498 19583 20501
rect 22142 20498 22202 20952
rect 19517 20496 22202 20498
rect 19517 20440 19522 20496
rect 19578 20440 22202 20496
rect 19517 20438 22202 20440
rect 19517 20435 19583 20438
rect 0 20272 480 20392
rect 62 19818 122 20272
rect 8459 20160 8779 20161
rect 8459 20096 8467 20160
rect 8531 20096 8547 20160
rect 8611 20096 8627 20160
rect 8691 20096 8707 20160
rect 8771 20096 8779 20160
rect 8459 20095 8779 20096
rect 15974 20160 16294 20161
rect 15974 20096 15982 20160
rect 16046 20096 16062 20160
rect 16126 20096 16142 20160
rect 16206 20096 16222 20160
rect 16286 20096 16294 20160
rect 15974 20095 16294 20096
rect 22066 20000 22546 20120
rect 1577 19818 1643 19821
rect 62 19816 1643 19818
rect 62 19760 1582 19816
rect 1638 19760 1643 19816
rect 62 19758 1643 19760
rect 1577 19755 1643 19758
rect 18965 19818 19031 19821
rect 22142 19818 22202 20000
rect 18965 19816 22202 19818
rect 18965 19760 18970 19816
rect 19026 19760 22202 19816
rect 18965 19758 22202 19760
rect 18965 19755 19031 19758
rect 4701 19616 5021 19617
rect 4701 19552 4709 19616
rect 4773 19552 4789 19616
rect 4853 19552 4869 19616
rect 4933 19552 4949 19616
rect 5013 19552 5021 19616
rect 4701 19551 5021 19552
rect 12217 19616 12537 19617
rect 12217 19552 12225 19616
rect 12289 19552 12305 19616
rect 12369 19552 12385 19616
rect 12449 19552 12465 19616
rect 12529 19552 12537 19616
rect 12217 19551 12537 19552
rect 19732 19616 20052 19617
rect 19732 19552 19740 19616
rect 19804 19552 19820 19616
rect 19884 19552 19900 19616
rect 19964 19552 19980 19616
rect 20044 19552 20052 19616
rect 19732 19551 20052 19552
rect 7373 19274 7439 19277
rect 19609 19274 19675 19277
rect 20161 19274 20227 19277
rect 7373 19272 20227 19274
rect 7373 19216 7378 19272
rect 7434 19216 19614 19272
rect 19670 19216 20166 19272
rect 20222 19216 20227 19272
rect 7373 19214 20227 19216
rect 7373 19211 7439 19214
rect 19609 19211 19675 19214
rect 20161 19211 20227 19214
rect 0 19136 480 19168
rect 0 19080 110 19136
rect 166 19080 480 19136
rect 0 19048 480 19080
rect 8459 19072 8779 19073
rect 8459 19008 8467 19072
rect 8531 19008 8547 19072
rect 8611 19008 8627 19072
rect 8691 19008 8707 19072
rect 8771 19008 8779 19072
rect 8459 19007 8779 19008
rect 15974 19072 16294 19073
rect 15974 19008 15982 19072
rect 16046 19008 16062 19072
rect 16126 19008 16142 19072
rect 16206 19008 16222 19072
rect 16286 19008 16294 19072
rect 15974 19007 16294 19008
rect 22066 19002 22546 19032
rect 22012 19000 22546 19002
rect 22012 18944 22098 19000
rect 22154 18944 22546 19000
rect 22012 18942 22546 18944
rect 22066 18912 22546 18942
rect 4701 18528 5021 18529
rect 4701 18464 4709 18528
rect 4773 18464 4789 18528
rect 4853 18464 4869 18528
rect 4933 18464 4949 18528
rect 5013 18464 5021 18528
rect 4701 18463 5021 18464
rect 12217 18528 12537 18529
rect 12217 18464 12225 18528
rect 12289 18464 12305 18528
rect 12369 18464 12385 18528
rect 12449 18464 12465 18528
rect 12529 18464 12537 18528
rect 12217 18463 12537 18464
rect 19732 18528 20052 18529
rect 19732 18464 19740 18528
rect 19804 18464 19820 18528
rect 19884 18464 19900 18528
rect 19964 18464 19980 18528
rect 20044 18464 20052 18528
rect 19732 18463 20052 18464
rect 8459 17984 8779 17985
rect 0 17824 480 17944
rect 8459 17920 8467 17984
rect 8531 17920 8547 17984
rect 8611 17920 8627 17984
rect 8691 17920 8707 17984
rect 8771 17920 8779 17984
rect 8459 17919 8779 17920
rect 15974 17984 16294 17985
rect 15974 17920 15982 17984
rect 16046 17920 16062 17984
rect 16126 17920 16142 17984
rect 16206 17920 16222 17984
rect 16286 17920 16294 17984
rect 15974 17919 16294 17920
rect 22066 17824 22546 17944
rect 62 17370 122 17824
rect 19425 17642 19491 17645
rect 22142 17642 22202 17824
rect 19425 17640 22202 17642
rect 19425 17584 19430 17640
rect 19486 17584 22202 17640
rect 19425 17582 22202 17584
rect 19425 17579 19491 17582
rect 4701 17440 5021 17441
rect 4701 17376 4709 17440
rect 4773 17376 4789 17440
rect 4853 17376 4869 17440
rect 4933 17376 4949 17440
rect 5013 17376 5021 17440
rect 4701 17375 5021 17376
rect 12217 17440 12537 17441
rect 12217 17376 12225 17440
rect 12289 17376 12305 17440
rect 12369 17376 12385 17440
rect 12449 17376 12465 17440
rect 12529 17376 12537 17440
rect 12217 17375 12537 17376
rect 19732 17440 20052 17441
rect 19732 17376 19740 17440
rect 19804 17376 19820 17440
rect 19884 17376 19900 17440
rect 19964 17376 19980 17440
rect 20044 17376 20052 17440
rect 19732 17375 20052 17376
rect 2773 17370 2839 17373
rect 62 17368 2839 17370
rect 62 17312 2778 17368
rect 2834 17312 2839 17368
rect 62 17310 2839 17312
rect 2773 17307 2839 17310
rect 22093 17234 22159 17237
rect 19290 17232 22159 17234
rect 19290 17176 22098 17232
rect 22154 17176 22159 17232
rect 19290 17174 22159 17176
rect 8385 17098 8451 17101
rect 19290 17098 19350 17174
rect 22093 17171 22159 17174
rect 8385 17096 19350 17098
rect 8385 17040 8390 17096
rect 8446 17040 19350 17096
rect 8385 17038 19350 17040
rect 8385 17035 8451 17038
rect 8459 16896 8779 16897
rect 8459 16832 8467 16896
rect 8531 16832 8547 16896
rect 8611 16832 8627 16896
rect 8691 16832 8707 16896
rect 8771 16832 8779 16896
rect 8459 16831 8779 16832
rect 15974 16896 16294 16897
rect 15974 16832 15982 16896
rect 16046 16832 16062 16896
rect 16126 16832 16142 16896
rect 16206 16832 16222 16896
rect 16286 16832 16294 16896
rect 22066 16872 22546 16992
rect 15974 16831 16294 16832
rect 0 16600 480 16720
rect 62 16146 122 16600
rect 15469 16554 15535 16557
rect 22142 16554 22202 16872
rect 15469 16552 22202 16554
rect 15469 16496 15474 16552
rect 15530 16496 22202 16552
rect 15469 16494 22202 16496
rect 15469 16491 15535 16494
rect 4701 16352 5021 16353
rect 4701 16288 4709 16352
rect 4773 16288 4789 16352
rect 4853 16288 4869 16352
rect 4933 16288 4949 16352
rect 5013 16288 5021 16352
rect 4701 16287 5021 16288
rect 12217 16352 12537 16353
rect 12217 16288 12225 16352
rect 12289 16288 12305 16352
rect 12369 16288 12385 16352
rect 12449 16288 12465 16352
rect 12529 16288 12537 16352
rect 12217 16287 12537 16288
rect 19732 16352 20052 16353
rect 19732 16288 19740 16352
rect 19804 16288 19820 16352
rect 19884 16288 19900 16352
rect 19964 16288 19980 16352
rect 20044 16288 20052 16352
rect 19732 16287 20052 16288
rect 9305 16146 9371 16149
rect 62 16144 9371 16146
rect 62 16088 9310 16144
rect 9366 16088 9371 16144
rect 62 16086 9371 16088
rect 9305 16083 9371 16086
rect 8459 15808 8779 15809
rect 8459 15744 8467 15808
rect 8531 15744 8547 15808
rect 8611 15744 8627 15808
rect 8691 15744 8707 15808
rect 8771 15744 8779 15808
rect 8459 15743 8779 15744
rect 15974 15808 16294 15809
rect 15974 15744 15982 15808
rect 16046 15744 16062 15808
rect 16126 15744 16142 15808
rect 16206 15744 16222 15808
rect 16286 15744 16294 15808
rect 22066 15784 22546 15904
rect 15974 15743 16294 15744
rect 0 15376 480 15496
rect 17493 15466 17559 15469
rect 22142 15466 22202 15784
rect 17493 15464 22202 15466
rect 17493 15408 17498 15464
rect 17554 15408 22202 15464
rect 17493 15406 22202 15408
rect 17493 15403 17559 15406
rect 62 15058 122 15376
rect 4701 15264 5021 15265
rect 4701 15200 4709 15264
rect 4773 15200 4789 15264
rect 4853 15200 4869 15264
rect 4933 15200 4949 15264
rect 5013 15200 5021 15264
rect 4701 15199 5021 15200
rect 12217 15264 12537 15265
rect 12217 15200 12225 15264
rect 12289 15200 12305 15264
rect 12369 15200 12385 15264
rect 12449 15200 12465 15264
rect 12529 15200 12537 15264
rect 12217 15199 12537 15200
rect 19732 15264 20052 15265
rect 19732 15200 19740 15264
rect 19804 15200 19820 15264
rect 19884 15200 19900 15264
rect 19964 15200 19980 15264
rect 20044 15200 20052 15264
rect 19732 15199 20052 15200
rect 4613 15058 4679 15061
rect 62 15056 4679 15058
rect 62 15000 4618 15056
rect 4674 15000 4679 15056
rect 62 14998 4679 15000
rect 4613 14995 4679 14998
rect 7373 14922 7439 14925
rect 22066 14922 22546 14952
rect 7373 14920 22546 14922
rect 7373 14864 7378 14920
rect 7434 14864 22546 14920
rect 7373 14862 22546 14864
rect 7373 14859 7439 14862
rect 22066 14832 22546 14862
rect 8459 14720 8779 14721
rect 8459 14656 8467 14720
rect 8531 14656 8547 14720
rect 8611 14656 8627 14720
rect 8691 14656 8707 14720
rect 8771 14656 8779 14720
rect 8459 14655 8779 14656
rect 15974 14720 16294 14721
rect 15974 14656 15982 14720
rect 16046 14656 16062 14720
rect 16126 14656 16142 14720
rect 16206 14656 16222 14720
rect 16286 14656 16294 14720
rect 15974 14655 16294 14656
rect 0 14152 480 14272
rect 4701 14176 5021 14177
rect 62 13698 122 14152
rect 4701 14112 4709 14176
rect 4773 14112 4789 14176
rect 4853 14112 4869 14176
rect 4933 14112 4949 14176
rect 5013 14112 5021 14176
rect 4701 14111 5021 14112
rect 12217 14176 12537 14177
rect 12217 14112 12225 14176
rect 12289 14112 12305 14176
rect 12369 14112 12385 14176
rect 12449 14112 12465 14176
rect 12529 14112 12537 14176
rect 12217 14111 12537 14112
rect 19732 14176 20052 14177
rect 19732 14112 19740 14176
rect 19804 14112 19820 14176
rect 19884 14112 19900 14176
rect 19964 14112 19980 14176
rect 20044 14112 20052 14176
rect 19732 14111 20052 14112
rect 22066 13834 22546 13864
rect 22012 13832 22546 13834
rect 22012 13776 22098 13832
rect 22154 13776 22546 13832
rect 22012 13774 22546 13776
rect 22066 13744 22546 13774
rect 4245 13698 4311 13701
rect 62 13696 4311 13698
rect 62 13640 4250 13696
rect 4306 13640 4311 13696
rect 62 13638 4311 13640
rect 4245 13635 4311 13638
rect 8459 13632 8779 13633
rect 8459 13568 8467 13632
rect 8531 13568 8547 13632
rect 8611 13568 8627 13632
rect 8691 13568 8707 13632
rect 8771 13568 8779 13632
rect 8459 13567 8779 13568
rect 15974 13632 16294 13633
rect 15974 13568 15982 13632
rect 16046 13568 16062 13632
rect 16126 13568 16142 13632
rect 16206 13568 16222 13632
rect 16286 13568 16294 13632
rect 15974 13567 16294 13568
rect 21081 13154 21147 13157
rect 22134 13154 22140 13156
rect 21081 13152 22140 13154
rect 21081 13096 21086 13152
rect 21142 13096 22140 13152
rect 21081 13094 22140 13096
rect 21081 13091 21147 13094
rect 22134 13092 22140 13094
rect 22204 13092 22210 13156
rect 4701 13088 5021 13089
rect 0 13016 480 13048
rect 4701 13024 4709 13088
rect 4773 13024 4789 13088
rect 4853 13024 4869 13088
rect 4933 13024 4949 13088
rect 5013 13024 5021 13088
rect 4701 13023 5021 13024
rect 12217 13088 12537 13089
rect 12217 13024 12225 13088
rect 12289 13024 12305 13088
rect 12369 13024 12385 13088
rect 12449 13024 12465 13088
rect 12529 13024 12537 13088
rect 12217 13023 12537 13024
rect 19732 13088 20052 13089
rect 19732 13024 19740 13088
rect 19804 13024 19820 13088
rect 19884 13024 19900 13088
rect 19964 13024 19980 13088
rect 20044 13024 20052 13088
rect 19732 13023 20052 13024
rect 0 12960 110 13016
rect 166 12960 480 13016
rect 0 12928 480 12960
rect 22066 12884 22546 12912
rect 22066 12882 22140 12884
rect 22012 12822 22140 12882
rect 22066 12820 22140 12822
rect 22204 12820 22546 12884
rect 22066 12792 22546 12820
rect 8459 12544 8779 12545
rect 8459 12480 8467 12544
rect 8531 12480 8547 12544
rect 8611 12480 8627 12544
rect 8691 12480 8707 12544
rect 8771 12480 8779 12544
rect 8459 12479 8779 12480
rect 15974 12544 16294 12545
rect 15974 12480 15982 12544
rect 16046 12480 16062 12544
rect 16126 12480 16142 12544
rect 16206 12480 16222 12544
rect 16286 12480 16294 12544
rect 15974 12479 16294 12480
rect 4701 12000 5021 12001
rect 4701 11936 4709 12000
rect 4773 11936 4789 12000
rect 4853 11936 4869 12000
rect 4933 11936 4949 12000
rect 5013 11936 5021 12000
rect 4701 11935 5021 11936
rect 12217 12000 12537 12001
rect 12217 11936 12225 12000
rect 12289 11936 12305 12000
rect 12369 11936 12385 12000
rect 12449 11936 12465 12000
rect 12529 11936 12537 12000
rect 12217 11935 12537 11936
rect 19732 12000 20052 12001
rect 19732 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20052 12000
rect 19732 11935 20052 11936
rect 54 11868 60 11932
rect 124 11930 130 11932
rect 2497 11930 2563 11933
rect 124 11928 2563 11930
rect 124 11872 2502 11928
rect 2558 11872 2563 11928
rect 124 11870 2563 11872
rect 124 11868 130 11870
rect 2497 11867 2563 11870
rect 22066 11704 22546 11824
rect 0 11660 480 11688
rect 0 11596 60 11660
rect 124 11596 480 11660
rect 0 11568 480 11596
rect 8459 11456 8779 11457
rect 8459 11392 8467 11456
rect 8531 11392 8547 11456
rect 8611 11392 8627 11456
rect 8691 11392 8707 11456
rect 8771 11392 8779 11456
rect 8459 11391 8779 11392
rect 15974 11456 16294 11457
rect 15974 11392 15982 11456
rect 16046 11392 16062 11456
rect 16126 11392 16142 11456
rect 16206 11392 16222 11456
rect 16286 11392 16294 11456
rect 15974 11391 16294 11392
rect 20161 11250 20227 11253
rect 22142 11250 22202 11704
rect 20161 11248 22202 11250
rect 20161 11192 20166 11248
rect 20222 11192 22202 11248
rect 20161 11190 22202 11192
rect 20161 11187 20227 11190
rect 4701 10912 5021 10913
rect 4701 10848 4709 10912
rect 4773 10848 4789 10912
rect 4853 10848 4869 10912
rect 4933 10848 4949 10912
rect 5013 10848 5021 10912
rect 4701 10847 5021 10848
rect 12217 10912 12537 10913
rect 12217 10848 12225 10912
rect 12289 10848 12305 10912
rect 12369 10848 12385 10912
rect 12449 10848 12465 10912
rect 12529 10848 12537 10912
rect 12217 10847 12537 10848
rect 19732 10912 20052 10913
rect 19732 10848 19740 10912
rect 19804 10848 19820 10912
rect 19884 10848 19900 10912
rect 19964 10848 19980 10912
rect 20044 10848 20052 10912
rect 19732 10847 20052 10848
rect 22066 10708 22546 10736
rect 22066 10706 22140 10708
rect 22012 10646 22140 10706
rect 22066 10644 22140 10646
rect 22204 10644 22546 10708
rect 22066 10616 22546 10644
rect 3877 10570 3943 10573
rect 9949 10570 10015 10573
rect 3877 10568 10015 10570
rect 3877 10512 3882 10568
rect 3938 10512 9954 10568
rect 10010 10512 10015 10568
rect 3877 10510 10015 10512
rect 3877 10507 3943 10510
rect 9949 10507 10015 10510
rect 14273 10570 14339 10573
rect 14273 10568 19350 10570
rect 14273 10512 14278 10568
rect 14334 10512 19350 10568
rect 14273 10510 19350 10512
rect 14273 10507 14339 10510
rect 0 10344 480 10464
rect 19290 10434 19350 10510
rect 22134 10434 22140 10436
rect 19290 10374 22140 10434
rect 22134 10372 22140 10374
rect 22204 10372 22210 10436
rect 8459 10368 8779 10369
rect 62 9890 122 10344
rect 8459 10304 8467 10368
rect 8531 10304 8547 10368
rect 8611 10304 8627 10368
rect 8691 10304 8707 10368
rect 8771 10304 8779 10368
rect 8459 10303 8779 10304
rect 15974 10368 16294 10369
rect 15974 10304 15982 10368
rect 16046 10304 16062 10368
rect 16126 10304 16142 10368
rect 16206 10304 16222 10368
rect 16286 10304 16294 10368
rect 15974 10303 16294 10304
rect 1393 9890 1459 9893
rect 62 9888 1459 9890
rect 62 9832 1398 9888
rect 1454 9832 1459 9888
rect 62 9830 1459 9832
rect 1393 9827 1459 9830
rect 4701 9824 5021 9825
rect 4701 9760 4709 9824
rect 4773 9760 4789 9824
rect 4853 9760 4869 9824
rect 4933 9760 4949 9824
rect 5013 9760 5021 9824
rect 4701 9759 5021 9760
rect 12217 9824 12537 9825
rect 12217 9760 12225 9824
rect 12289 9760 12305 9824
rect 12369 9760 12385 9824
rect 12449 9760 12465 9824
rect 12529 9760 12537 9824
rect 12217 9759 12537 9760
rect 19732 9824 20052 9825
rect 19732 9760 19740 9824
rect 19804 9760 19820 9824
rect 19884 9760 19900 9824
rect 19964 9760 19980 9824
rect 20044 9760 20052 9824
rect 19732 9759 20052 9760
rect 22066 9664 22546 9784
rect 5717 9482 5783 9485
rect 13353 9482 13419 9485
rect 14641 9482 14707 9485
rect 5717 9480 14707 9482
rect 5717 9424 5722 9480
rect 5778 9424 13358 9480
rect 13414 9424 14646 9480
rect 14702 9424 14707 9480
rect 5717 9422 14707 9424
rect 5717 9419 5783 9422
rect 13353 9419 13419 9422
rect 14641 9419 14707 9422
rect 20161 9346 20227 9349
rect 22142 9346 22202 9664
rect 20161 9344 22202 9346
rect 20161 9288 20166 9344
rect 20222 9288 22202 9344
rect 20161 9286 22202 9288
rect 20161 9283 20227 9286
rect 8459 9280 8779 9281
rect 0 9120 480 9240
rect 8459 9216 8467 9280
rect 8531 9216 8547 9280
rect 8611 9216 8627 9280
rect 8691 9216 8707 9280
rect 8771 9216 8779 9280
rect 8459 9215 8779 9216
rect 15974 9280 16294 9281
rect 15974 9216 15982 9280
rect 16046 9216 16062 9280
rect 16126 9216 16142 9280
rect 16206 9216 16222 9280
rect 16286 9216 16294 9280
rect 15974 9215 16294 9216
rect 62 8666 122 9120
rect 4701 8736 5021 8737
rect 4701 8672 4709 8736
rect 4773 8672 4789 8736
rect 4853 8672 4869 8736
rect 4933 8672 4949 8736
rect 5013 8672 5021 8736
rect 4701 8671 5021 8672
rect 12217 8736 12537 8737
rect 12217 8672 12225 8736
rect 12289 8672 12305 8736
rect 12369 8672 12385 8736
rect 12449 8672 12465 8736
rect 12529 8672 12537 8736
rect 12217 8671 12537 8672
rect 19732 8736 20052 8737
rect 19732 8672 19740 8736
rect 19804 8672 19820 8736
rect 19884 8672 19900 8736
rect 19964 8672 19980 8736
rect 20044 8672 20052 8736
rect 19732 8671 20052 8672
rect 2589 8666 2655 8669
rect 62 8664 2655 8666
rect 62 8608 2594 8664
rect 2650 8608 2655 8664
rect 62 8606 2655 8608
rect 2589 8603 2655 8606
rect 20161 8666 20227 8669
rect 22066 8666 22546 8696
rect 20161 8664 22546 8666
rect 20161 8608 20166 8664
rect 20222 8608 22546 8664
rect 20161 8606 22546 8608
rect 20161 8603 20227 8606
rect 22066 8576 22546 8606
rect 8459 8192 8779 8193
rect 8459 8128 8467 8192
rect 8531 8128 8547 8192
rect 8611 8128 8627 8192
rect 8691 8128 8707 8192
rect 8771 8128 8779 8192
rect 8459 8127 8779 8128
rect 15974 8192 16294 8193
rect 15974 8128 15982 8192
rect 16046 8128 16062 8192
rect 16126 8128 16142 8192
rect 16206 8128 16222 8192
rect 16286 8128 16294 8192
rect 15974 8127 16294 8128
rect 0 7896 480 8016
rect 5349 7986 5415 7989
rect 18597 7986 18663 7989
rect 5349 7984 18663 7986
rect 5349 7928 5354 7984
rect 5410 7928 18602 7984
rect 18658 7928 18663 7984
rect 5349 7926 18663 7928
rect 5349 7923 5415 7926
rect 18597 7923 18663 7926
rect 62 7442 122 7896
rect 4701 7648 5021 7649
rect 4701 7584 4709 7648
rect 4773 7584 4789 7648
rect 4853 7584 4869 7648
rect 4933 7584 4949 7648
rect 5013 7584 5021 7648
rect 4701 7583 5021 7584
rect 12217 7648 12537 7649
rect 12217 7584 12225 7648
rect 12289 7584 12305 7648
rect 12369 7584 12385 7648
rect 12449 7584 12465 7648
rect 12529 7584 12537 7648
rect 12217 7583 12537 7584
rect 19732 7648 20052 7649
rect 19732 7584 19740 7648
rect 19804 7584 19820 7648
rect 19884 7584 19900 7648
rect 19964 7584 19980 7648
rect 20044 7584 20052 7648
rect 22066 7624 22546 7744
rect 19732 7583 20052 7584
rect 5165 7442 5231 7445
rect 62 7440 5231 7442
rect 62 7384 5170 7440
rect 5226 7384 5231 7440
rect 62 7382 5231 7384
rect 5165 7379 5231 7382
rect 2681 7306 2747 7309
rect 62 7304 2747 7306
rect 62 7248 2686 7304
rect 2742 7248 2747 7304
rect 62 7246 2747 7248
rect 62 6792 122 7246
rect 2681 7243 2747 7246
rect 10961 7306 11027 7309
rect 22142 7306 22202 7624
rect 10961 7304 22202 7306
rect 10961 7248 10966 7304
rect 11022 7248 22202 7304
rect 10961 7246 22202 7248
rect 10961 7243 11027 7246
rect 8459 7104 8779 7105
rect 8459 7040 8467 7104
rect 8531 7040 8547 7104
rect 8611 7040 8627 7104
rect 8691 7040 8707 7104
rect 8771 7040 8779 7104
rect 8459 7039 8779 7040
rect 15974 7104 16294 7105
rect 15974 7040 15982 7104
rect 16046 7040 16062 7104
rect 16126 7040 16142 7104
rect 16206 7040 16222 7104
rect 16286 7040 16294 7104
rect 15974 7039 16294 7040
rect 0 6672 480 6792
rect 4701 6560 5021 6561
rect 4701 6496 4709 6560
rect 4773 6496 4789 6560
rect 4853 6496 4869 6560
rect 4933 6496 4949 6560
rect 5013 6496 5021 6560
rect 4701 6495 5021 6496
rect 12217 6560 12537 6561
rect 12217 6496 12225 6560
rect 12289 6496 12305 6560
rect 12369 6496 12385 6560
rect 12449 6496 12465 6560
rect 12529 6496 12537 6560
rect 12217 6495 12537 6496
rect 19732 6560 20052 6561
rect 19732 6496 19740 6560
rect 19804 6496 19820 6560
rect 19884 6496 19900 6560
rect 19964 6496 19980 6560
rect 20044 6496 20052 6560
rect 22066 6536 22546 6656
rect 19732 6495 20052 6496
rect 16941 6354 17007 6357
rect 22142 6354 22202 6536
rect 16941 6352 22202 6354
rect 16941 6296 16946 6352
rect 17002 6296 22202 6352
rect 16941 6294 22202 6296
rect 16941 6291 17007 6294
rect 8459 6016 8779 6017
rect 8459 5952 8467 6016
rect 8531 5952 8547 6016
rect 8611 5952 8627 6016
rect 8691 5952 8707 6016
rect 8771 5952 8779 6016
rect 8459 5951 8779 5952
rect 15974 6016 16294 6017
rect 15974 5952 15982 6016
rect 16046 5952 16062 6016
rect 16126 5952 16142 6016
rect 16206 5952 16222 6016
rect 16286 5952 16294 6016
rect 15974 5951 16294 5952
rect 0 5536 480 5568
rect 0 5480 110 5536
rect 166 5480 480 5536
rect 0 5448 480 5480
rect 20161 5538 20227 5541
rect 22066 5538 22546 5568
rect 20161 5536 22546 5538
rect 20161 5480 20166 5536
rect 20222 5480 22546 5536
rect 20161 5478 22546 5480
rect 20161 5475 20227 5478
rect 4701 5472 5021 5473
rect 4701 5408 4709 5472
rect 4773 5408 4789 5472
rect 4853 5408 4869 5472
rect 4933 5408 4949 5472
rect 5013 5408 5021 5472
rect 4701 5407 5021 5408
rect 12217 5472 12537 5473
rect 12217 5408 12225 5472
rect 12289 5408 12305 5472
rect 12369 5408 12385 5472
rect 12449 5408 12465 5472
rect 12529 5408 12537 5472
rect 12217 5407 12537 5408
rect 19732 5472 20052 5473
rect 19732 5408 19740 5472
rect 19804 5408 19820 5472
rect 19884 5408 19900 5472
rect 19964 5408 19980 5472
rect 20044 5408 20052 5472
rect 22066 5448 22546 5478
rect 19732 5407 20052 5408
rect 6453 5266 6519 5269
rect 16297 5266 16363 5269
rect 6453 5264 16363 5266
rect 6453 5208 6458 5264
rect 6514 5208 16302 5264
rect 16358 5208 16363 5264
rect 6453 5206 16363 5208
rect 6453 5203 6519 5206
rect 16297 5203 16363 5206
rect 20253 5130 20319 5133
rect 20253 5128 22202 5130
rect 20253 5072 20258 5128
rect 20314 5072 22202 5128
rect 20253 5070 22202 5072
rect 20253 5067 20319 5070
rect 8459 4928 8779 4929
rect 8459 4864 8467 4928
rect 8531 4864 8547 4928
rect 8611 4864 8627 4928
rect 8691 4864 8707 4928
rect 8771 4864 8779 4928
rect 8459 4863 8779 4864
rect 15974 4928 16294 4929
rect 15974 4864 15982 4928
rect 16046 4864 16062 4928
rect 16126 4864 16142 4928
rect 16206 4864 16222 4928
rect 16286 4864 16294 4928
rect 15974 4863 16294 4864
rect 22142 4616 22202 5070
rect 22066 4496 22546 4616
rect 4701 4384 5021 4385
rect 0 4224 480 4344
rect 4701 4320 4709 4384
rect 4773 4320 4789 4384
rect 4853 4320 4869 4384
rect 4933 4320 4949 4384
rect 5013 4320 5021 4384
rect 4701 4319 5021 4320
rect 12217 4384 12537 4385
rect 12217 4320 12225 4384
rect 12289 4320 12305 4384
rect 12369 4320 12385 4384
rect 12449 4320 12465 4384
rect 12529 4320 12537 4384
rect 12217 4319 12537 4320
rect 19732 4384 20052 4385
rect 19732 4320 19740 4384
rect 19804 4320 19820 4384
rect 19884 4320 19900 4384
rect 19964 4320 19980 4384
rect 20044 4320 20052 4384
rect 19732 4319 20052 4320
rect 62 4042 122 4224
rect 8293 4178 8359 4181
rect 8293 4176 8586 4178
rect 8293 4120 8298 4176
rect 8354 4120 8586 4176
rect 8293 4118 8586 4120
rect 8293 4115 8359 4118
rect 8385 4042 8451 4045
rect 62 4040 8451 4042
rect 62 3984 8390 4040
rect 8446 3984 8451 4040
rect 62 3982 8451 3984
rect 8526 4042 8586 4118
rect 20069 4042 20135 4045
rect 8526 4040 20135 4042
rect 8526 3984 20074 4040
rect 20130 3984 20135 4040
rect 8526 3982 20135 3984
rect 8385 3979 8451 3982
rect 20069 3979 20135 3982
rect 8459 3840 8779 3841
rect 8459 3776 8467 3840
rect 8531 3776 8547 3840
rect 8611 3776 8627 3840
rect 8691 3776 8707 3840
rect 8771 3776 8779 3840
rect 8459 3775 8779 3776
rect 15974 3840 16294 3841
rect 15974 3776 15982 3840
rect 16046 3776 16062 3840
rect 16126 3776 16142 3840
rect 16206 3776 16222 3840
rect 16286 3776 16294 3840
rect 15974 3775 16294 3776
rect 11973 3634 12039 3637
rect 62 3632 12039 3634
rect 62 3576 11978 3632
rect 12034 3576 12039 3632
rect 62 3574 12039 3576
rect 62 3120 122 3574
rect 11973 3571 12039 3574
rect 22066 3408 22546 3528
rect 4701 3296 5021 3297
rect 4701 3232 4709 3296
rect 4773 3232 4789 3296
rect 4853 3232 4869 3296
rect 4933 3232 4949 3296
rect 5013 3232 5021 3296
rect 4701 3231 5021 3232
rect 12217 3296 12537 3297
rect 12217 3232 12225 3296
rect 12289 3232 12305 3296
rect 12369 3232 12385 3296
rect 12449 3232 12465 3296
rect 12529 3232 12537 3296
rect 12217 3231 12537 3232
rect 19732 3296 20052 3297
rect 19732 3232 19740 3296
rect 19804 3232 19820 3296
rect 19884 3232 19900 3296
rect 19964 3232 19980 3296
rect 20044 3232 20052 3296
rect 19732 3231 20052 3232
rect 0 3000 480 3120
rect 8459 2752 8779 2753
rect 8459 2688 8467 2752
rect 8531 2688 8547 2752
rect 8611 2688 8627 2752
rect 8691 2688 8707 2752
rect 8771 2688 8779 2752
rect 8459 2687 8779 2688
rect 15974 2752 16294 2753
rect 15974 2688 15982 2752
rect 16046 2688 16062 2752
rect 16126 2688 16142 2752
rect 16206 2688 16222 2752
rect 16286 2688 16294 2752
rect 15974 2687 16294 2688
rect 22066 2456 22546 2576
rect 1301 2410 1367 2413
rect 62 2408 1367 2410
rect 62 2352 1306 2408
rect 1362 2352 1367 2408
rect 62 2350 1367 2352
rect 62 1896 122 2350
rect 1301 2347 1367 2350
rect 4701 2208 5021 2209
rect 4701 2144 4709 2208
rect 4773 2144 4789 2208
rect 4853 2144 4869 2208
rect 4933 2144 4949 2208
rect 5013 2144 5021 2208
rect 4701 2143 5021 2144
rect 12217 2208 12537 2209
rect 12217 2144 12225 2208
rect 12289 2144 12305 2208
rect 12369 2144 12385 2208
rect 12449 2144 12465 2208
rect 12529 2144 12537 2208
rect 12217 2143 12537 2144
rect 19732 2208 20052 2209
rect 19732 2144 19740 2208
rect 19804 2144 19820 2208
rect 19884 2144 19900 2208
rect 19964 2144 19980 2208
rect 20044 2144 20052 2208
rect 19732 2143 20052 2144
rect 0 1776 480 1896
rect 2221 1458 2287 1461
rect 11329 1458 11395 1461
rect 2221 1456 11395 1458
rect 2221 1400 2226 1456
rect 2282 1400 11334 1456
rect 11390 1400 11395 1456
rect 2221 1398 11395 1400
rect 2221 1395 2287 1398
rect 11329 1395 11395 1398
rect 22066 1368 22546 1488
rect 0 552 480 672
rect 22066 416 22546 536
<< via3 >>
rect 8467 22332 8531 22336
rect 8467 22276 8471 22332
rect 8471 22276 8527 22332
rect 8527 22276 8531 22332
rect 8467 22272 8531 22276
rect 8547 22332 8611 22336
rect 8547 22276 8551 22332
rect 8551 22276 8607 22332
rect 8607 22276 8611 22332
rect 8547 22272 8611 22276
rect 8627 22332 8691 22336
rect 8627 22276 8631 22332
rect 8631 22276 8687 22332
rect 8687 22276 8691 22332
rect 8627 22272 8691 22276
rect 8707 22332 8771 22336
rect 8707 22276 8711 22332
rect 8711 22276 8767 22332
rect 8767 22276 8771 22332
rect 8707 22272 8771 22276
rect 15982 22332 16046 22336
rect 15982 22276 15986 22332
rect 15986 22276 16042 22332
rect 16042 22276 16046 22332
rect 15982 22272 16046 22276
rect 16062 22332 16126 22336
rect 16062 22276 16066 22332
rect 16066 22276 16122 22332
rect 16122 22276 16126 22332
rect 16062 22272 16126 22276
rect 16142 22332 16206 22336
rect 16142 22276 16146 22332
rect 16146 22276 16202 22332
rect 16202 22276 16206 22332
rect 16142 22272 16206 22276
rect 16222 22332 16286 22336
rect 16222 22276 16226 22332
rect 16226 22276 16282 22332
rect 16282 22276 16286 22332
rect 16222 22272 16286 22276
rect 4709 21788 4773 21792
rect 4709 21732 4713 21788
rect 4713 21732 4769 21788
rect 4769 21732 4773 21788
rect 4709 21728 4773 21732
rect 4789 21788 4853 21792
rect 4789 21732 4793 21788
rect 4793 21732 4849 21788
rect 4849 21732 4853 21788
rect 4789 21728 4853 21732
rect 4869 21788 4933 21792
rect 4869 21732 4873 21788
rect 4873 21732 4929 21788
rect 4929 21732 4933 21788
rect 4869 21728 4933 21732
rect 4949 21788 5013 21792
rect 4949 21732 4953 21788
rect 4953 21732 5009 21788
rect 5009 21732 5013 21788
rect 4949 21728 5013 21732
rect 12225 21788 12289 21792
rect 12225 21732 12229 21788
rect 12229 21732 12285 21788
rect 12285 21732 12289 21788
rect 12225 21728 12289 21732
rect 12305 21788 12369 21792
rect 12305 21732 12309 21788
rect 12309 21732 12365 21788
rect 12365 21732 12369 21788
rect 12305 21728 12369 21732
rect 12385 21788 12449 21792
rect 12385 21732 12389 21788
rect 12389 21732 12445 21788
rect 12445 21732 12449 21788
rect 12385 21728 12449 21732
rect 12465 21788 12529 21792
rect 12465 21732 12469 21788
rect 12469 21732 12525 21788
rect 12525 21732 12529 21788
rect 12465 21728 12529 21732
rect 19740 21788 19804 21792
rect 19740 21732 19744 21788
rect 19744 21732 19800 21788
rect 19800 21732 19804 21788
rect 19740 21728 19804 21732
rect 19820 21788 19884 21792
rect 19820 21732 19824 21788
rect 19824 21732 19880 21788
rect 19880 21732 19884 21788
rect 19820 21728 19884 21732
rect 19900 21788 19964 21792
rect 19900 21732 19904 21788
rect 19904 21732 19960 21788
rect 19960 21732 19964 21788
rect 19900 21728 19964 21732
rect 19980 21788 20044 21792
rect 19980 21732 19984 21788
rect 19984 21732 20040 21788
rect 20040 21732 20044 21788
rect 19980 21728 20044 21732
rect 8467 21244 8531 21248
rect 8467 21188 8471 21244
rect 8471 21188 8527 21244
rect 8527 21188 8531 21244
rect 8467 21184 8531 21188
rect 8547 21244 8611 21248
rect 8547 21188 8551 21244
rect 8551 21188 8607 21244
rect 8607 21188 8611 21244
rect 8547 21184 8611 21188
rect 8627 21244 8691 21248
rect 8627 21188 8631 21244
rect 8631 21188 8687 21244
rect 8687 21188 8691 21244
rect 8627 21184 8691 21188
rect 8707 21244 8771 21248
rect 8707 21188 8711 21244
rect 8711 21188 8767 21244
rect 8767 21188 8771 21244
rect 8707 21184 8771 21188
rect 15982 21244 16046 21248
rect 15982 21188 15986 21244
rect 15986 21188 16042 21244
rect 16042 21188 16046 21244
rect 15982 21184 16046 21188
rect 16062 21244 16126 21248
rect 16062 21188 16066 21244
rect 16066 21188 16122 21244
rect 16122 21188 16126 21244
rect 16062 21184 16126 21188
rect 16142 21244 16206 21248
rect 16142 21188 16146 21244
rect 16146 21188 16202 21244
rect 16202 21188 16206 21244
rect 16142 21184 16206 21188
rect 16222 21244 16286 21248
rect 16222 21188 16226 21244
rect 16226 21188 16282 21244
rect 16282 21188 16286 21244
rect 16222 21184 16286 21188
rect 4709 20700 4773 20704
rect 4709 20644 4713 20700
rect 4713 20644 4769 20700
rect 4769 20644 4773 20700
rect 4709 20640 4773 20644
rect 4789 20700 4853 20704
rect 4789 20644 4793 20700
rect 4793 20644 4849 20700
rect 4849 20644 4853 20700
rect 4789 20640 4853 20644
rect 4869 20700 4933 20704
rect 4869 20644 4873 20700
rect 4873 20644 4929 20700
rect 4929 20644 4933 20700
rect 4869 20640 4933 20644
rect 4949 20700 5013 20704
rect 4949 20644 4953 20700
rect 4953 20644 5009 20700
rect 5009 20644 5013 20700
rect 4949 20640 5013 20644
rect 12225 20700 12289 20704
rect 12225 20644 12229 20700
rect 12229 20644 12285 20700
rect 12285 20644 12289 20700
rect 12225 20640 12289 20644
rect 12305 20700 12369 20704
rect 12305 20644 12309 20700
rect 12309 20644 12365 20700
rect 12365 20644 12369 20700
rect 12305 20640 12369 20644
rect 12385 20700 12449 20704
rect 12385 20644 12389 20700
rect 12389 20644 12445 20700
rect 12445 20644 12449 20700
rect 12385 20640 12449 20644
rect 12465 20700 12529 20704
rect 12465 20644 12469 20700
rect 12469 20644 12525 20700
rect 12525 20644 12529 20700
rect 12465 20640 12529 20644
rect 19740 20700 19804 20704
rect 19740 20644 19744 20700
rect 19744 20644 19800 20700
rect 19800 20644 19804 20700
rect 19740 20640 19804 20644
rect 19820 20700 19884 20704
rect 19820 20644 19824 20700
rect 19824 20644 19880 20700
rect 19880 20644 19884 20700
rect 19820 20640 19884 20644
rect 19900 20700 19964 20704
rect 19900 20644 19904 20700
rect 19904 20644 19960 20700
rect 19960 20644 19964 20700
rect 19900 20640 19964 20644
rect 19980 20700 20044 20704
rect 19980 20644 19984 20700
rect 19984 20644 20040 20700
rect 20040 20644 20044 20700
rect 19980 20640 20044 20644
rect 8467 20156 8531 20160
rect 8467 20100 8471 20156
rect 8471 20100 8527 20156
rect 8527 20100 8531 20156
rect 8467 20096 8531 20100
rect 8547 20156 8611 20160
rect 8547 20100 8551 20156
rect 8551 20100 8607 20156
rect 8607 20100 8611 20156
rect 8547 20096 8611 20100
rect 8627 20156 8691 20160
rect 8627 20100 8631 20156
rect 8631 20100 8687 20156
rect 8687 20100 8691 20156
rect 8627 20096 8691 20100
rect 8707 20156 8771 20160
rect 8707 20100 8711 20156
rect 8711 20100 8767 20156
rect 8767 20100 8771 20156
rect 8707 20096 8771 20100
rect 15982 20156 16046 20160
rect 15982 20100 15986 20156
rect 15986 20100 16042 20156
rect 16042 20100 16046 20156
rect 15982 20096 16046 20100
rect 16062 20156 16126 20160
rect 16062 20100 16066 20156
rect 16066 20100 16122 20156
rect 16122 20100 16126 20156
rect 16062 20096 16126 20100
rect 16142 20156 16206 20160
rect 16142 20100 16146 20156
rect 16146 20100 16202 20156
rect 16202 20100 16206 20156
rect 16142 20096 16206 20100
rect 16222 20156 16286 20160
rect 16222 20100 16226 20156
rect 16226 20100 16282 20156
rect 16282 20100 16286 20156
rect 16222 20096 16286 20100
rect 4709 19612 4773 19616
rect 4709 19556 4713 19612
rect 4713 19556 4769 19612
rect 4769 19556 4773 19612
rect 4709 19552 4773 19556
rect 4789 19612 4853 19616
rect 4789 19556 4793 19612
rect 4793 19556 4849 19612
rect 4849 19556 4853 19612
rect 4789 19552 4853 19556
rect 4869 19612 4933 19616
rect 4869 19556 4873 19612
rect 4873 19556 4929 19612
rect 4929 19556 4933 19612
rect 4869 19552 4933 19556
rect 4949 19612 5013 19616
rect 4949 19556 4953 19612
rect 4953 19556 5009 19612
rect 5009 19556 5013 19612
rect 4949 19552 5013 19556
rect 12225 19612 12289 19616
rect 12225 19556 12229 19612
rect 12229 19556 12285 19612
rect 12285 19556 12289 19612
rect 12225 19552 12289 19556
rect 12305 19612 12369 19616
rect 12305 19556 12309 19612
rect 12309 19556 12365 19612
rect 12365 19556 12369 19612
rect 12305 19552 12369 19556
rect 12385 19612 12449 19616
rect 12385 19556 12389 19612
rect 12389 19556 12445 19612
rect 12445 19556 12449 19612
rect 12385 19552 12449 19556
rect 12465 19612 12529 19616
rect 12465 19556 12469 19612
rect 12469 19556 12525 19612
rect 12525 19556 12529 19612
rect 12465 19552 12529 19556
rect 19740 19612 19804 19616
rect 19740 19556 19744 19612
rect 19744 19556 19800 19612
rect 19800 19556 19804 19612
rect 19740 19552 19804 19556
rect 19820 19612 19884 19616
rect 19820 19556 19824 19612
rect 19824 19556 19880 19612
rect 19880 19556 19884 19612
rect 19820 19552 19884 19556
rect 19900 19612 19964 19616
rect 19900 19556 19904 19612
rect 19904 19556 19960 19612
rect 19960 19556 19964 19612
rect 19900 19552 19964 19556
rect 19980 19612 20044 19616
rect 19980 19556 19984 19612
rect 19984 19556 20040 19612
rect 20040 19556 20044 19612
rect 19980 19552 20044 19556
rect 8467 19068 8531 19072
rect 8467 19012 8471 19068
rect 8471 19012 8527 19068
rect 8527 19012 8531 19068
rect 8467 19008 8531 19012
rect 8547 19068 8611 19072
rect 8547 19012 8551 19068
rect 8551 19012 8607 19068
rect 8607 19012 8611 19068
rect 8547 19008 8611 19012
rect 8627 19068 8691 19072
rect 8627 19012 8631 19068
rect 8631 19012 8687 19068
rect 8687 19012 8691 19068
rect 8627 19008 8691 19012
rect 8707 19068 8771 19072
rect 8707 19012 8711 19068
rect 8711 19012 8767 19068
rect 8767 19012 8771 19068
rect 8707 19008 8771 19012
rect 15982 19068 16046 19072
rect 15982 19012 15986 19068
rect 15986 19012 16042 19068
rect 16042 19012 16046 19068
rect 15982 19008 16046 19012
rect 16062 19068 16126 19072
rect 16062 19012 16066 19068
rect 16066 19012 16122 19068
rect 16122 19012 16126 19068
rect 16062 19008 16126 19012
rect 16142 19068 16206 19072
rect 16142 19012 16146 19068
rect 16146 19012 16202 19068
rect 16202 19012 16206 19068
rect 16142 19008 16206 19012
rect 16222 19068 16286 19072
rect 16222 19012 16226 19068
rect 16226 19012 16282 19068
rect 16282 19012 16286 19068
rect 16222 19008 16286 19012
rect 4709 18524 4773 18528
rect 4709 18468 4713 18524
rect 4713 18468 4769 18524
rect 4769 18468 4773 18524
rect 4709 18464 4773 18468
rect 4789 18524 4853 18528
rect 4789 18468 4793 18524
rect 4793 18468 4849 18524
rect 4849 18468 4853 18524
rect 4789 18464 4853 18468
rect 4869 18524 4933 18528
rect 4869 18468 4873 18524
rect 4873 18468 4929 18524
rect 4929 18468 4933 18524
rect 4869 18464 4933 18468
rect 4949 18524 5013 18528
rect 4949 18468 4953 18524
rect 4953 18468 5009 18524
rect 5009 18468 5013 18524
rect 4949 18464 5013 18468
rect 12225 18524 12289 18528
rect 12225 18468 12229 18524
rect 12229 18468 12285 18524
rect 12285 18468 12289 18524
rect 12225 18464 12289 18468
rect 12305 18524 12369 18528
rect 12305 18468 12309 18524
rect 12309 18468 12365 18524
rect 12365 18468 12369 18524
rect 12305 18464 12369 18468
rect 12385 18524 12449 18528
rect 12385 18468 12389 18524
rect 12389 18468 12445 18524
rect 12445 18468 12449 18524
rect 12385 18464 12449 18468
rect 12465 18524 12529 18528
rect 12465 18468 12469 18524
rect 12469 18468 12525 18524
rect 12525 18468 12529 18524
rect 12465 18464 12529 18468
rect 19740 18524 19804 18528
rect 19740 18468 19744 18524
rect 19744 18468 19800 18524
rect 19800 18468 19804 18524
rect 19740 18464 19804 18468
rect 19820 18524 19884 18528
rect 19820 18468 19824 18524
rect 19824 18468 19880 18524
rect 19880 18468 19884 18524
rect 19820 18464 19884 18468
rect 19900 18524 19964 18528
rect 19900 18468 19904 18524
rect 19904 18468 19960 18524
rect 19960 18468 19964 18524
rect 19900 18464 19964 18468
rect 19980 18524 20044 18528
rect 19980 18468 19984 18524
rect 19984 18468 20040 18524
rect 20040 18468 20044 18524
rect 19980 18464 20044 18468
rect 8467 17980 8531 17984
rect 8467 17924 8471 17980
rect 8471 17924 8527 17980
rect 8527 17924 8531 17980
rect 8467 17920 8531 17924
rect 8547 17980 8611 17984
rect 8547 17924 8551 17980
rect 8551 17924 8607 17980
rect 8607 17924 8611 17980
rect 8547 17920 8611 17924
rect 8627 17980 8691 17984
rect 8627 17924 8631 17980
rect 8631 17924 8687 17980
rect 8687 17924 8691 17980
rect 8627 17920 8691 17924
rect 8707 17980 8771 17984
rect 8707 17924 8711 17980
rect 8711 17924 8767 17980
rect 8767 17924 8771 17980
rect 8707 17920 8771 17924
rect 15982 17980 16046 17984
rect 15982 17924 15986 17980
rect 15986 17924 16042 17980
rect 16042 17924 16046 17980
rect 15982 17920 16046 17924
rect 16062 17980 16126 17984
rect 16062 17924 16066 17980
rect 16066 17924 16122 17980
rect 16122 17924 16126 17980
rect 16062 17920 16126 17924
rect 16142 17980 16206 17984
rect 16142 17924 16146 17980
rect 16146 17924 16202 17980
rect 16202 17924 16206 17980
rect 16142 17920 16206 17924
rect 16222 17980 16286 17984
rect 16222 17924 16226 17980
rect 16226 17924 16282 17980
rect 16282 17924 16286 17980
rect 16222 17920 16286 17924
rect 4709 17436 4773 17440
rect 4709 17380 4713 17436
rect 4713 17380 4769 17436
rect 4769 17380 4773 17436
rect 4709 17376 4773 17380
rect 4789 17436 4853 17440
rect 4789 17380 4793 17436
rect 4793 17380 4849 17436
rect 4849 17380 4853 17436
rect 4789 17376 4853 17380
rect 4869 17436 4933 17440
rect 4869 17380 4873 17436
rect 4873 17380 4929 17436
rect 4929 17380 4933 17436
rect 4869 17376 4933 17380
rect 4949 17436 5013 17440
rect 4949 17380 4953 17436
rect 4953 17380 5009 17436
rect 5009 17380 5013 17436
rect 4949 17376 5013 17380
rect 12225 17436 12289 17440
rect 12225 17380 12229 17436
rect 12229 17380 12285 17436
rect 12285 17380 12289 17436
rect 12225 17376 12289 17380
rect 12305 17436 12369 17440
rect 12305 17380 12309 17436
rect 12309 17380 12365 17436
rect 12365 17380 12369 17436
rect 12305 17376 12369 17380
rect 12385 17436 12449 17440
rect 12385 17380 12389 17436
rect 12389 17380 12445 17436
rect 12445 17380 12449 17436
rect 12385 17376 12449 17380
rect 12465 17436 12529 17440
rect 12465 17380 12469 17436
rect 12469 17380 12525 17436
rect 12525 17380 12529 17436
rect 12465 17376 12529 17380
rect 19740 17436 19804 17440
rect 19740 17380 19744 17436
rect 19744 17380 19800 17436
rect 19800 17380 19804 17436
rect 19740 17376 19804 17380
rect 19820 17436 19884 17440
rect 19820 17380 19824 17436
rect 19824 17380 19880 17436
rect 19880 17380 19884 17436
rect 19820 17376 19884 17380
rect 19900 17436 19964 17440
rect 19900 17380 19904 17436
rect 19904 17380 19960 17436
rect 19960 17380 19964 17436
rect 19900 17376 19964 17380
rect 19980 17436 20044 17440
rect 19980 17380 19984 17436
rect 19984 17380 20040 17436
rect 20040 17380 20044 17436
rect 19980 17376 20044 17380
rect 8467 16892 8531 16896
rect 8467 16836 8471 16892
rect 8471 16836 8527 16892
rect 8527 16836 8531 16892
rect 8467 16832 8531 16836
rect 8547 16892 8611 16896
rect 8547 16836 8551 16892
rect 8551 16836 8607 16892
rect 8607 16836 8611 16892
rect 8547 16832 8611 16836
rect 8627 16892 8691 16896
rect 8627 16836 8631 16892
rect 8631 16836 8687 16892
rect 8687 16836 8691 16892
rect 8627 16832 8691 16836
rect 8707 16892 8771 16896
rect 8707 16836 8711 16892
rect 8711 16836 8767 16892
rect 8767 16836 8771 16892
rect 8707 16832 8771 16836
rect 15982 16892 16046 16896
rect 15982 16836 15986 16892
rect 15986 16836 16042 16892
rect 16042 16836 16046 16892
rect 15982 16832 16046 16836
rect 16062 16892 16126 16896
rect 16062 16836 16066 16892
rect 16066 16836 16122 16892
rect 16122 16836 16126 16892
rect 16062 16832 16126 16836
rect 16142 16892 16206 16896
rect 16142 16836 16146 16892
rect 16146 16836 16202 16892
rect 16202 16836 16206 16892
rect 16142 16832 16206 16836
rect 16222 16892 16286 16896
rect 16222 16836 16226 16892
rect 16226 16836 16282 16892
rect 16282 16836 16286 16892
rect 16222 16832 16286 16836
rect 4709 16348 4773 16352
rect 4709 16292 4713 16348
rect 4713 16292 4769 16348
rect 4769 16292 4773 16348
rect 4709 16288 4773 16292
rect 4789 16348 4853 16352
rect 4789 16292 4793 16348
rect 4793 16292 4849 16348
rect 4849 16292 4853 16348
rect 4789 16288 4853 16292
rect 4869 16348 4933 16352
rect 4869 16292 4873 16348
rect 4873 16292 4929 16348
rect 4929 16292 4933 16348
rect 4869 16288 4933 16292
rect 4949 16348 5013 16352
rect 4949 16292 4953 16348
rect 4953 16292 5009 16348
rect 5009 16292 5013 16348
rect 4949 16288 5013 16292
rect 12225 16348 12289 16352
rect 12225 16292 12229 16348
rect 12229 16292 12285 16348
rect 12285 16292 12289 16348
rect 12225 16288 12289 16292
rect 12305 16348 12369 16352
rect 12305 16292 12309 16348
rect 12309 16292 12365 16348
rect 12365 16292 12369 16348
rect 12305 16288 12369 16292
rect 12385 16348 12449 16352
rect 12385 16292 12389 16348
rect 12389 16292 12445 16348
rect 12445 16292 12449 16348
rect 12385 16288 12449 16292
rect 12465 16348 12529 16352
rect 12465 16292 12469 16348
rect 12469 16292 12525 16348
rect 12525 16292 12529 16348
rect 12465 16288 12529 16292
rect 19740 16348 19804 16352
rect 19740 16292 19744 16348
rect 19744 16292 19800 16348
rect 19800 16292 19804 16348
rect 19740 16288 19804 16292
rect 19820 16348 19884 16352
rect 19820 16292 19824 16348
rect 19824 16292 19880 16348
rect 19880 16292 19884 16348
rect 19820 16288 19884 16292
rect 19900 16348 19964 16352
rect 19900 16292 19904 16348
rect 19904 16292 19960 16348
rect 19960 16292 19964 16348
rect 19900 16288 19964 16292
rect 19980 16348 20044 16352
rect 19980 16292 19984 16348
rect 19984 16292 20040 16348
rect 20040 16292 20044 16348
rect 19980 16288 20044 16292
rect 8467 15804 8531 15808
rect 8467 15748 8471 15804
rect 8471 15748 8527 15804
rect 8527 15748 8531 15804
rect 8467 15744 8531 15748
rect 8547 15804 8611 15808
rect 8547 15748 8551 15804
rect 8551 15748 8607 15804
rect 8607 15748 8611 15804
rect 8547 15744 8611 15748
rect 8627 15804 8691 15808
rect 8627 15748 8631 15804
rect 8631 15748 8687 15804
rect 8687 15748 8691 15804
rect 8627 15744 8691 15748
rect 8707 15804 8771 15808
rect 8707 15748 8711 15804
rect 8711 15748 8767 15804
rect 8767 15748 8771 15804
rect 8707 15744 8771 15748
rect 15982 15804 16046 15808
rect 15982 15748 15986 15804
rect 15986 15748 16042 15804
rect 16042 15748 16046 15804
rect 15982 15744 16046 15748
rect 16062 15804 16126 15808
rect 16062 15748 16066 15804
rect 16066 15748 16122 15804
rect 16122 15748 16126 15804
rect 16062 15744 16126 15748
rect 16142 15804 16206 15808
rect 16142 15748 16146 15804
rect 16146 15748 16202 15804
rect 16202 15748 16206 15804
rect 16142 15744 16206 15748
rect 16222 15804 16286 15808
rect 16222 15748 16226 15804
rect 16226 15748 16282 15804
rect 16282 15748 16286 15804
rect 16222 15744 16286 15748
rect 4709 15260 4773 15264
rect 4709 15204 4713 15260
rect 4713 15204 4769 15260
rect 4769 15204 4773 15260
rect 4709 15200 4773 15204
rect 4789 15260 4853 15264
rect 4789 15204 4793 15260
rect 4793 15204 4849 15260
rect 4849 15204 4853 15260
rect 4789 15200 4853 15204
rect 4869 15260 4933 15264
rect 4869 15204 4873 15260
rect 4873 15204 4929 15260
rect 4929 15204 4933 15260
rect 4869 15200 4933 15204
rect 4949 15260 5013 15264
rect 4949 15204 4953 15260
rect 4953 15204 5009 15260
rect 5009 15204 5013 15260
rect 4949 15200 5013 15204
rect 12225 15260 12289 15264
rect 12225 15204 12229 15260
rect 12229 15204 12285 15260
rect 12285 15204 12289 15260
rect 12225 15200 12289 15204
rect 12305 15260 12369 15264
rect 12305 15204 12309 15260
rect 12309 15204 12365 15260
rect 12365 15204 12369 15260
rect 12305 15200 12369 15204
rect 12385 15260 12449 15264
rect 12385 15204 12389 15260
rect 12389 15204 12445 15260
rect 12445 15204 12449 15260
rect 12385 15200 12449 15204
rect 12465 15260 12529 15264
rect 12465 15204 12469 15260
rect 12469 15204 12525 15260
rect 12525 15204 12529 15260
rect 12465 15200 12529 15204
rect 19740 15260 19804 15264
rect 19740 15204 19744 15260
rect 19744 15204 19800 15260
rect 19800 15204 19804 15260
rect 19740 15200 19804 15204
rect 19820 15260 19884 15264
rect 19820 15204 19824 15260
rect 19824 15204 19880 15260
rect 19880 15204 19884 15260
rect 19820 15200 19884 15204
rect 19900 15260 19964 15264
rect 19900 15204 19904 15260
rect 19904 15204 19960 15260
rect 19960 15204 19964 15260
rect 19900 15200 19964 15204
rect 19980 15260 20044 15264
rect 19980 15204 19984 15260
rect 19984 15204 20040 15260
rect 20040 15204 20044 15260
rect 19980 15200 20044 15204
rect 8467 14716 8531 14720
rect 8467 14660 8471 14716
rect 8471 14660 8527 14716
rect 8527 14660 8531 14716
rect 8467 14656 8531 14660
rect 8547 14716 8611 14720
rect 8547 14660 8551 14716
rect 8551 14660 8607 14716
rect 8607 14660 8611 14716
rect 8547 14656 8611 14660
rect 8627 14716 8691 14720
rect 8627 14660 8631 14716
rect 8631 14660 8687 14716
rect 8687 14660 8691 14716
rect 8627 14656 8691 14660
rect 8707 14716 8771 14720
rect 8707 14660 8711 14716
rect 8711 14660 8767 14716
rect 8767 14660 8771 14716
rect 8707 14656 8771 14660
rect 15982 14716 16046 14720
rect 15982 14660 15986 14716
rect 15986 14660 16042 14716
rect 16042 14660 16046 14716
rect 15982 14656 16046 14660
rect 16062 14716 16126 14720
rect 16062 14660 16066 14716
rect 16066 14660 16122 14716
rect 16122 14660 16126 14716
rect 16062 14656 16126 14660
rect 16142 14716 16206 14720
rect 16142 14660 16146 14716
rect 16146 14660 16202 14716
rect 16202 14660 16206 14716
rect 16142 14656 16206 14660
rect 16222 14716 16286 14720
rect 16222 14660 16226 14716
rect 16226 14660 16282 14716
rect 16282 14660 16286 14716
rect 16222 14656 16286 14660
rect 4709 14172 4773 14176
rect 4709 14116 4713 14172
rect 4713 14116 4769 14172
rect 4769 14116 4773 14172
rect 4709 14112 4773 14116
rect 4789 14172 4853 14176
rect 4789 14116 4793 14172
rect 4793 14116 4849 14172
rect 4849 14116 4853 14172
rect 4789 14112 4853 14116
rect 4869 14172 4933 14176
rect 4869 14116 4873 14172
rect 4873 14116 4929 14172
rect 4929 14116 4933 14172
rect 4869 14112 4933 14116
rect 4949 14172 5013 14176
rect 4949 14116 4953 14172
rect 4953 14116 5009 14172
rect 5009 14116 5013 14172
rect 4949 14112 5013 14116
rect 12225 14172 12289 14176
rect 12225 14116 12229 14172
rect 12229 14116 12285 14172
rect 12285 14116 12289 14172
rect 12225 14112 12289 14116
rect 12305 14172 12369 14176
rect 12305 14116 12309 14172
rect 12309 14116 12365 14172
rect 12365 14116 12369 14172
rect 12305 14112 12369 14116
rect 12385 14172 12449 14176
rect 12385 14116 12389 14172
rect 12389 14116 12445 14172
rect 12445 14116 12449 14172
rect 12385 14112 12449 14116
rect 12465 14172 12529 14176
rect 12465 14116 12469 14172
rect 12469 14116 12525 14172
rect 12525 14116 12529 14172
rect 12465 14112 12529 14116
rect 19740 14172 19804 14176
rect 19740 14116 19744 14172
rect 19744 14116 19800 14172
rect 19800 14116 19804 14172
rect 19740 14112 19804 14116
rect 19820 14172 19884 14176
rect 19820 14116 19824 14172
rect 19824 14116 19880 14172
rect 19880 14116 19884 14172
rect 19820 14112 19884 14116
rect 19900 14172 19964 14176
rect 19900 14116 19904 14172
rect 19904 14116 19960 14172
rect 19960 14116 19964 14172
rect 19900 14112 19964 14116
rect 19980 14172 20044 14176
rect 19980 14116 19984 14172
rect 19984 14116 20040 14172
rect 20040 14116 20044 14172
rect 19980 14112 20044 14116
rect 8467 13628 8531 13632
rect 8467 13572 8471 13628
rect 8471 13572 8527 13628
rect 8527 13572 8531 13628
rect 8467 13568 8531 13572
rect 8547 13628 8611 13632
rect 8547 13572 8551 13628
rect 8551 13572 8607 13628
rect 8607 13572 8611 13628
rect 8547 13568 8611 13572
rect 8627 13628 8691 13632
rect 8627 13572 8631 13628
rect 8631 13572 8687 13628
rect 8687 13572 8691 13628
rect 8627 13568 8691 13572
rect 8707 13628 8771 13632
rect 8707 13572 8711 13628
rect 8711 13572 8767 13628
rect 8767 13572 8771 13628
rect 8707 13568 8771 13572
rect 15982 13628 16046 13632
rect 15982 13572 15986 13628
rect 15986 13572 16042 13628
rect 16042 13572 16046 13628
rect 15982 13568 16046 13572
rect 16062 13628 16126 13632
rect 16062 13572 16066 13628
rect 16066 13572 16122 13628
rect 16122 13572 16126 13628
rect 16062 13568 16126 13572
rect 16142 13628 16206 13632
rect 16142 13572 16146 13628
rect 16146 13572 16202 13628
rect 16202 13572 16206 13628
rect 16142 13568 16206 13572
rect 16222 13628 16286 13632
rect 16222 13572 16226 13628
rect 16226 13572 16282 13628
rect 16282 13572 16286 13628
rect 16222 13568 16286 13572
rect 22140 13092 22204 13156
rect 4709 13084 4773 13088
rect 4709 13028 4713 13084
rect 4713 13028 4769 13084
rect 4769 13028 4773 13084
rect 4709 13024 4773 13028
rect 4789 13084 4853 13088
rect 4789 13028 4793 13084
rect 4793 13028 4849 13084
rect 4849 13028 4853 13084
rect 4789 13024 4853 13028
rect 4869 13084 4933 13088
rect 4869 13028 4873 13084
rect 4873 13028 4929 13084
rect 4929 13028 4933 13084
rect 4869 13024 4933 13028
rect 4949 13084 5013 13088
rect 4949 13028 4953 13084
rect 4953 13028 5009 13084
rect 5009 13028 5013 13084
rect 4949 13024 5013 13028
rect 12225 13084 12289 13088
rect 12225 13028 12229 13084
rect 12229 13028 12285 13084
rect 12285 13028 12289 13084
rect 12225 13024 12289 13028
rect 12305 13084 12369 13088
rect 12305 13028 12309 13084
rect 12309 13028 12365 13084
rect 12365 13028 12369 13084
rect 12305 13024 12369 13028
rect 12385 13084 12449 13088
rect 12385 13028 12389 13084
rect 12389 13028 12445 13084
rect 12445 13028 12449 13084
rect 12385 13024 12449 13028
rect 12465 13084 12529 13088
rect 12465 13028 12469 13084
rect 12469 13028 12525 13084
rect 12525 13028 12529 13084
rect 12465 13024 12529 13028
rect 19740 13084 19804 13088
rect 19740 13028 19744 13084
rect 19744 13028 19800 13084
rect 19800 13028 19804 13084
rect 19740 13024 19804 13028
rect 19820 13084 19884 13088
rect 19820 13028 19824 13084
rect 19824 13028 19880 13084
rect 19880 13028 19884 13084
rect 19820 13024 19884 13028
rect 19900 13084 19964 13088
rect 19900 13028 19904 13084
rect 19904 13028 19960 13084
rect 19960 13028 19964 13084
rect 19900 13024 19964 13028
rect 19980 13084 20044 13088
rect 19980 13028 19984 13084
rect 19984 13028 20040 13084
rect 20040 13028 20044 13084
rect 19980 13024 20044 13028
rect 22140 12820 22204 12884
rect 8467 12540 8531 12544
rect 8467 12484 8471 12540
rect 8471 12484 8527 12540
rect 8527 12484 8531 12540
rect 8467 12480 8531 12484
rect 8547 12540 8611 12544
rect 8547 12484 8551 12540
rect 8551 12484 8607 12540
rect 8607 12484 8611 12540
rect 8547 12480 8611 12484
rect 8627 12540 8691 12544
rect 8627 12484 8631 12540
rect 8631 12484 8687 12540
rect 8687 12484 8691 12540
rect 8627 12480 8691 12484
rect 8707 12540 8771 12544
rect 8707 12484 8711 12540
rect 8711 12484 8767 12540
rect 8767 12484 8771 12540
rect 8707 12480 8771 12484
rect 15982 12540 16046 12544
rect 15982 12484 15986 12540
rect 15986 12484 16042 12540
rect 16042 12484 16046 12540
rect 15982 12480 16046 12484
rect 16062 12540 16126 12544
rect 16062 12484 16066 12540
rect 16066 12484 16122 12540
rect 16122 12484 16126 12540
rect 16062 12480 16126 12484
rect 16142 12540 16206 12544
rect 16142 12484 16146 12540
rect 16146 12484 16202 12540
rect 16202 12484 16206 12540
rect 16142 12480 16206 12484
rect 16222 12540 16286 12544
rect 16222 12484 16226 12540
rect 16226 12484 16282 12540
rect 16282 12484 16286 12540
rect 16222 12480 16286 12484
rect 4709 11996 4773 12000
rect 4709 11940 4713 11996
rect 4713 11940 4769 11996
rect 4769 11940 4773 11996
rect 4709 11936 4773 11940
rect 4789 11996 4853 12000
rect 4789 11940 4793 11996
rect 4793 11940 4849 11996
rect 4849 11940 4853 11996
rect 4789 11936 4853 11940
rect 4869 11996 4933 12000
rect 4869 11940 4873 11996
rect 4873 11940 4929 11996
rect 4929 11940 4933 11996
rect 4869 11936 4933 11940
rect 4949 11996 5013 12000
rect 4949 11940 4953 11996
rect 4953 11940 5009 11996
rect 5009 11940 5013 11996
rect 4949 11936 5013 11940
rect 12225 11996 12289 12000
rect 12225 11940 12229 11996
rect 12229 11940 12285 11996
rect 12285 11940 12289 11996
rect 12225 11936 12289 11940
rect 12305 11996 12369 12000
rect 12305 11940 12309 11996
rect 12309 11940 12365 11996
rect 12365 11940 12369 11996
rect 12305 11936 12369 11940
rect 12385 11996 12449 12000
rect 12385 11940 12389 11996
rect 12389 11940 12445 11996
rect 12445 11940 12449 11996
rect 12385 11936 12449 11940
rect 12465 11996 12529 12000
rect 12465 11940 12469 11996
rect 12469 11940 12525 11996
rect 12525 11940 12529 11996
rect 12465 11936 12529 11940
rect 19740 11996 19804 12000
rect 19740 11940 19744 11996
rect 19744 11940 19800 11996
rect 19800 11940 19804 11996
rect 19740 11936 19804 11940
rect 19820 11996 19884 12000
rect 19820 11940 19824 11996
rect 19824 11940 19880 11996
rect 19880 11940 19884 11996
rect 19820 11936 19884 11940
rect 19900 11996 19964 12000
rect 19900 11940 19904 11996
rect 19904 11940 19960 11996
rect 19960 11940 19964 11996
rect 19900 11936 19964 11940
rect 19980 11996 20044 12000
rect 19980 11940 19984 11996
rect 19984 11940 20040 11996
rect 20040 11940 20044 11996
rect 19980 11936 20044 11940
rect 60 11868 124 11932
rect 60 11596 124 11660
rect 8467 11452 8531 11456
rect 8467 11396 8471 11452
rect 8471 11396 8527 11452
rect 8527 11396 8531 11452
rect 8467 11392 8531 11396
rect 8547 11452 8611 11456
rect 8547 11396 8551 11452
rect 8551 11396 8607 11452
rect 8607 11396 8611 11452
rect 8547 11392 8611 11396
rect 8627 11452 8691 11456
rect 8627 11396 8631 11452
rect 8631 11396 8687 11452
rect 8687 11396 8691 11452
rect 8627 11392 8691 11396
rect 8707 11452 8771 11456
rect 8707 11396 8711 11452
rect 8711 11396 8767 11452
rect 8767 11396 8771 11452
rect 8707 11392 8771 11396
rect 15982 11452 16046 11456
rect 15982 11396 15986 11452
rect 15986 11396 16042 11452
rect 16042 11396 16046 11452
rect 15982 11392 16046 11396
rect 16062 11452 16126 11456
rect 16062 11396 16066 11452
rect 16066 11396 16122 11452
rect 16122 11396 16126 11452
rect 16062 11392 16126 11396
rect 16142 11452 16206 11456
rect 16142 11396 16146 11452
rect 16146 11396 16202 11452
rect 16202 11396 16206 11452
rect 16142 11392 16206 11396
rect 16222 11452 16286 11456
rect 16222 11396 16226 11452
rect 16226 11396 16282 11452
rect 16282 11396 16286 11452
rect 16222 11392 16286 11396
rect 4709 10908 4773 10912
rect 4709 10852 4713 10908
rect 4713 10852 4769 10908
rect 4769 10852 4773 10908
rect 4709 10848 4773 10852
rect 4789 10908 4853 10912
rect 4789 10852 4793 10908
rect 4793 10852 4849 10908
rect 4849 10852 4853 10908
rect 4789 10848 4853 10852
rect 4869 10908 4933 10912
rect 4869 10852 4873 10908
rect 4873 10852 4929 10908
rect 4929 10852 4933 10908
rect 4869 10848 4933 10852
rect 4949 10908 5013 10912
rect 4949 10852 4953 10908
rect 4953 10852 5009 10908
rect 5009 10852 5013 10908
rect 4949 10848 5013 10852
rect 12225 10908 12289 10912
rect 12225 10852 12229 10908
rect 12229 10852 12285 10908
rect 12285 10852 12289 10908
rect 12225 10848 12289 10852
rect 12305 10908 12369 10912
rect 12305 10852 12309 10908
rect 12309 10852 12365 10908
rect 12365 10852 12369 10908
rect 12305 10848 12369 10852
rect 12385 10908 12449 10912
rect 12385 10852 12389 10908
rect 12389 10852 12445 10908
rect 12445 10852 12449 10908
rect 12385 10848 12449 10852
rect 12465 10908 12529 10912
rect 12465 10852 12469 10908
rect 12469 10852 12525 10908
rect 12525 10852 12529 10908
rect 12465 10848 12529 10852
rect 19740 10908 19804 10912
rect 19740 10852 19744 10908
rect 19744 10852 19800 10908
rect 19800 10852 19804 10908
rect 19740 10848 19804 10852
rect 19820 10908 19884 10912
rect 19820 10852 19824 10908
rect 19824 10852 19880 10908
rect 19880 10852 19884 10908
rect 19820 10848 19884 10852
rect 19900 10908 19964 10912
rect 19900 10852 19904 10908
rect 19904 10852 19960 10908
rect 19960 10852 19964 10908
rect 19900 10848 19964 10852
rect 19980 10908 20044 10912
rect 19980 10852 19984 10908
rect 19984 10852 20040 10908
rect 20040 10852 20044 10908
rect 19980 10848 20044 10852
rect 22140 10644 22204 10708
rect 22140 10372 22204 10436
rect 8467 10364 8531 10368
rect 8467 10308 8471 10364
rect 8471 10308 8527 10364
rect 8527 10308 8531 10364
rect 8467 10304 8531 10308
rect 8547 10364 8611 10368
rect 8547 10308 8551 10364
rect 8551 10308 8607 10364
rect 8607 10308 8611 10364
rect 8547 10304 8611 10308
rect 8627 10364 8691 10368
rect 8627 10308 8631 10364
rect 8631 10308 8687 10364
rect 8687 10308 8691 10364
rect 8627 10304 8691 10308
rect 8707 10364 8771 10368
rect 8707 10308 8711 10364
rect 8711 10308 8767 10364
rect 8767 10308 8771 10364
rect 8707 10304 8771 10308
rect 15982 10364 16046 10368
rect 15982 10308 15986 10364
rect 15986 10308 16042 10364
rect 16042 10308 16046 10364
rect 15982 10304 16046 10308
rect 16062 10364 16126 10368
rect 16062 10308 16066 10364
rect 16066 10308 16122 10364
rect 16122 10308 16126 10364
rect 16062 10304 16126 10308
rect 16142 10364 16206 10368
rect 16142 10308 16146 10364
rect 16146 10308 16202 10364
rect 16202 10308 16206 10364
rect 16142 10304 16206 10308
rect 16222 10364 16286 10368
rect 16222 10308 16226 10364
rect 16226 10308 16282 10364
rect 16282 10308 16286 10364
rect 16222 10304 16286 10308
rect 4709 9820 4773 9824
rect 4709 9764 4713 9820
rect 4713 9764 4769 9820
rect 4769 9764 4773 9820
rect 4709 9760 4773 9764
rect 4789 9820 4853 9824
rect 4789 9764 4793 9820
rect 4793 9764 4849 9820
rect 4849 9764 4853 9820
rect 4789 9760 4853 9764
rect 4869 9820 4933 9824
rect 4869 9764 4873 9820
rect 4873 9764 4929 9820
rect 4929 9764 4933 9820
rect 4869 9760 4933 9764
rect 4949 9820 5013 9824
rect 4949 9764 4953 9820
rect 4953 9764 5009 9820
rect 5009 9764 5013 9820
rect 4949 9760 5013 9764
rect 12225 9820 12289 9824
rect 12225 9764 12229 9820
rect 12229 9764 12285 9820
rect 12285 9764 12289 9820
rect 12225 9760 12289 9764
rect 12305 9820 12369 9824
rect 12305 9764 12309 9820
rect 12309 9764 12365 9820
rect 12365 9764 12369 9820
rect 12305 9760 12369 9764
rect 12385 9820 12449 9824
rect 12385 9764 12389 9820
rect 12389 9764 12445 9820
rect 12445 9764 12449 9820
rect 12385 9760 12449 9764
rect 12465 9820 12529 9824
rect 12465 9764 12469 9820
rect 12469 9764 12525 9820
rect 12525 9764 12529 9820
rect 12465 9760 12529 9764
rect 19740 9820 19804 9824
rect 19740 9764 19744 9820
rect 19744 9764 19800 9820
rect 19800 9764 19804 9820
rect 19740 9760 19804 9764
rect 19820 9820 19884 9824
rect 19820 9764 19824 9820
rect 19824 9764 19880 9820
rect 19880 9764 19884 9820
rect 19820 9760 19884 9764
rect 19900 9820 19964 9824
rect 19900 9764 19904 9820
rect 19904 9764 19960 9820
rect 19960 9764 19964 9820
rect 19900 9760 19964 9764
rect 19980 9820 20044 9824
rect 19980 9764 19984 9820
rect 19984 9764 20040 9820
rect 20040 9764 20044 9820
rect 19980 9760 20044 9764
rect 8467 9276 8531 9280
rect 8467 9220 8471 9276
rect 8471 9220 8527 9276
rect 8527 9220 8531 9276
rect 8467 9216 8531 9220
rect 8547 9276 8611 9280
rect 8547 9220 8551 9276
rect 8551 9220 8607 9276
rect 8607 9220 8611 9276
rect 8547 9216 8611 9220
rect 8627 9276 8691 9280
rect 8627 9220 8631 9276
rect 8631 9220 8687 9276
rect 8687 9220 8691 9276
rect 8627 9216 8691 9220
rect 8707 9276 8771 9280
rect 8707 9220 8711 9276
rect 8711 9220 8767 9276
rect 8767 9220 8771 9276
rect 8707 9216 8771 9220
rect 15982 9276 16046 9280
rect 15982 9220 15986 9276
rect 15986 9220 16042 9276
rect 16042 9220 16046 9276
rect 15982 9216 16046 9220
rect 16062 9276 16126 9280
rect 16062 9220 16066 9276
rect 16066 9220 16122 9276
rect 16122 9220 16126 9276
rect 16062 9216 16126 9220
rect 16142 9276 16206 9280
rect 16142 9220 16146 9276
rect 16146 9220 16202 9276
rect 16202 9220 16206 9276
rect 16142 9216 16206 9220
rect 16222 9276 16286 9280
rect 16222 9220 16226 9276
rect 16226 9220 16282 9276
rect 16282 9220 16286 9276
rect 16222 9216 16286 9220
rect 4709 8732 4773 8736
rect 4709 8676 4713 8732
rect 4713 8676 4769 8732
rect 4769 8676 4773 8732
rect 4709 8672 4773 8676
rect 4789 8732 4853 8736
rect 4789 8676 4793 8732
rect 4793 8676 4849 8732
rect 4849 8676 4853 8732
rect 4789 8672 4853 8676
rect 4869 8732 4933 8736
rect 4869 8676 4873 8732
rect 4873 8676 4929 8732
rect 4929 8676 4933 8732
rect 4869 8672 4933 8676
rect 4949 8732 5013 8736
rect 4949 8676 4953 8732
rect 4953 8676 5009 8732
rect 5009 8676 5013 8732
rect 4949 8672 5013 8676
rect 12225 8732 12289 8736
rect 12225 8676 12229 8732
rect 12229 8676 12285 8732
rect 12285 8676 12289 8732
rect 12225 8672 12289 8676
rect 12305 8732 12369 8736
rect 12305 8676 12309 8732
rect 12309 8676 12365 8732
rect 12365 8676 12369 8732
rect 12305 8672 12369 8676
rect 12385 8732 12449 8736
rect 12385 8676 12389 8732
rect 12389 8676 12445 8732
rect 12445 8676 12449 8732
rect 12385 8672 12449 8676
rect 12465 8732 12529 8736
rect 12465 8676 12469 8732
rect 12469 8676 12525 8732
rect 12525 8676 12529 8732
rect 12465 8672 12529 8676
rect 19740 8732 19804 8736
rect 19740 8676 19744 8732
rect 19744 8676 19800 8732
rect 19800 8676 19804 8732
rect 19740 8672 19804 8676
rect 19820 8732 19884 8736
rect 19820 8676 19824 8732
rect 19824 8676 19880 8732
rect 19880 8676 19884 8732
rect 19820 8672 19884 8676
rect 19900 8732 19964 8736
rect 19900 8676 19904 8732
rect 19904 8676 19960 8732
rect 19960 8676 19964 8732
rect 19900 8672 19964 8676
rect 19980 8732 20044 8736
rect 19980 8676 19984 8732
rect 19984 8676 20040 8732
rect 20040 8676 20044 8732
rect 19980 8672 20044 8676
rect 8467 8188 8531 8192
rect 8467 8132 8471 8188
rect 8471 8132 8527 8188
rect 8527 8132 8531 8188
rect 8467 8128 8531 8132
rect 8547 8188 8611 8192
rect 8547 8132 8551 8188
rect 8551 8132 8607 8188
rect 8607 8132 8611 8188
rect 8547 8128 8611 8132
rect 8627 8188 8691 8192
rect 8627 8132 8631 8188
rect 8631 8132 8687 8188
rect 8687 8132 8691 8188
rect 8627 8128 8691 8132
rect 8707 8188 8771 8192
rect 8707 8132 8711 8188
rect 8711 8132 8767 8188
rect 8767 8132 8771 8188
rect 8707 8128 8771 8132
rect 15982 8188 16046 8192
rect 15982 8132 15986 8188
rect 15986 8132 16042 8188
rect 16042 8132 16046 8188
rect 15982 8128 16046 8132
rect 16062 8188 16126 8192
rect 16062 8132 16066 8188
rect 16066 8132 16122 8188
rect 16122 8132 16126 8188
rect 16062 8128 16126 8132
rect 16142 8188 16206 8192
rect 16142 8132 16146 8188
rect 16146 8132 16202 8188
rect 16202 8132 16206 8188
rect 16142 8128 16206 8132
rect 16222 8188 16286 8192
rect 16222 8132 16226 8188
rect 16226 8132 16282 8188
rect 16282 8132 16286 8188
rect 16222 8128 16286 8132
rect 4709 7644 4773 7648
rect 4709 7588 4713 7644
rect 4713 7588 4769 7644
rect 4769 7588 4773 7644
rect 4709 7584 4773 7588
rect 4789 7644 4853 7648
rect 4789 7588 4793 7644
rect 4793 7588 4849 7644
rect 4849 7588 4853 7644
rect 4789 7584 4853 7588
rect 4869 7644 4933 7648
rect 4869 7588 4873 7644
rect 4873 7588 4929 7644
rect 4929 7588 4933 7644
rect 4869 7584 4933 7588
rect 4949 7644 5013 7648
rect 4949 7588 4953 7644
rect 4953 7588 5009 7644
rect 5009 7588 5013 7644
rect 4949 7584 5013 7588
rect 12225 7644 12289 7648
rect 12225 7588 12229 7644
rect 12229 7588 12285 7644
rect 12285 7588 12289 7644
rect 12225 7584 12289 7588
rect 12305 7644 12369 7648
rect 12305 7588 12309 7644
rect 12309 7588 12365 7644
rect 12365 7588 12369 7644
rect 12305 7584 12369 7588
rect 12385 7644 12449 7648
rect 12385 7588 12389 7644
rect 12389 7588 12445 7644
rect 12445 7588 12449 7644
rect 12385 7584 12449 7588
rect 12465 7644 12529 7648
rect 12465 7588 12469 7644
rect 12469 7588 12525 7644
rect 12525 7588 12529 7644
rect 12465 7584 12529 7588
rect 19740 7644 19804 7648
rect 19740 7588 19744 7644
rect 19744 7588 19800 7644
rect 19800 7588 19804 7644
rect 19740 7584 19804 7588
rect 19820 7644 19884 7648
rect 19820 7588 19824 7644
rect 19824 7588 19880 7644
rect 19880 7588 19884 7644
rect 19820 7584 19884 7588
rect 19900 7644 19964 7648
rect 19900 7588 19904 7644
rect 19904 7588 19960 7644
rect 19960 7588 19964 7644
rect 19900 7584 19964 7588
rect 19980 7644 20044 7648
rect 19980 7588 19984 7644
rect 19984 7588 20040 7644
rect 20040 7588 20044 7644
rect 19980 7584 20044 7588
rect 8467 7100 8531 7104
rect 8467 7044 8471 7100
rect 8471 7044 8527 7100
rect 8527 7044 8531 7100
rect 8467 7040 8531 7044
rect 8547 7100 8611 7104
rect 8547 7044 8551 7100
rect 8551 7044 8607 7100
rect 8607 7044 8611 7100
rect 8547 7040 8611 7044
rect 8627 7100 8691 7104
rect 8627 7044 8631 7100
rect 8631 7044 8687 7100
rect 8687 7044 8691 7100
rect 8627 7040 8691 7044
rect 8707 7100 8771 7104
rect 8707 7044 8711 7100
rect 8711 7044 8767 7100
rect 8767 7044 8771 7100
rect 8707 7040 8771 7044
rect 15982 7100 16046 7104
rect 15982 7044 15986 7100
rect 15986 7044 16042 7100
rect 16042 7044 16046 7100
rect 15982 7040 16046 7044
rect 16062 7100 16126 7104
rect 16062 7044 16066 7100
rect 16066 7044 16122 7100
rect 16122 7044 16126 7100
rect 16062 7040 16126 7044
rect 16142 7100 16206 7104
rect 16142 7044 16146 7100
rect 16146 7044 16202 7100
rect 16202 7044 16206 7100
rect 16142 7040 16206 7044
rect 16222 7100 16286 7104
rect 16222 7044 16226 7100
rect 16226 7044 16282 7100
rect 16282 7044 16286 7100
rect 16222 7040 16286 7044
rect 4709 6556 4773 6560
rect 4709 6500 4713 6556
rect 4713 6500 4769 6556
rect 4769 6500 4773 6556
rect 4709 6496 4773 6500
rect 4789 6556 4853 6560
rect 4789 6500 4793 6556
rect 4793 6500 4849 6556
rect 4849 6500 4853 6556
rect 4789 6496 4853 6500
rect 4869 6556 4933 6560
rect 4869 6500 4873 6556
rect 4873 6500 4929 6556
rect 4929 6500 4933 6556
rect 4869 6496 4933 6500
rect 4949 6556 5013 6560
rect 4949 6500 4953 6556
rect 4953 6500 5009 6556
rect 5009 6500 5013 6556
rect 4949 6496 5013 6500
rect 12225 6556 12289 6560
rect 12225 6500 12229 6556
rect 12229 6500 12285 6556
rect 12285 6500 12289 6556
rect 12225 6496 12289 6500
rect 12305 6556 12369 6560
rect 12305 6500 12309 6556
rect 12309 6500 12365 6556
rect 12365 6500 12369 6556
rect 12305 6496 12369 6500
rect 12385 6556 12449 6560
rect 12385 6500 12389 6556
rect 12389 6500 12445 6556
rect 12445 6500 12449 6556
rect 12385 6496 12449 6500
rect 12465 6556 12529 6560
rect 12465 6500 12469 6556
rect 12469 6500 12525 6556
rect 12525 6500 12529 6556
rect 12465 6496 12529 6500
rect 19740 6556 19804 6560
rect 19740 6500 19744 6556
rect 19744 6500 19800 6556
rect 19800 6500 19804 6556
rect 19740 6496 19804 6500
rect 19820 6556 19884 6560
rect 19820 6500 19824 6556
rect 19824 6500 19880 6556
rect 19880 6500 19884 6556
rect 19820 6496 19884 6500
rect 19900 6556 19964 6560
rect 19900 6500 19904 6556
rect 19904 6500 19960 6556
rect 19960 6500 19964 6556
rect 19900 6496 19964 6500
rect 19980 6556 20044 6560
rect 19980 6500 19984 6556
rect 19984 6500 20040 6556
rect 20040 6500 20044 6556
rect 19980 6496 20044 6500
rect 8467 6012 8531 6016
rect 8467 5956 8471 6012
rect 8471 5956 8527 6012
rect 8527 5956 8531 6012
rect 8467 5952 8531 5956
rect 8547 6012 8611 6016
rect 8547 5956 8551 6012
rect 8551 5956 8607 6012
rect 8607 5956 8611 6012
rect 8547 5952 8611 5956
rect 8627 6012 8691 6016
rect 8627 5956 8631 6012
rect 8631 5956 8687 6012
rect 8687 5956 8691 6012
rect 8627 5952 8691 5956
rect 8707 6012 8771 6016
rect 8707 5956 8711 6012
rect 8711 5956 8767 6012
rect 8767 5956 8771 6012
rect 8707 5952 8771 5956
rect 15982 6012 16046 6016
rect 15982 5956 15986 6012
rect 15986 5956 16042 6012
rect 16042 5956 16046 6012
rect 15982 5952 16046 5956
rect 16062 6012 16126 6016
rect 16062 5956 16066 6012
rect 16066 5956 16122 6012
rect 16122 5956 16126 6012
rect 16062 5952 16126 5956
rect 16142 6012 16206 6016
rect 16142 5956 16146 6012
rect 16146 5956 16202 6012
rect 16202 5956 16206 6012
rect 16142 5952 16206 5956
rect 16222 6012 16286 6016
rect 16222 5956 16226 6012
rect 16226 5956 16282 6012
rect 16282 5956 16286 6012
rect 16222 5952 16286 5956
rect 4709 5468 4773 5472
rect 4709 5412 4713 5468
rect 4713 5412 4769 5468
rect 4769 5412 4773 5468
rect 4709 5408 4773 5412
rect 4789 5468 4853 5472
rect 4789 5412 4793 5468
rect 4793 5412 4849 5468
rect 4849 5412 4853 5468
rect 4789 5408 4853 5412
rect 4869 5468 4933 5472
rect 4869 5412 4873 5468
rect 4873 5412 4929 5468
rect 4929 5412 4933 5468
rect 4869 5408 4933 5412
rect 4949 5468 5013 5472
rect 4949 5412 4953 5468
rect 4953 5412 5009 5468
rect 5009 5412 5013 5468
rect 4949 5408 5013 5412
rect 12225 5468 12289 5472
rect 12225 5412 12229 5468
rect 12229 5412 12285 5468
rect 12285 5412 12289 5468
rect 12225 5408 12289 5412
rect 12305 5468 12369 5472
rect 12305 5412 12309 5468
rect 12309 5412 12365 5468
rect 12365 5412 12369 5468
rect 12305 5408 12369 5412
rect 12385 5468 12449 5472
rect 12385 5412 12389 5468
rect 12389 5412 12445 5468
rect 12445 5412 12449 5468
rect 12385 5408 12449 5412
rect 12465 5468 12529 5472
rect 12465 5412 12469 5468
rect 12469 5412 12525 5468
rect 12525 5412 12529 5468
rect 12465 5408 12529 5412
rect 19740 5468 19804 5472
rect 19740 5412 19744 5468
rect 19744 5412 19800 5468
rect 19800 5412 19804 5468
rect 19740 5408 19804 5412
rect 19820 5468 19884 5472
rect 19820 5412 19824 5468
rect 19824 5412 19880 5468
rect 19880 5412 19884 5468
rect 19820 5408 19884 5412
rect 19900 5468 19964 5472
rect 19900 5412 19904 5468
rect 19904 5412 19960 5468
rect 19960 5412 19964 5468
rect 19900 5408 19964 5412
rect 19980 5468 20044 5472
rect 19980 5412 19984 5468
rect 19984 5412 20040 5468
rect 20040 5412 20044 5468
rect 19980 5408 20044 5412
rect 8467 4924 8531 4928
rect 8467 4868 8471 4924
rect 8471 4868 8527 4924
rect 8527 4868 8531 4924
rect 8467 4864 8531 4868
rect 8547 4924 8611 4928
rect 8547 4868 8551 4924
rect 8551 4868 8607 4924
rect 8607 4868 8611 4924
rect 8547 4864 8611 4868
rect 8627 4924 8691 4928
rect 8627 4868 8631 4924
rect 8631 4868 8687 4924
rect 8687 4868 8691 4924
rect 8627 4864 8691 4868
rect 8707 4924 8771 4928
rect 8707 4868 8711 4924
rect 8711 4868 8767 4924
rect 8767 4868 8771 4924
rect 8707 4864 8771 4868
rect 15982 4924 16046 4928
rect 15982 4868 15986 4924
rect 15986 4868 16042 4924
rect 16042 4868 16046 4924
rect 15982 4864 16046 4868
rect 16062 4924 16126 4928
rect 16062 4868 16066 4924
rect 16066 4868 16122 4924
rect 16122 4868 16126 4924
rect 16062 4864 16126 4868
rect 16142 4924 16206 4928
rect 16142 4868 16146 4924
rect 16146 4868 16202 4924
rect 16202 4868 16206 4924
rect 16142 4864 16206 4868
rect 16222 4924 16286 4928
rect 16222 4868 16226 4924
rect 16226 4868 16282 4924
rect 16282 4868 16286 4924
rect 16222 4864 16286 4868
rect 4709 4380 4773 4384
rect 4709 4324 4713 4380
rect 4713 4324 4769 4380
rect 4769 4324 4773 4380
rect 4709 4320 4773 4324
rect 4789 4380 4853 4384
rect 4789 4324 4793 4380
rect 4793 4324 4849 4380
rect 4849 4324 4853 4380
rect 4789 4320 4853 4324
rect 4869 4380 4933 4384
rect 4869 4324 4873 4380
rect 4873 4324 4929 4380
rect 4929 4324 4933 4380
rect 4869 4320 4933 4324
rect 4949 4380 5013 4384
rect 4949 4324 4953 4380
rect 4953 4324 5009 4380
rect 5009 4324 5013 4380
rect 4949 4320 5013 4324
rect 12225 4380 12289 4384
rect 12225 4324 12229 4380
rect 12229 4324 12285 4380
rect 12285 4324 12289 4380
rect 12225 4320 12289 4324
rect 12305 4380 12369 4384
rect 12305 4324 12309 4380
rect 12309 4324 12365 4380
rect 12365 4324 12369 4380
rect 12305 4320 12369 4324
rect 12385 4380 12449 4384
rect 12385 4324 12389 4380
rect 12389 4324 12445 4380
rect 12445 4324 12449 4380
rect 12385 4320 12449 4324
rect 12465 4380 12529 4384
rect 12465 4324 12469 4380
rect 12469 4324 12525 4380
rect 12525 4324 12529 4380
rect 12465 4320 12529 4324
rect 19740 4380 19804 4384
rect 19740 4324 19744 4380
rect 19744 4324 19800 4380
rect 19800 4324 19804 4380
rect 19740 4320 19804 4324
rect 19820 4380 19884 4384
rect 19820 4324 19824 4380
rect 19824 4324 19880 4380
rect 19880 4324 19884 4380
rect 19820 4320 19884 4324
rect 19900 4380 19964 4384
rect 19900 4324 19904 4380
rect 19904 4324 19960 4380
rect 19960 4324 19964 4380
rect 19900 4320 19964 4324
rect 19980 4380 20044 4384
rect 19980 4324 19984 4380
rect 19984 4324 20040 4380
rect 20040 4324 20044 4380
rect 19980 4320 20044 4324
rect 8467 3836 8531 3840
rect 8467 3780 8471 3836
rect 8471 3780 8527 3836
rect 8527 3780 8531 3836
rect 8467 3776 8531 3780
rect 8547 3836 8611 3840
rect 8547 3780 8551 3836
rect 8551 3780 8607 3836
rect 8607 3780 8611 3836
rect 8547 3776 8611 3780
rect 8627 3836 8691 3840
rect 8627 3780 8631 3836
rect 8631 3780 8687 3836
rect 8687 3780 8691 3836
rect 8627 3776 8691 3780
rect 8707 3836 8771 3840
rect 8707 3780 8711 3836
rect 8711 3780 8767 3836
rect 8767 3780 8771 3836
rect 8707 3776 8771 3780
rect 15982 3836 16046 3840
rect 15982 3780 15986 3836
rect 15986 3780 16042 3836
rect 16042 3780 16046 3836
rect 15982 3776 16046 3780
rect 16062 3836 16126 3840
rect 16062 3780 16066 3836
rect 16066 3780 16122 3836
rect 16122 3780 16126 3836
rect 16062 3776 16126 3780
rect 16142 3836 16206 3840
rect 16142 3780 16146 3836
rect 16146 3780 16202 3836
rect 16202 3780 16206 3836
rect 16142 3776 16206 3780
rect 16222 3836 16286 3840
rect 16222 3780 16226 3836
rect 16226 3780 16282 3836
rect 16282 3780 16286 3836
rect 16222 3776 16286 3780
rect 4709 3292 4773 3296
rect 4709 3236 4713 3292
rect 4713 3236 4769 3292
rect 4769 3236 4773 3292
rect 4709 3232 4773 3236
rect 4789 3292 4853 3296
rect 4789 3236 4793 3292
rect 4793 3236 4849 3292
rect 4849 3236 4853 3292
rect 4789 3232 4853 3236
rect 4869 3292 4933 3296
rect 4869 3236 4873 3292
rect 4873 3236 4929 3292
rect 4929 3236 4933 3292
rect 4869 3232 4933 3236
rect 4949 3292 5013 3296
rect 4949 3236 4953 3292
rect 4953 3236 5009 3292
rect 5009 3236 5013 3292
rect 4949 3232 5013 3236
rect 12225 3292 12289 3296
rect 12225 3236 12229 3292
rect 12229 3236 12285 3292
rect 12285 3236 12289 3292
rect 12225 3232 12289 3236
rect 12305 3292 12369 3296
rect 12305 3236 12309 3292
rect 12309 3236 12365 3292
rect 12365 3236 12369 3292
rect 12305 3232 12369 3236
rect 12385 3292 12449 3296
rect 12385 3236 12389 3292
rect 12389 3236 12445 3292
rect 12445 3236 12449 3292
rect 12385 3232 12449 3236
rect 12465 3292 12529 3296
rect 12465 3236 12469 3292
rect 12469 3236 12525 3292
rect 12525 3236 12529 3292
rect 12465 3232 12529 3236
rect 19740 3292 19804 3296
rect 19740 3236 19744 3292
rect 19744 3236 19800 3292
rect 19800 3236 19804 3292
rect 19740 3232 19804 3236
rect 19820 3292 19884 3296
rect 19820 3236 19824 3292
rect 19824 3236 19880 3292
rect 19880 3236 19884 3292
rect 19820 3232 19884 3236
rect 19900 3292 19964 3296
rect 19900 3236 19904 3292
rect 19904 3236 19960 3292
rect 19960 3236 19964 3292
rect 19900 3232 19964 3236
rect 19980 3292 20044 3296
rect 19980 3236 19984 3292
rect 19984 3236 20040 3292
rect 20040 3236 20044 3292
rect 19980 3232 20044 3236
rect 8467 2748 8531 2752
rect 8467 2692 8471 2748
rect 8471 2692 8527 2748
rect 8527 2692 8531 2748
rect 8467 2688 8531 2692
rect 8547 2748 8611 2752
rect 8547 2692 8551 2748
rect 8551 2692 8607 2748
rect 8607 2692 8611 2748
rect 8547 2688 8611 2692
rect 8627 2748 8691 2752
rect 8627 2692 8631 2748
rect 8631 2692 8687 2748
rect 8687 2692 8691 2748
rect 8627 2688 8691 2692
rect 8707 2748 8771 2752
rect 8707 2692 8711 2748
rect 8711 2692 8767 2748
rect 8767 2692 8771 2748
rect 8707 2688 8771 2692
rect 15982 2748 16046 2752
rect 15982 2692 15986 2748
rect 15986 2692 16042 2748
rect 16042 2692 16046 2748
rect 15982 2688 16046 2692
rect 16062 2748 16126 2752
rect 16062 2692 16066 2748
rect 16066 2692 16122 2748
rect 16122 2692 16126 2748
rect 16062 2688 16126 2692
rect 16142 2748 16206 2752
rect 16142 2692 16146 2748
rect 16146 2692 16202 2748
rect 16202 2692 16206 2748
rect 16142 2688 16206 2692
rect 16222 2748 16286 2752
rect 16222 2692 16226 2748
rect 16226 2692 16282 2748
rect 16282 2692 16286 2748
rect 16222 2688 16286 2692
rect 4709 2204 4773 2208
rect 4709 2148 4713 2204
rect 4713 2148 4769 2204
rect 4769 2148 4773 2204
rect 4709 2144 4773 2148
rect 4789 2204 4853 2208
rect 4789 2148 4793 2204
rect 4793 2148 4849 2204
rect 4849 2148 4853 2204
rect 4789 2144 4853 2148
rect 4869 2204 4933 2208
rect 4869 2148 4873 2204
rect 4873 2148 4929 2204
rect 4929 2148 4933 2204
rect 4869 2144 4933 2148
rect 4949 2204 5013 2208
rect 4949 2148 4953 2204
rect 4953 2148 5009 2204
rect 5009 2148 5013 2204
rect 4949 2144 5013 2148
rect 12225 2204 12289 2208
rect 12225 2148 12229 2204
rect 12229 2148 12285 2204
rect 12285 2148 12289 2204
rect 12225 2144 12289 2148
rect 12305 2204 12369 2208
rect 12305 2148 12309 2204
rect 12309 2148 12365 2204
rect 12365 2148 12369 2204
rect 12305 2144 12369 2148
rect 12385 2204 12449 2208
rect 12385 2148 12389 2204
rect 12389 2148 12445 2204
rect 12445 2148 12449 2204
rect 12385 2144 12449 2148
rect 12465 2204 12529 2208
rect 12465 2148 12469 2204
rect 12469 2148 12525 2204
rect 12525 2148 12529 2204
rect 12465 2144 12529 2148
rect 19740 2204 19804 2208
rect 19740 2148 19744 2204
rect 19744 2148 19800 2204
rect 19800 2148 19804 2204
rect 19740 2144 19804 2148
rect 19820 2204 19884 2208
rect 19820 2148 19824 2204
rect 19824 2148 19880 2204
rect 19880 2148 19884 2204
rect 19820 2144 19884 2148
rect 19900 2204 19964 2208
rect 19900 2148 19904 2204
rect 19904 2148 19960 2204
rect 19960 2148 19964 2204
rect 19900 2144 19964 2148
rect 19980 2204 20044 2208
rect 19980 2148 19984 2204
rect 19984 2148 20040 2204
rect 20040 2148 20044 2204
rect 19980 2144 20044 2148
<< metal4 >>
rect 4701 21792 5022 22352
rect 4701 21728 4709 21792
rect 4773 21728 4789 21792
rect 4853 21728 4869 21792
rect 4933 21728 4949 21792
rect 5013 21728 5022 21792
rect 4701 20704 5022 21728
rect 4701 20640 4709 20704
rect 4773 20640 4789 20704
rect 4853 20640 4869 20704
rect 4933 20640 4949 20704
rect 5013 20640 5022 20704
rect 4701 19616 5022 20640
rect 4701 19552 4709 19616
rect 4773 19552 4789 19616
rect 4853 19552 4869 19616
rect 4933 19552 4949 19616
rect 5013 19552 5022 19616
rect 4701 18528 5022 19552
rect 4701 18464 4709 18528
rect 4773 18464 4789 18528
rect 4853 18464 4869 18528
rect 4933 18464 4949 18528
rect 5013 18464 5022 18528
rect 4701 17440 5022 18464
rect 4701 17376 4709 17440
rect 4773 17376 4789 17440
rect 4853 17376 4869 17440
rect 4933 17376 4949 17440
rect 5013 17376 5022 17440
rect 4701 16352 5022 17376
rect 4701 16288 4709 16352
rect 4773 16288 4789 16352
rect 4853 16288 4869 16352
rect 4933 16288 4949 16352
rect 5013 16288 5022 16352
rect 4701 15264 5022 16288
rect 4701 15200 4709 15264
rect 4773 15200 4789 15264
rect 4853 15200 4869 15264
rect 4933 15200 4949 15264
rect 5013 15200 5022 15264
rect 4701 14176 5022 15200
rect 4701 14112 4709 14176
rect 4773 14112 4789 14176
rect 4853 14112 4869 14176
rect 4933 14112 4949 14176
rect 5013 14112 5022 14176
rect 4701 13088 5022 14112
rect 4701 13024 4709 13088
rect 4773 13024 4789 13088
rect 4853 13024 4869 13088
rect 4933 13024 4949 13088
rect 5013 13024 5022 13088
rect 4701 12000 5022 13024
rect 4701 11936 4709 12000
rect 4773 11936 4789 12000
rect 4853 11936 4869 12000
rect 4933 11936 4949 12000
rect 5013 11936 5022 12000
rect 59 11932 125 11933
rect 59 11868 60 11932
rect 124 11868 125 11932
rect 59 11867 125 11868
rect 62 11661 122 11867
rect 59 11660 125 11661
rect 59 11596 60 11660
rect 124 11596 125 11660
rect 59 11595 125 11596
rect 4701 10912 5022 11936
rect 4701 10848 4709 10912
rect 4773 10848 4789 10912
rect 4853 10848 4869 10912
rect 4933 10848 4949 10912
rect 5013 10848 5022 10912
rect 4701 9824 5022 10848
rect 4701 9760 4709 9824
rect 4773 9760 4789 9824
rect 4853 9760 4869 9824
rect 4933 9760 4949 9824
rect 5013 9760 5022 9824
rect 4701 8736 5022 9760
rect 4701 8672 4709 8736
rect 4773 8672 4789 8736
rect 4853 8672 4869 8736
rect 4933 8672 4949 8736
rect 5013 8672 5022 8736
rect 4701 7648 5022 8672
rect 4701 7584 4709 7648
rect 4773 7584 4789 7648
rect 4853 7584 4869 7648
rect 4933 7584 4949 7648
rect 5013 7584 5022 7648
rect 4701 6560 5022 7584
rect 4701 6496 4709 6560
rect 4773 6496 4789 6560
rect 4853 6496 4869 6560
rect 4933 6496 4949 6560
rect 5013 6496 5022 6560
rect 4701 5472 5022 6496
rect 4701 5408 4709 5472
rect 4773 5408 4789 5472
rect 4853 5408 4869 5472
rect 4933 5408 4949 5472
rect 5013 5408 5022 5472
rect 4701 4384 5022 5408
rect 4701 4320 4709 4384
rect 4773 4320 4789 4384
rect 4853 4320 4869 4384
rect 4933 4320 4949 4384
rect 5013 4320 5022 4384
rect 4701 3296 5022 4320
rect 4701 3232 4709 3296
rect 4773 3232 4789 3296
rect 4853 3232 4869 3296
rect 4933 3232 4949 3296
rect 5013 3232 5022 3296
rect 4701 2208 5022 3232
rect 4701 2144 4709 2208
rect 4773 2144 4789 2208
rect 4853 2144 4869 2208
rect 4933 2144 4949 2208
rect 5013 2144 5022 2208
rect 4701 2128 5022 2144
rect 8459 22336 8779 22352
rect 8459 22272 8467 22336
rect 8531 22272 8547 22336
rect 8611 22272 8627 22336
rect 8691 22272 8707 22336
rect 8771 22272 8779 22336
rect 8459 21248 8779 22272
rect 8459 21184 8467 21248
rect 8531 21184 8547 21248
rect 8611 21184 8627 21248
rect 8691 21184 8707 21248
rect 8771 21184 8779 21248
rect 8459 20160 8779 21184
rect 8459 20096 8467 20160
rect 8531 20096 8547 20160
rect 8611 20096 8627 20160
rect 8691 20096 8707 20160
rect 8771 20096 8779 20160
rect 8459 19072 8779 20096
rect 8459 19008 8467 19072
rect 8531 19008 8547 19072
rect 8611 19008 8627 19072
rect 8691 19008 8707 19072
rect 8771 19008 8779 19072
rect 8459 17984 8779 19008
rect 8459 17920 8467 17984
rect 8531 17920 8547 17984
rect 8611 17920 8627 17984
rect 8691 17920 8707 17984
rect 8771 17920 8779 17984
rect 8459 16896 8779 17920
rect 8459 16832 8467 16896
rect 8531 16832 8547 16896
rect 8611 16832 8627 16896
rect 8691 16832 8707 16896
rect 8771 16832 8779 16896
rect 8459 15808 8779 16832
rect 8459 15744 8467 15808
rect 8531 15744 8547 15808
rect 8611 15744 8627 15808
rect 8691 15744 8707 15808
rect 8771 15744 8779 15808
rect 8459 14720 8779 15744
rect 8459 14656 8467 14720
rect 8531 14656 8547 14720
rect 8611 14656 8627 14720
rect 8691 14656 8707 14720
rect 8771 14656 8779 14720
rect 8459 13632 8779 14656
rect 8459 13568 8467 13632
rect 8531 13568 8547 13632
rect 8611 13568 8627 13632
rect 8691 13568 8707 13632
rect 8771 13568 8779 13632
rect 8459 12544 8779 13568
rect 8459 12480 8467 12544
rect 8531 12480 8547 12544
rect 8611 12480 8627 12544
rect 8691 12480 8707 12544
rect 8771 12480 8779 12544
rect 8459 11456 8779 12480
rect 8459 11392 8467 11456
rect 8531 11392 8547 11456
rect 8611 11392 8627 11456
rect 8691 11392 8707 11456
rect 8771 11392 8779 11456
rect 8459 10368 8779 11392
rect 8459 10304 8467 10368
rect 8531 10304 8547 10368
rect 8611 10304 8627 10368
rect 8691 10304 8707 10368
rect 8771 10304 8779 10368
rect 8459 9280 8779 10304
rect 8459 9216 8467 9280
rect 8531 9216 8547 9280
rect 8611 9216 8627 9280
rect 8691 9216 8707 9280
rect 8771 9216 8779 9280
rect 8459 8192 8779 9216
rect 8459 8128 8467 8192
rect 8531 8128 8547 8192
rect 8611 8128 8627 8192
rect 8691 8128 8707 8192
rect 8771 8128 8779 8192
rect 8459 7104 8779 8128
rect 8459 7040 8467 7104
rect 8531 7040 8547 7104
rect 8611 7040 8627 7104
rect 8691 7040 8707 7104
rect 8771 7040 8779 7104
rect 8459 6016 8779 7040
rect 8459 5952 8467 6016
rect 8531 5952 8547 6016
rect 8611 5952 8627 6016
rect 8691 5952 8707 6016
rect 8771 5952 8779 6016
rect 8459 4928 8779 5952
rect 8459 4864 8467 4928
rect 8531 4864 8547 4928
rect 8611 4864 8627 4928
rect 8691 4864 8707 4928
rect 8771 4864 8779 4928
rect 8459 3840 8779 4864
rect 8459 3776 8467 3840
rect 8531 3776 8547 3840
rect 8611 3776 8627 3840
rect 8691 3776 8707 3840
rect 8771 3776 8779 3840
rect 8459 2752 8779 3776
rect 8459 2688 8467 2752
rect 8531 2688 8547 2752
rect 8611 2688 8627 2752
rect 8691 2688 8707 2752
rect 8771 2688 8779 2752
rect 8459 2128 8779 2688
rect 12217 21792 12537 22352
rect 12217 21728 12225 21792
rect 12289 21728 12305 21792
rect 12369 21728 12385 21792
rect 12449 21728 12465 21792
rect 12529 21728 12537 21792
rect 12217 20704 12537 21728
rect 12217 20640 12225 20704
rect 12289 20640 12305 20704
rect 12369 20640 12385 20704
rect 12449 20640 12465 20704
rect 12529 20640 12537 20704
rect 12217 19616 12537 20640
rect 12217 19552 12225 19616
rect 12289 19552 12305 19616
rect 12369 19552 12385 19616
rect 12449 19552 12465 19616
rect 12529 19552 12537 19616
rect 12217 18528 12537 19552
rect 12217 18464 12225 18528
rect 12289 18464 12305 18528
rect 12369 18464 12385 18528
rect 12449 18464 12465 18528
rect 12529 18464 12537 18528
rect 12217 17440 12537 18464
rect 12217 17376 12225 17440
rect 12289 17376 12305 17440
rect 12369 17376 12385 17440
rect 12449 17376 12465 17440
rect 12529 17376 12537 17440
rect 12217 16352 12537 17376
rect 12217 16288 12225 16352
rect 12289 16288 12305 16352
rect 12369 16288 12385 16352
rect 12449 16288 12465 16352
rect 12529 16288 12537 16352
rect 12217 15264 12537 16288
rect 12217 15200 12225 15264
rect 12289 15200 12305 15264
rect 12369 15200 12385 15264
rect 12449 15200 12465 15264
rect 12529 15200 12537 15264
rect 12217 14176 12537 15200
rect 12217 14112 12225 14176
rect 12289 14112 12305 14176
rect 12369 14112 12385 14176
rect 12449 14112 12465 14176
rect 12529 14112 12537 14176
rect 12217 13088 12537 14112
rect 12217 13024 12225 13088
rect 12289 13024 12305 13088
rect 12369 13024 12385 13088
rect 12449 13024 12465 13088
rect 12529 13024 12537 13088
rect 12217 12000 12537 13024
rect 12217 11936 12225 12000
rect 12289 11936 12305 12000
rect 12369 11936 12385 12000
rect 12449 11936 12465 12000
rect 12529 11936 12537 12000
rect 12217 10912 12537 11936
rect 12217 10848 12225 10912
rect 12289 10848 12305 10912
rect 12369 10848 12385 10912
rect 12449 10848 12465 10912
rect 12529 10848 12537 10912
rect 12217 9824 12537 10848
rect 12217 9760 12225 9824
rect 12289 9760 12305 9824
rect 12369 9760 12385 9824
rect 12449 9760 12465 9824
rect 12529 9760 12537 9824
rect 12217 8736 12537 9760
rect 12217 8672 12225 8736
rect 12289 8672 12305 8736
rect 12369 8672 12385 8736
rect 12449 8672 12465 8736
rect 12529 8672 12537 8736
rect 12217 7648 12537 8672
rect 12217 7584 12225 7648
rect 12289 7584 12305 7648
rect 12369 7584 12385 7648
rect 12449 7584 12465 7648
rect 12529 7584 12537 7648
rect 12217 6560 12537 7584
rect 12217 6496 12225 6560
rect 12289 6496 12305 6560
rect 12369 6496 12385 6560
rect 12449 6496 12465 6560
rect 12529 6496 12537 6560
rect 12217 5472 12537 6496
rect 12217 5408 12225 5472
rect 12289 5408 12305 5472
rect 12369 5408 12385 5472
rect 12449 5408 12465 5472
rect 12529 5408 12537 5472
rect 12217 4384 12537 5408
rect 12217 4320 12225 4384
rect 12289 4320 12305 4384
rect 12369 4320 12385 4384
rect 12449 4320 12465 4384
rect 12529 4320 12537 4384
rect 12217 3296 12537 4320
rect 12217 3232 12225 3296
rect 12289 3232 12305 3296
rect 12369 3232 12385 3296
rect 12449 3232 12465 3296
rect 12529 3232 12537 3296
rect 12217 2208 12537 3232
rect 12217 2144 12225 2208
rect 12289 2144 12305 2208
rect 12369 2144 12385 2208
rect 12449 2144 12465 2208
rect 12529 2144 12537 2208
rect 12217 2128 12537 2144
rect 15974 22336 16294 22352
rect 15974 22272 15982 22336
rect 16046 22272 16062 22336
rect 16126 22272 16142 22336
rect 16206 22272 16222 22336
rect 16286 22272 16294 22336
rect 15974 21248 16294 22272
rect 15974 21184 15982 21248
rect 16046 21184 16062 21248
rect 16126 21184 16142 21248
rect 16206 21184 16222 21248
rect 16286 21184 16294 21248
rect 15974 20160 16294 21184
rect 15974 20096 15982 20160
rect 16046 20096 16062 20160
rect 16126 20096 16142 20160
rect 16206 20096 16222 20160
rect 16286 20096 16294 20160
rect 15974 19072 16294 20096
rect 15974 19008 15982 19072
rect 16046 19008 16062 19072
rect 16126 19008 16142 19072
rect 16206 19008 16222 19072
rect 16286 19008 16294 19072
rect 15974 17984 16294 19008
rect 15974 17920 15982 17984
rect 16046 17920 16062 17984
rect 16126 17920 16142 17984
rect 16206 17920 16222 17984
rect 16286 17920 16294 17984
rect 15974 16896 16294 17920
rect 15974 16832 15982 16896
rect 16046 16832 16062 16896
rect 16126 16832 16142 16896
rect 16206 16832 16222 16896
rect 16286 16832 16294 16896
rect 15974 15808 16294 16832
rect 15974 15744 15982 15808
rect 16046 15744 16062 15808
rect 16126 15744 16142 15808
rect 16206 15744 16222 15808
rect 16286 15744 16294 15808
rect 15974 14720 16294 15744
rect 15974 14656 15982 14720
rect 16046 14656 16062 14720
rect 16126 14656 16142 14720
rect 16206 14656 16222 14720
rect 16286 14656 16294 14720
rect 15974 13632 16294 14656
rect 15974 13568 15982 13632
rect 16046 13568 16062 13632
rect 16126 13568 16142 13632
rect 16206 13568 16222 13632
rect 16286 13568 16294 13632
rect 15974 12544 16294 13568
rect 15974 12480 15982 12544
rect 16046 12480 16062 12544
rect 16126 12480 16142 12544
rect 16206 12480 16222 12544
rect 16286 12480 16294 12544
rect 15974 11456 16294 12480
rect 15974 11392 15982 11456
rect 16046 11392 16062 11456
rect 16126 11392 16142 11456
rect 16206 11392 16222 11456
rect 16286 11392 16294 11456
rect 15974 10368 16294 11392
rect 15974 10304 15982 10368
rect 16046 10304 16062 10368
rect 16126 10304 16142 10368
rect 16206 10304 16222 10368
rect 16286 10304 16294 10368
rect 15974 9280 16294 10304
rect 15974 9216 15982 9280
rect 16046 9216 16062 9280
rect 16126 9216 16142 9280
rect 16206 9216 16222 9280
rect 16286 9216 16294 9280
rect 15974 8192 16294 9216
rect 15974 8128 15982 8192
rect 16046 8128 16062 8192
rect 16126 8128 16142 8192
rect 16206 8128 16222 8192
rect 16286 8128 16294 8192
rect 15974 7104 16294 8128
rect 15974 7040 15982 7104
rect 16046 7040 16062 7104
rect 16126 7040 16142 7104
rect 16206 7040 16222 7104
rect 16286 7040 16294 7104
rect 15974 6016 16294 7040
rect 15974 5952 15982 6016
rect 16046 5952 16062 6016
rect 16126 5952 16142 6016
rect 16206 5952 16222 6016
rect 16286 5952 16294 6016
rect 15974 4928 16294 5952
rect 15974 4864 15982 4928
rect 16046 4864 16062 4928
rect 16126 4864 16142 4928
rect 16206 4864 16222 4928
rect 16286 4864 16294 4928
rect 15974 3840 16294 4864
rect 15974 3776 15982 3840
rect 16046 3776 16062 3840
rect 16126 3776 16142 3840
rect 16206 3776 16222 3840
rect 16286 3776 16294 3840
rect 15974 2752 16294 3776
rect 15974 2688 15982 2752
rect 16046 2688 16062 2752
rect 16126 2688 16142 2752
rect 16206 2688 16222 2752
rect 16286 2688 16294 2752
rect 15974 2128 16294 2688
rect 19732 21792 20052 22352
rect 19732 21728 19740 21792
rect 19804 21728 19820 21792
rect 19884 21728 19900 21792
rect 19964 21728 19980 21792
rect 20044 21728 20052 21792
rect 19732 20704 20052 21728
rect 19732 20640 19740 20704
rect 19804 20640 19820 20704
rect 19884 20640 19900 20704
rect 19964 20640 19980 20704
rect 20044 20640 20052 20704
rect 19732 19616 20052 20640
rect 19732 19552 19740 19616
rect 19804 19552 19820 19616
rect 19884 19552 19900 19616
rect 19964 19552 19980 19616
rect 20044 19552 20052 19616
rect 19732 18528 20052 19552
rect 19732 18464 19740 18528
rect 19804 18464 19820 18528
rect 19884 18464 19900 18528
rect 19964 18464 19980 18528
rect 20044 18464 20052 18528
rect 19732 17440 20052 18464
rect 19732 17376 19740 17440
rect 19804 17376 19820 17440
rect 19884 17376 19900 17440
rect 19964 17376 19980 17440
rect 20044 17376 20052 17440
rect 19732 16352 20052 17376
rect 19732 16288 19740 16352
rect 19804 16288 19820 16352
rect 19884 16288 19900 16352
rect 19964 16288 19980 16352
rect 20044 16288 20052 16352
rect 19732 15264 20052 16288
rect 19732 15200 19740 15264
rect 19804 15200 19820 15264
rect 19884 15200 19900 15264
rect 19964 15200 19980 15264
rect 20044 15200 20052 15264
rect 19732 14176 20052 15200
rect 19732 14112 19740 14176
rect 19804 14112 19820 14176
rect 19884 14112 19900 14176
rect 19964 14112 19980 14176
rect 20044 14112 20052 14176
rect 19732 13088 20052 14112
rect 22139 13156 22205 13157
rect 22139 13092 22140 13156
rect 22204 13092 22205 13156
rect 22139 13091 22205 13092
rect 19732 13024 19740 13088
rect 19804 13024 19820 13088
rect 19884 13024 19900 13088
rect 19964 13024 19980 13088
rect 20044 13024 20052 13088
rect 19732 12000 20052 13024
rect 22142 12885 22202 13091
rect 22139 12884 22205 12885
rect 22139 12820 22140 12884
rect 22204 12820 22205 12884
rect 22139 12819 22205 12820
rect 19732 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20052 12000
rect 19732 10912 20052 11936
rect 19732 10848 19740 10912
rect 19804 10848 19820 10912
rect 19884 10848 19900 10912
rect 19964 10848 19980 10912
rect 20044 10848 20052 10912
rect 19732 9824 20052 10848
rect 22139 10708 22205 10709
rect 22139 10644 22140 10708
rect 22204 10644 22205 10708
rect 22139 10643 22205 10644
rect 22142 10437 22202 10643
rect 22139 10436 22205 10437
rect 22139 10372 22140 10436
rect 22204 10372 22205 10436
rect 22139 10371 22205 10372
rect 19732 9760 19740 9824
rect 19804 9760 19820 9824
rect 19884 9760 19900 9824
rect 19964 9760 19980 9824
rect 20044 9760 20052 9824
rect 19732 8736 20052 9760
rect 19732 8672 19740 8736
rect 19804 8672 19820 8736
rect 19884 8672 19900 8736
rect 19964 8672 19980 8736
rect 20044 8672 20052 8736
rect 19732 7648 20052 8672
rect 19732 7584 19740 7648
rect 19804 7584 19820 7648
rect 19884 7584 19900 7648
rect 19964 7584 19980 7648
rect 20044 7584 20052 7648
rect 19732 6560 20052 7584
rect 19732 6496 19740 6560
rect 19804 6496 19820 6560
rect 19884 6496 19900 6560
rect 19964 6496 19980 6560
rect 20044 6496 20052 6560
rect 19732 5472 20052 6496
rect 19732 5408 19740 5472
rect 19804 5408 19820 5472
rect 19884 5408 19900 5472
rect 19964 5408 19980 5472
rect 20044 5408 20052 5472
rect 19732 4384 20052 5408
rect 19732 4320 19740 4384
rect 19804 4320 19820 4384
rect 19884 4320 19900 4384
rect 19964 4320 19980 4384
rect 20044 4320 20052 4384
rect 19732 3296 20052 4320
rect 19732 3232 19740 3296
rect 19804 3232 19820 3296
rect 19884 3232 19900 3296
rect 19964 3232 19980 3296
rect 20044 3232 20052 3296
rect 19732 2208 20052 3232
rect 19732 2144 19740 2208
rect 19804 2144 19820 2208
rect 19884 2144 19900 2208
rect 19964 2144 19980 2208
rect 20044 2144 20052 2208
rect 19732 2128 20052 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_78 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_81
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _38_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 774 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_136
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_184
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_190
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 866 592
use scs8hd_decap_12  FILLER_0_194
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 21436 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 21436 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_206
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_214
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_209
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_177
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 21436 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_82
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use scs8hd_conb_1  _24_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 21436 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_170
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 21436 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 774 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 866 592
use scs8hd_decap_6  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_181
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 21436 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 774 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 21436 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 21436 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_48
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_72
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_99
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_137
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _15_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 21436 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _16_
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_26
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_45
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_49
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 590 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 18216 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_189
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 21436 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_206
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_25
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_43
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_78
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 21436 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_47
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_82
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_133
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 21436 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 21436 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_78
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_82
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 21436 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 21436 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_8
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_50
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_137
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 21436 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_111
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 314 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_172
timestamp 1586364061
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_189
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 21436 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_91
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_95
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 1142 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_151
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 21436 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_13
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 21436 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_131
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_173
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_181
timestamp 1586364061
transform 1 0 17756 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_191
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_203
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 21436 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 21436 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_133
timestamp 1586364061
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_163
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 21436 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_38
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_120
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_137
timestamp 1586364061
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_164
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_22_172
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 21436 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_89
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_103
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 21436 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_216
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_90
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_182
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_194
timestamp 1586364061
transform 1 0 18952 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 21436 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_38
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 21436 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_216
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_33
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_39
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_41
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_104
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 21436 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 21436 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_216
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 21436 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_31
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 21436 0 1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_29_211
timestamp 1586364061
transform 1 0 20516 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_17
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_196
timestamp 1586364061
transform 1 0 19136 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 21436 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_129
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_133
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_137
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_191
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 21436 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_71
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 21436 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_20
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_28
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_42
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_34_40
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 7912 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_76
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_70
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_83
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_78
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_99
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_90
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_33_139
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_151
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 774 592
use scs8hd_decap_6  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_163
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_160
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_164
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_188
timestamp 1586364061
transform 1 0 18400 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_181
timestamp 1586364061
transform 1 0 17756 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_203
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 21436 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 21436 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_209
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_217
timestamp 1586364061
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_207
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_197
timestamp 1586364061
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 21436 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_210
timestamp 1586364061
transform 1 0 20424 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_94
timestamp 1586364061
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_118
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_156
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18492 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_180
timestamp 1586364061
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_192
timestamp 1586364061
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 21436 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_209
timestamp 1586364061
transform 1 0 20332 0 -1 22304
box -38 -48 774 592
<< labels >>
rlabel metal3 s 22066 416 22546 536 6 address[0]
port 0 nsew default input
rlabel metal2 s 754 24210 810 24690 6 address[1]
port 1 nsew default input
rlabel metal2 s 2226 24210 2282 24690 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 552 480 672 6 address[3]
port 3 nsew default input
rlabel metal3 s 22066 1368 22546 1488 6 address[4]
port 4 nsew default input
rlabel metal3 s 22066 2456 22546 2576 6 address[5]
port 5 nsew default input
rlabel metal3 s 22066 3408 22546 3528 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 1776 480 1896 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 3698 24210 3754 24690 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal2 s 5262 24210 5318 24690 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 22066 4496 22546 4616 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 22066 5448 22546 5568 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal2 s 3238 0 3294 480 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 22066 6536 22546 6656 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal2 s 6734 24210 6790 24690 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 5170 0 5226 480 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 7930 0 7986 480 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 8850 0 8906 480 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 8206 24210 8262 24690 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal2 s 9862 0 9918 480 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 0 7896 480 8016 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 22066 7624 22546 7744 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 22066 8576 22546 8696 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 12622 0 12678 480 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 22066 9664 22546 9784 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 22066 10616 22546 10736 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 22066 11704 22546 11824 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 22066 12792 22546 12912 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal3 s 22066 13744 22546 13864 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal3 s 22066 14832 22546 14952 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 9770 24210 9826 24690 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal3 s 22066 15784 22546 15904 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 11242 24210 11298 24690 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 12714 24210 12770 24690 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 14278 24210 14334 24690 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal3 s 22066 16872 22546 16992 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 15750 24210 15806 24690 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 17222 24210 17278 24690 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal3 s 22066 17824 22546 17944 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 63 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 64 nsew default input
rlabel metal2 s 18786 24210 18842 24690 6 left_bottom_grid_pin_12_
port 65 nsew default input
rlabel metal3 s 22066 20000 22546 20120 6 left_top_grid_pin_11_
port 66 nsew default input
rlabel metal2 s 20258 24210 20314 24690 6 left_top_grid_pin_13_
port 67 nsew default input
rlabel metal2 s 20166 0 20222 480 6 left_top_grid_pin_15_
port 68 nsew default input
rlabel metal2 s 17314 0 17370 480 6 left_top_grid_pin_1_
port 69 nsew default input
rlabel metal3 s 22066 18912 22546 19032 6 left_top_grid_pin_3_
port 70 nsew default input
rlabel metal2 s 18234 0 18290 480 6 left_top_grid_pin_5_
port 71 nsew default input
rlabel metal2 s 19246 0 19302 480 6 left_top_grid_pin_7_
port 72 nsew default input
rlabel metal3 s 0 21496 480 21616 6 left_top_grid_pin_9_
port 73 nsew default input
rlabel metal3 s 0 22720 480 22840 6 right_bottom_grid_pin_12_
port 74 nsew default input
rlabel metal2 s 21730 24210 21786 24690 6 right_top_grid_pin_11_
port 75 nsew default input
rlabel metal3 s 22066 22992 22546 23112 6 right_top_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 22066 24080 22546 24200 6 right_top_grid_pin_15_
port 77 nsew default input
rlabel metal2 s 21086 0 21142 480 6 right_top_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 22066 20952 22546 21072 6 right_top_grid_pin_3_
port 79 nsew default input
rlabel metal2 s 22006 0 22062 480 6 right_top_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 22066 22040 22546 22160 6 right_top_grid_pin_7_
port 81 nsew default input
rlabel metal3 s 0 23944 480 24064 6 right_top_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 4702 2128 5022 22352 6 vpwr
port 83 nsew default input
rlabel metal4 s 8459 2128 8779 22352 6 vgnd
port 84 nsew default input
<< end >>
