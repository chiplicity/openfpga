VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right
  CLASS BLOCK ;
  FOREIGN grid_io_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 193.760 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END address[3]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 2.400 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 12.280 80.000 12.880 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 36.760 80.000 37.360 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 61.920 80.000 62.520 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 87.080 80.000 87.680 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 112.240 80.000 112.840 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 136.720 80.000 137.320 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 161.880 80.000 162.480 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 187.040 80.000 187.640 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END left_width_0_height_0__pin_10_
  PIN left_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 2.400 144.120 ;
    END
  END left_width_0_height_0__pin_11_
  PIN left_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 2.400 156.360 ;
    END
  END left_width_0_height_0__pin_12_
  PIN left_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 2.400 168.600 ;
    END
  END left_width_0_height_0__pin_13_
  PIN left_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 2.400 181.520 ;
    END
  END left_width_0_height_0__pin_14_
  PIN left_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 2.400 193.760 ;
    END
  END left_width_0_height_0__pin_15_
  PIN left_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END left_width_0_height_0__pin_1_
  PIN left_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END left_width_0_height_0__pin_2_
  PIN left_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END left_width_0_height_0__pin_3_
  PIN left_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END left_width_0_height_0__pin_4_
  PIN left_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END left_width_0_height_0__pin_5_
  PIN left_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END left_width_0_height_0__pin_6_
  PIN left_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END left_width_0_height_0__pin_7_
  PIN left_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END left_width_0_height_0__pin_8_
  PIN left_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END left_width_0_height_0__pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 5.520 10.640 74.060 187.920 ;
      LAYER met2 ;
        RECT 6.530 2.680 73.510 193.645 ;
        RECT 7.090 2.400 19.590 2.680 ;
        RECT 20.430 2.400 32.930 2.680 ;
        RECT 33.770 2.400 46.270 2.680 ;
        RECT 47.110 2.400 59.610 2.680 ;
        RECT 60.450 2.400 72.950 2.680 ;
      LAYER met3 ;
        RECT 2.800 192.760 77.600 193.625 ;
        RECT 2.400 188.040 77.600 192.760 ;
        RECT 2.400 186.640 77.200 188.040 ;
        RECT 2.400 181.920 77.600 186.640 ;
        RECT 2.800 180.520 77.600 181.920 ;
        RECT 2.400 169.000 77.600 180.520 ;
        RECT 2.800 167.600 77.600 169.000 ;
        RECT 2.400 162.880 77.600 167.600 ;
        RECT 2.400 161.480 77.200 162.880 ;
        RECT 2.400 156.760 77.600 161.480 ;
        RECT 2.800 155.360 77.600 156.760 ;
        RECT 2.400 144.520 77.600 155.360 ;
        RECT 2.800 143.120 77.600 144.520 ;
        RECT 2.400 137.720 77.600 143.120 ;
        RECT 2.400 136.320 77.200 137.720 ;
        RECT 2.400 131.600 77.600 136.320 ;
        RECT 2.800 130.200 77.600 131.600 ;
        RECT 2.400 119.360 77.600 130.200 ;
        RECT 2.800 117.960 77.600 119.360 ;
        RECT 2.400 113.240 77.600 117.960 ;
        RECT 2.400 111.840 77.200 113.240 ;
        RECT 2.400 107.120 77.600 111.840 ;
        RECT 2.800 105.720 77.600 107.120 ;
        RECT 2.400 94.200 77.600 105.720 ;
        RECT 2.800 92.800 77.600 94.200 ;
        RECT 2.400 88.080 77.600 92.800 ;
        RECT 2.400 86.680 77.200 88.080 ;
        RECT 2.400 81.960 77.600 86.680 ;
        RECT 2.800 80.560 77.600 81.960 ;
        RECT 2.400 69.040 77.600 80.560 ;
        RECT 2.800 67.640 77.600 69.040 ;
        RECT 2.400 62.920 77.600 67.640 ;
        RECT 2.400 61.520 77.200 62.920 ;
        RECT 2.400 56.800 77.600 61.520 ;
        RECT 2.800 55.400 77.600 56.800 ;
        RECT 2.400 44.560 77.600 55.400 ;
        RECT 2.800 43.160 77.600 44.560 ;
        RECT 2.400 37.760 77.600 43.160 ;
        RECT 2.400 36.360 77.200 37.760 ;
        RECT 2.400 31.640 77.600 36.360 ;
        RECT 2.800 30.240 77.600 31.640 ;
        RECT 2.400 19.400 77.600 30.240 ;
        RECT 2.800 18.000 77.600 19.400 ;
        RECT 2.400 13.280 77.600 18.000 ;
        RECT 2.400 11.880 77.200 13.280 ;
        RECT 2.400 7.160 77.600 11.880 ;
        RECT 2.800 6.295 77.600 7.160 ;
      LAYER met4 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END grid_io_right
END LIBRARY

