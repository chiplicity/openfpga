magic
tech sky130A
magscale 1 2
timestamp 1605123239
<< locali >>
rect 14933 12087 14967 12257
rect 3709 11679 3743 11849
rect 12633 10999 12667 11169
rect 8861 3519 8895 3689
rect 13093 3519 13127 3689
rect 6101 2839 6135 3077
rect 4997 2295 5031 2397
rect 11805 2295 11839 2465
rect 12633 2363 12667 2533
<< viali >>
rect 9965 25449 9999 25483
rect 11069 25449 11103 25483
rect 2053 25381 2087 25415
rect 1777 25313 1811 25347
rect 4077 25313 4111 25347
rect 5181 25313 5215 25347
rect 7573 25313 7607 25347
rect 7665 25313 7699 25347
rect 9781 25313 9815 25347
rect 10885 25313 10919 25347
rect 12633 25313 12667 25347
rect 13737 25313 13771 25347
rect 15485 25313 15519 25347
rect 7757 25245 7791 25279
rect 1685 25177 1719 25211
rect 7205 25177 7239 25211
rect 11437 25177 11471 25211
rect 13921 25177 13955 25211
rect 4261 25109 4295 25143
rect 5365 25109 5399 25143
rect 5733 25109 5767 25143
rect 6745 25109 6779 25143
rect 12817 25109 12851 25143
rect 13553 25109 13587 25143
rect 15669 25109 15703 25143
rect 2421 24905 2455 24939
rect 7021 24905 7055 24939
rect 10609 24905 10643 24939
rect 12633 24905 12667 24939
rect 13369 24905 13403 24939
rect 13737 24905 13771 24939
rect 16037 24905 16071 24939
rect 8033 24837 8067 24871
rect 1869 24769 1903 24803
rect 4721 24769 4755 24803
rect 5641 24769 5675 24803
rect 5825 24769 5859 24803
rect 7573 24769 7607 24803
rect 11253 24769 11287 24803
rect 1593 24701 1627 24735
rect 2881 24701 2915 24735
rect 6653 24701 6687 24735
rect 8585 24701 8619 24735
rect 9137 24701 9171 24735
rect 9689 24701 9723 24735
rect 10241 24701 10275 24735
rect 11069 24701 11103 24735
rect 12449 24701 12483 24735
rect 13001 24701 13035 24735
rect 13553 24701 13587 24735
rect 15485 24701 15519 24735
rect 16865 24701 16899 24735
rect 3157 24633 3191 24667
rect 4169 24633 4203 24667
rect 5089 24633 5123 24667
rect 7481 24633 7515 24667
rect 15393 24633 15427 24667
rect 3709 24565 3743 24599
rect 5181 24565 5215 24599
rect 5549 24565 5583 24599
rect 6285 24565 6319 24599
rect 7389 24565 7423 24599
rect 8401 24565 8435 24599
rect 8769 24565 8803 24599
rect 9873 24565 9907 24599
rect 11897 24565 11931 24599
rect 14105 24565 14139 24599
rect 15669 24565 15703 24599
rect 17049 24565 17083 24599
rect 17509 24565 17543 24599
rect 12265 24361 12299 24395
rect 15485 24361 15519 24395
rect 17693 24361 17727 24395
rect 18797 24361 18831 24395
rect 19901 24361 19935 24395
rect 21097 24361 21131 24395
rect 22201 24361 22235 24395
rect 4905 24293 4939 24327
rect 1685 24225 1719 24259
rect 1961 24225 1995 24259
rect 6837 24225 6871 24259
rect 7196 24225 7230 24259
rect 10129 24225 10163 24259
rect 12081 24225 12115 24259
rect 13553 24225 13587 24259
rect 13829 24225 13863 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 18613 24225 18647 24259
rect 19717 24225 19751 24259
rect 20913 24225 20947 24259
rect 22017 24225 22051 24259
rect 2973 24157 3007 24191
rect 4997 24157 5031 24191
rect 5089 24157 5123 24191
rect 6929 24157 6963 24191
rect 9873 24157 9907 24191
rect 4537 24089 4571 24123
rect 16589 24089 16623 24123
rect 2513 24021 2547 24055
rect 4353 24021 4387 24055
rect 5641 24021 5675 24055
rect 8309 24021 8343 24055
rect 8585 24021 8619 24055
rect 9137 24021 9171 24055
rect 9505 24021 9539 24055
rect 11253 24021 11287 24055
rect 11621 24021 11655 24055
rect 12725 24021 12759 24055
rect 14289 24021 14323 24055
rect 2421 23817 2455 23851
rect 2881 23817 2915 23851
rect 4077 23817 4111 23851
rect 5917 23817 5951 23851
rect 6285 23817 6319 23851
rect 6653 23817 6687 23851
rect 12449 23817 12483 23851
rect 15669 23817 15703 23851
rect 16405 23817 16439 23851
rect 18245 23817 18279 23851
rect 19349 23817 19383 23851
rect 20453 23817 20487 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 23857 23817 23891 23851
rect 4445 23749 4479 23783
rect 3525 23681 3559 23715
rect 6837 23681 6871 23715
rect 12909 23681 12943 23715
rect 13093 23681 13127 23715
rect 14013 23681 14047 23715
rect 20913 23681 20947 23715
rect 1593 23613 1627 23647
rect 3341 23613 3375 23647
rect 3433 23613 3467 23647
rect 4537 23613 4571 23647
rect 7757 23613 7791 23647
rect 7849 23613 7883 23647
rect 8105 23613 8139 23647
rect 10149 23613 10183 23647
rect 11897 23613 11931 23647
rect 16221 23613 16255 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 21373 23613 21407 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 1869 23545 1903 23579
rect 4782 23545 4816 23579
rect 7389 23545 7423 23579
rect 9597 23545 9631 23579
rect 10394 23545 10428 23579
rect 13461 23545 13495 23579
rect 14258 23545 14292 23579
rect 18981 23545 19015 23579
rect 2973 23477 3007 23511
rect 9229 23477 9263 23511
rect 9965 23477 9999 23511
rect 11529 23477 11563 23511
rect 12265 23477 12299 23511
rect 12817 23477 12851 23511
rect 13921 23477 13955 23511
rect 15393 23477 15427 23511
rect 16037 23477 16071 23511
rect 16773 23477 16807 23511
rect 17509 23477 17543 23511
rect 20085 23477 20119 23511
rect 22017 23477 22051 23511
rect 3433 23273 3467 23307
rect 8677 23273 8711 23307
rect 9137 23273 9171 23307
rect 10793 23273 10827 23307
rect 12633 23273 12667 23307
rect 13461 23273 13495 23307
rect 14473 23273 14507 23307
rect 19349 23273 19383 23307
rect 2053 23205 2087 23239
rect 11520 23205 11554 23239
rect 13829 23205 13863 23239
rect 16589 23205 16623 23239
rect 22661 23205 22695 23239
rect 1777 23137 1811 23171
rect 4344 23137 4378 23171
rect 7297 23137 7331 23171
rect 7553 23137 7587 23171
rect 10057 23137 10091 23171
rect 11253 23137 11287 23171
rect 15301 23137 15335 23171
rect 16313 23137 16347 23171
rect 17877 23137 17911 23171
rect 18153 23137 18187 23171
rect 19165 23137 19199 23171
rect 22385 23137 22419 23171
rect 4077 23069 4111 23103
rect 6285 23069 6319 23103
rect 9505 23069 9539 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 13921 23069 13955 23103
rect 14105 23069 14139 23103
rect 1685 22933 1719 22967
rect 2513 22933 2547 22967
rect 3065 22933 3099 22967
rect 3893 22933 3927 22967
rect 5457 22933 5491 22967
rect 9689 22933 9723 22967
rect 12909 22933 12943 22967
rect 13277 22933 13311 22967
rect 20269 22933 20303 22967
rect 21373 22933 21407 22967
rect 1685 22729 1719 22763
rect 2145 22729 2179 22763
rect 5641 22729 5675 22763
rect 6009 22729 6043 22763
rect 6653 22729 6687 22763
rect 7389 22729 7423 22763
rect 7849 22729 7883 22763
rect 8861 22729 8895 22763
rect 9321 22729 9355 22763
rect 10793 22729 10827 22763
rect 11897 22729 11931 22763
rect 12173 22729 12207 22763
rect 13461 22729 13495 22763
rect 14933 22729 14967 22763
rect 15301 22729 15335 22763
rect 19165 22729 19199 22763
rect 22385 22729 22419 22763
rect 10241 22661 10275 22695
rect 12633 22661 12667 22695
rect 2605 22593 2639 22627
rect 2789 22593 2823 22627
rect 3801 22593 3835 22627
rect 6837 22593 6871 22627
rect 7757 22593 7791 22627
rect 8309 22593 8343 22627
rect 8493 22593 8527 22627
rect 9689 22593 9723 22627
rect 10701 22593 10735 22627
rect 11253 22593 11287 22627
rect 11345 22593 11379 22627
rect 16037 22593 16071 22627
rect 2053 22525 2087 22559
rect 3893 22525 3927 22559
rect 4160 22525 4194 22559
rect 9413 22525 9447 22559
rect 12449 22525 12483 22559
rect 13553 22525 13587 22559
rect 13820 22525 13854 22559
rect 15761 22525 15795 22559
rect 16497 22525 16531 22559
rect 2513 22457 2547 22491
rect 3157 22457 3191 22491
rect 13093 22457 13127 22491
rect 18245 22457 18279 22491
rect 5273 22389 5307 22423
rect 8217 22389 8251 22423
rect 11161 22389 11195 22423
rect 16865 22389 16899 22423
rect 4353 22185 4387 22219
rect 9137 22185 9171 22219
rect 14657 22185 14691 22219
rect 2789 22117 2823 22151
rect 5080 22117 5114 22151
rect 7021 22117 7055 22151
rect 8401 22117 8435 22151
rect 14013 22117 14047 22151
rect 10057 22049 10091 22083
rect 11713 22049 11747 22083
rect 12541 22049 12575 22083
rect 13553 22049 13587 22083
rect 15301 22049 15335 22083
rect 15568 22049 15602 22083
rect 2881 21981 2915 22015
rect 3065 21981 3099 22015
rect 3525 21981 3559 22015
rect 4721 21981 4755 22015
rect 4813 21981 4847 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 11805 21981 11839 22015
rect 11897 21981 11931 22015
rect 13185 21981 13219 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 1685 21913 1719 21947
rect 2421 21913 2455 21947
rect 3801 21913 3835 21947
rect 7849 21913 7883 21947
rect 9689 21913 9723 21947
rect 11253 21913 11287 21947
rect 1961 21845 1995 21879
rect 6193 21845 6227 21879
rect 6561 21845 6595 21879
rect 6837 21845 6871 21879
rect 7573 21845 7607 21879
rect 8033 21845 8067 21879
rect 9505 21845 9539 21879
rect 10885 21845 10919 21879
rect 11345 21845 11379 21879
rect 13645 21845 13679 21879
rect 16681 21845 16715 21879
rect 1409 21641 1443 21675
rect 2513 21641 2547 21675
rect 3249 21641 3283 21675
rect 4905 21641 4939 21675
rect 8033 21641 8067 21675
rect 9505 21641 9539 21675
rect 10333 21641 10367 21675
rect 11897 21641 11931 21675
rect 12633 21641 12667 21675
rect 13277 21641 13311 21675
rect 15945 21641 15979 21675
rect 3709 21573 3743 21607
rect 10241 21573 10275 21607
rect 15117 21573 15151 21607
rect 1961 21505 1995 21539
rect 4261 21505 4295 21539
rect 4445 21505 4479 21539
rect 5549 21505 5583 21539
rect 7021 21505 7055 21539
rect 10977 21505 11011 21539
rect 13737 21505 13771 21539
rect 15485 21505 15519 21539
rect 16589 21505 16623 21539
rect 16957 21505 16991 21539
rect 1777 21437 1811 21471
rect 4169 21437 4203 21471
rect 5365 21437 5399 21471
rect 6101 21437 6135 21471
rect 6653 21437 6687 21471
rect 6837 21437 6871 21471
rect 8125 21437 8159 21471
rect 8392 21437 8426 21471
rect 10793 21437 10827 21471
rect 12081 21437 12115 21471
rect 12449 21437 12483 21471
rect 7665 21369 7699 21403
rect 13982 21369 14016 21403
rect 1869 21301 1903 21335
rect 2881 21301 2915 21335
rect 3801 21301 3835 21335
rect 5273 21301 5307 21335
rect 9873 21301 9907 21335
rect 10701 21301 10735 21335
rect 11437 21301 11471 21335
rect 11805 21301 11839 21335
rect 13645 21301 13679 21335
rect 15761 21301 15795 21335
rect 16313 21301 16347 21335
rect 16405 21301 16439 21335
rect 1409 21097 1443 21131
rect 3893 21097 3927 21131
rect 4905 21097 4939 21131
rect 5457 21097 5491 21131
rect 8401 21097 8435 21131
rect 8769 21097 8803 21131
rect 9137 21097 9171 21131
rect 11069 21097 11103 21131
rect 11713 21097 11747 21131
rect 12081 21097 12115 21131
rect 13645 21097 13679 21131
rect 14657 21097 14691 21131
rect 15025 21097 15059 21131
rect 4353 21029 4387 21063
rect 5917 21029 5951 21063
rect 7266 21029 7300 21063
rect 9934 21029 9968 21063
rect 11437 21029 11471 21063
rect 13553 21029 13587 21063
rect 1777 20961 1811 20995
rect 4077 20961 4111 20995
rect 5825 20961 5859 20995
rect 6929 20961 6963 20995
rect 9413 20961 9447 20995
rect 9689 20961 9723 20995
rect 12449 20961 12483 20995
rect 14013 20961 14047 20995
rect 1869 20893 1903 20927
rect 1961 20893 1995 20927
rect 6101 20893 6135 20927
rect 7021 20893 7055 20927
rect 12541 20893 12575 20927
rect 12633 20893 12667 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 15301 20893 15335 20927
rect 16313 20893 16347 20927
rect 2789 20825 2823 20859
rect 9229 20825 9263 20859
rect 2513 20757 2547 20791
rect 3525 20757 3559 20791
rect 5273 20757 5307 20791
rect 6561 20757 6595 20791
rect 13185 20757 13219 20791
rect 15945 20757 15979 20791
rect 6285 20553 6319 20587
rect 6653 20553 6687 20587
rect 8217 20553 8251 20587
rect 9229 20553 9263 20587
rect 9781 20553 9815 20587
rect 12173 20553 12207 20587
rect 13829 20553 13863 20587
rect 14105 20553 14139 20587
rect 14565 20553 14599 20587
rect 15209 20553 15243 20587
rect 16037 20553 16071 20587
rect 8585 20485 8619 20519
rect 15485 20485 15519 20519
rect 2697 20417 2731 20451
rect 4169 20417 4203 20451
rect 4721 20417 4755 20451
rect 5825 20417 5859 20451
rect 12449 20417 12483 20451
rect 14657 20417 14691 20451
rect 4077 20349 4111 20383
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 7104 20349 7138 20383
rect 9045 20349 9079 20383
rect 10149 20349 10183 20383
rect 15853 20349 15887 20383
rect 16405 20349 16439 20383
rect 2513 20281 2547 20315
rect 3525 20281 3559 20315
rect 5549 20281 5583 20315
rect 10416 20281 10450 20315
rect 12716 20281 12750 20315
rect 1593 20213 1627 20247
rect 2053 20213 2087 20247
rect 2421 20213 2455 20247
rect 3065 20213 3099 20247
rect 3617 20213 3651 20247
rect 3985 20213 4019 20247
rect 4997 20213 5031 20247
rect 5181 20213 5215 20247
rect 8953 20213 8987 20247
rect 11529 20213 11563 20247
rect 2053 20009 2087 20043
rect 2881 20009 2915 20043
rect 3709 20009 3743 20043
rect 5825 20009 5859 20043
rect 6745 20009 6779 20043
rect 7205 20009 7239 20043
rect 7941 20009 7975 20043
rect 9689 20009 9723 20043
rect 10793 20009 10827 20043
rect 13461 20009 13495 20043
rect 13829 20009 13863 20043
rect 14933 20009 14967 20043
rect 16681 20009 16715 20043
rect 4322 19941 4356 19975
rect 6101 19941 6135 19975
rect 6561 19941 6595 19975
rect 10149 19941 10183 19975
rect 13277 19941 13311 19975
rect 2789 19873 2823 19907
rect 7113 19873 7147 19907
rect 8309 19873 8343 19907
rect 8861 19873 8895 19907
rect 10057 19873 10091 19907
rect 11253 19873 11287 19907
rect 11509 19873 11543 19907
rect 15301 19873 15335 19907
rect 15557 19873 15591 19907
rect 3065 19805 3099 19839
rect 4077 19805 4111 19839
rect 7297 19805 7331 19839
rect 10333 19805 10367 19839
rect 13921 19805 13955 19839
rect 14013 19805 14047 19839
rect 8493 19737 8527 19771
rect 12633 19737 12667 19771
rect 13001 19737 13035 19771
rect 1593 19669 1627 19703
rect 2421 19669 2455 19703
rect 5457 19669 5491 19703
rect 9413 19669 9447 19703
rect 11161 19669 11195 19703
rect 14473 19669 14507 19703
rect 3801 19465 3835 19499
rect 6285 19465 6319 19499
rect 7389 19465 7423 19499
rect 10977 19465 11011 19499
rect 12449 19465 12483 19499
rect 16681 19465 16715 19499
rect 13921 19397 13955 19431
rect 3341 19329 3375 19363
rect 6837 19329 6871 19363
rect 8401 19329 8435 19363
rect 9965 19329 9999 19363
rect 13093 19329 13127 19363
rect 14473 19329 14507 19363
rect 14657 19329 14691 19363
rect 15853 19329 15887 19363
rect 1409 19261 1443 19295
rect 3065 19261 3099 19295
rect 4261 19261 4295 19295
rect 6653 19261 6687 19295
rect 7665 19261 7699 19295
rect 8309 19261 8343 19295
rect 8953 19261 8987 19295
rect 10425 19261 10459 19295
rect 11069 19261 11103 19295
rect 12909 19261 12943 19295
rect 13553 19261 13587 19295
rect 15577 19261 15611 19295
rect 16313 19261 16347 19295
rect 1685 19193 1719 19227
rect 2513 19193 2547 19227
rect 4528 19193 4562 19227
rect 9873 19193 9907 19227
rect 11345 19193 11379 19227
rect 14381 19193 14415 19227
rect 15025 19193 15059 19227
rect 2697 19125 2731 19159
rect 3157 19125 3191 19159
rect 4077 19125 4111 19159
rect 5641 19125 5675 19159
rect 7849 19125 7883 19159
rect 8217 19125 8251 19159
rect 9229 19125 9263 19159
rect 9413 19125 9447 19159
rect 9781 19125 9815 19159
rect 11897 19125 11931 19159
rect 12173 19125 12207 19159
rect 12817 19125 12851 19159
rect 14013 19125 14047 19159
rect 15393 19125 15427 19159
rect 2789 18921 2823 18955
rect 3893 18921 3927 18955
rect 4261 18921 4295 18955
rect 4721 18921 4755 18955
rect 5641 18921 5675 18955
rect 7849 18921 7883 18955
rect 8493 18921 8527 18955
rect 9689 18921 9723 18955
rect 10149 18921 10183 18955
rect 12909 18921 12943 18955
rect 13461 18921 13495 18955
rect 13645 18921 13679 18955
rect 14105 18921 14139 18955
rect 15301 18921 15335 18955
rect 2329 18853 2363 18887
rect 4629 18785 4663 18819
rect 6081 18785 6115 18819
rect 8401 18785 8435 18819
rect 10957 18785 10991 18819
rect 14013 18785 14047 18819
rect 15669 18785 15703 18819
rect 2881 18717 2915 18751
rect 3065 18717 3099 18751
rect 4813 18717 4847 18751
rect 5825 18717 5859 18751
rect 8585 18717 8619 18751
rect 10701 18717 10735 18751
rect 12541 18717 12575 18751
rect 14197 18717 14231 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 2421 18649 2455 18683
rect 14749 18649 14783 18683
rect 1685 18581 1719 18615
rect 3433 18581 3467 18615
rect 5273 18581 5307 18615
rect 7205 18581 7239 18615
rect 7573 18581 7607 18615
rect 8033 18581 8067 18615
rect 9045 18581 9079 18615
rect 9413 18581 9447 18615
rect 10609 18581 10643 18615
rect 12081 18581 12115 18615
rect 1409 18377 1443 18411
rect 2513 18377 2547 18411
rect 4445 18377 4479 18411
rect 4813 18377 4847 18411
rect 5089 18377 5123 18411
rect 5457 18377 5491 18411
rect 7297 18377 7331 18411
rect 10333 18377 10367 18411
rect 10793 18377 10827 18411
rect 12173 18377 12207 18411
rect 13737 18377 13771 18411
rect 15761 18377 15795 18411
rect 5825 18309 5859 18343
rect 8309 18309 8343 18343
rect 8677 18309 8711 18343
rect 8861 18309 8895 18343
rect 9873 18309 9907 18343
rect 11805 18309 11839 18343
rect 12449 18309 12483 18343
rect 2053 18241 2087 18275
rect 3065 18241 3099 18275
rect 6653 18241 6687 18275
rect 7757 18241 7791 18275
rect 7849 18241 7883 18275
rect 9321 18241 9355 18275
rect 9505 18241 9539 18275
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 14289 18241 14323 18275
rect 5273 18173 5307 18207
rect 7205 18173 7239 18207
rect 10701 18173 10735 18207
rect 14381 18173 14415 18207
rect 14648 18173 14682 18207
rect 16773 18173 16807 18207
rect 1777 18105 1811 18139
rect 2973 18105 3007 18139
rect 3310 18105 3344 18139
rect 6193 18105 6227 18139
rect 16037 18105 16071 18139
rect 1869 18037 1903 18071
rect 7665 18037 7699 18071
rect 9229 18037 9263 18071
rect 11161 18037 11195 18071
rect 12817 18037 12851 18071
rect 16497 18037 16531 18071
rect 2421 17833 2455 17867
rect 3433 17833 3467 17867
rect 3801 17833 3835 17867
rect 4261 17833 4295 17867
rect 4445 17833 4479 17867
rect 5917 17833 5951 17867
rect 8769 17833 8803 17867
rect 11069 17833 11103 17867
rect 13737 17833 13771 17867
rect 14013 17833 14047 17867
rect 14197 17833 14231 17867
rect 14657 17833 14691 17867
rect 16681 17833 16715 17867
rect 2789 17765 2823 17799
rect 9934 17765 9968 17799
rect 2881 17697 2915 17731
rect 4813 17697 4847 17731
rect 5457 17697 5491 17731
rect 6009 17697 6043 17731
rect 7656 17697 7690 17731
rect 9689 17697 9723 17731
rect 12245 17697 12279 17731
rect 15301 17697 15335 17731
rect 15568 17697 15602 17731
rect 2973 17629 3007 17663
rect 4905 17629 4939 17663
rect 5089 17629 5123 17663
rect 6193 17629 6227 17663
rect 6929 17629 6963 17663
rect 7389 17629 7423 17663
rect 11989 17629 12023 17663
rect 1685 17561 1719 17595
rect 2053 17493 2087 17527
rect 7205 17493 7239 17527
rect 9137 17493 9171 17527
rect 9413 17493 9447 17527
rect 11345 17493 11379 17527
rect 11897 17493 11931 17527
rect 13369 17493 13403 17527
rect 1593 17289 1627 17323
rect 3525 17289 3559 17323
rect 3801 17289 3835 17323
rect 4261 17289 4295 17323
rect 4721 17289 4755 17323
rect 5733 17289 5767 17323
rect 7941 17289 7975 17323
rect 8125 17289 8159 17323
rect 9873 17289 9907 17323
rect 7021 17221 7055 17255
rect 9689 17221 9723 17255
rect 13921 17221 13955 17255
rect 2145 17153 2179 17187
rect 5273 17153 5307 17187
rect 8677 17153 8711 17187
rect 9413 17153 9447 17187
rect 10517 17153 10551 17187
rect 13001 17153 13035 17187
rect 13461 17153 13495 17187
rect 16865 17153 16899 17187
rect 2401 17085 2435 17119
rect 6837 17085 6871 17119
rect 8493 17085 8527 17119
rect 8585 17085 8619 17119
rect 12265 17085 12299 17119
rect 12817 17085 12851 17119
rect 14105 17085 14139 17119
rect 14361 17085 14395 17119
rect 16773 17085 16807 17119
rect 2053 17017 2087 17051
rect 5181 17017 5215 17051
rect 6561 17017 6595 17051
rect 10241 17017 10275 17051
rect 10885 17017 10919 17051
rect 11805 17017 11839 17051
rect 12909 17017 12943 17051
rect 16221 17017 16255 17051
rect 4629 16949 4663 16983
rect 5089 16949 5123 16983
rect 6101 16949 6135 16983
rect 7389 16949 7423 16983
rect 10333 16949 10367 16983
rect 11253 16949 11287 16983
rect 12449 16949 12483 16983
rect 15485 16949 15519 16983
rect 15853 16949 15887 16983
rect 16313 16949 16347 16983
rect 16681 16949 16715 16983
rect 1593 16745 1627 16779
rect 2237 16745 2271 16779
rect 2421 16745 2455 16779
rect 3433 16745 3467 16779
rect 4077 16745 4111 16779
rect 4813 16745 4847 16779
rect 5089 16745 5123 16779
rect 6193 16745 6227 16779
rect 6561 16745 6595 16779
rect 6929 16745 6963 16779
rect 7757 16745 7791 16779
rect 9137 16745 9171 16779
rect 9873 16745 9907 16779
rect 10885 16745 10919 16779
rect 11253 16745 11287 16779
rect 12081 16745 12115 16779
rect 12265 16745 12299 16779
rect 12725 16745 12759 16779
rect 15025 16745 15059 16779
rect 15301 16745 15335 16779
rect 16681 16745 16715 16779
rect 2789 16677 2823 16711
rect 3893 16677 3927 16711
rect 5549 16677 5583 16711
rect 8861 16677 8895 16711
rect 12633 16677 12667 16711
rect 15669 16677 15703 16711
rect 17049 16677 17083 16711
rect 2881 16609 2915 16643
rect 5457 16609 5491 16643
rect 10241 16609 10275 16643
rect 16313 16609 16347 16643
rect 3065 16541 3099 16575
rect 5641 16541 5675 16575
rect 7849 16541 7883 16575
rect 8033 16541 8067 16575
rect 10333 16541 10367 16575
rect 10517 16541 10551 16575
rect 12817 16541 12851 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 7389 16473 7423 16507
rect 7297 16405 7331 16439
rect 8401 16405 8435 16439
rect 13829 16405 13863 16439
rect 14197 16405 14231 16439
rect 2973 16201 3007 16235
rect 4721 16201 4755 16235
rect 5181 16201 5215 16235
rect 8309 16201 8343 16235
rect 8585 16201 8619 16235
rect 9229 16201 9263 16235
rect 9781 16201 9815 16235
rect 10885 16201 10919 16235
rect 11805 16201 11839 16235
rect 12265 16201 12299 16235
rect 15209 16201 15243 16235
rect 16037 16201 16071 16235
rect 17049 16201 17083 16235
rect 9689 16133 9723 16167
rect 15577 16133 15611 16167
rect 3341 16065 3375 16099
rect 4169 16065 4203 16099
rect 5825 16065 5859 16099
rect 7481 16065 7515 16099
rect 10333 16065 10367 16099
rect 11345 16065 11379 16099
rect 12633 16065 12667 16099
rect 13829 16065 13863 16099
rect 16589 16065 16623 16099
rect 1593 15997 1627 16031
rect 3893 15997 3927 16031
rect 5641 15997 5675 16031
rect 6193 15997 6227 16031
rect 6561 15997 6595 16031
rect 7297 15997 7331 16031
rect 8401 15997 8435 16031
rect 10241 15997 10275 16031
rect 12449 15997 12483 16031
rect 13185 15997 13219 16031
rect 1860 15929 1894 15963
rect 7849 15929 7883 15963
rect 10149 15929 10183 15963
rect 11161 15929 11195 15963
rect 14074 15929 14108 15963
rect 15945 15929 15979 15963
rect 3709 15861 3743 15895
rect 5089 15861 5123 15895
rect 5549 15861 5583 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 13645 15861 13679 15895
rect 16405 15861 16439 15895
rect 16497 15861 16531 15895
rect 17509 15861 17543 15895
rect 17785 15861 17819 15895
rect 1685 15657 1719 15691
rect 2237 15657 2271 15691
rect 2421 15657 2455 15691
rect 2789 15657 2823 15691
rect 4905 15657 4939 15691
rect 6101 15657 6135 15691
rect 6653 15657 6687 15691
rect 9505 15657 9539 15691
rect 10057 15657 10091 15691
rect 12357 15657 12391 15691
rect 14197 15657 14231 15691
rect 15761 15657 15795 15691
rect 16865 15657 16899 15691
rect 4629 15589 4663 15623
rect 8493 15589 8527 15623
rect 9045 15589 9079 15623
rect 9965 15589 9999 15623
rect 16681 15589 16715 15623
rect 17325 15589 17359 15623
rect 21189 15589 21223 15623
rect 2881 15521 2915 15555
rect 3433 15521 3467 15555
rect 5457 15521 5491 15555
rect 5549 15521 5583 15555
rect 7021 15521 7055 15555
rect 8033 15521 8067 15555
rect 8217 15521 8251 15555
rect 10425 15521 10459 15555
rect 13073 15521 13107 15555
rect 14473 15521 14507 15555
rect 15669 15521 15703 15555
rect 17233 15521 17267 15555
rect 20913 15521 20947 15555
rect 2973 15453 3007 15487
rect 5733 15453 5767 15487
rect 6561 15453 6595 15487
rect 7113 15453 7147 15487
rect 7297 15453 7331 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 11805 15453 11839 15487
rect 12817 15453 12851 15487
rect 15853 15453 15887 15487
rect 17417 15453 17451 15487
rect 3893 15385 3927 15419
rect 15301 15385 15335 15419
rect 5089 15317 5123 15351
rect 7757 15317 7791 15351
rect 11069 15317 11103 15351
rect 12725 15317 12759 15351
rect 15117 15317 15151 15351
rect 16405 15317 16439 15351
rect 18153 15317 18187 15351
rect 3249 15113 3283 15147
rect 3525 15113 3559 15147
rect 5917 15113 5951 15147
rect 9505 15113 9539 15147
rect 10057 15113 10091 15147
rect 11069 15113 11103 15147
rect 12449 15113 12483 15147
rect 13829 15113 13863 15147
rect 17785 15113 17819 15147
rect 18061 15113 18095 15147
rect 20913 15113 20947 15147
rect 5549 15045 5583 15079
rect 6193 15045 6227 15079
rect 13461 15045 13495 15079
rect 1869 14977 1903 15011
rect 10701 14977 10735 15011
rect 12265 14977 12299 15011
rect 13001 14977 13035 15011
rect 14565 14977 14599 15011
rect 18613 14977 18647 15011
rect 4169 14909 4203 14943
rect 6837 14909 6871 14943
rect 14381 14909 14415 14943
rect 14473 14909 14507 14943
rect 15761 14909 15795 14943
rect 1777 14841 1811 14875
rect 2114 14841 2148 14875
rect 4077 14841 4111 14875
rect 4436 14841 4470 14875
rect 7082 14841 7116 14875
rect 9229 14841 9263 14875
rect 10425 14841 10459 14875
rect 11897 14841 11931 14875
rect 12817 14841 12851 14875
rect 16028 14841 16062 14875
rect 17417 14841 17451 14875
rect 18429 14841 18463 14875
rect 6561 14773 6595 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 9873 14773 9907 14807
rect 10517 14773 10551 14807
rect 11529 14773 11563 14807
rect 12909 14773 12943 14807
rect 14013 14773 14047 14807
rect 15393 14773 15427 14807
rect 17141 14773 17175 14807
rect 18521 14773 18555 14807
rect 2237 14569 2271 14603
rect 2421 14569 2455 14603
rect 2789 14569 2823 14603
rect 4997 14569 5031 14603
rect 9045 14569 9079 14603
rect 10609 14569 10643 14603
rect 12541 14569 12575 14603
rect 15577 14569 15611 14603
rect 6929 14501 6963 14535
rect 7656 14501 7690 14535
rect 11038 14501 11072 14535
rect 16764 14501 16798 14535
rect 2881 14433 2915 14467
rect 3801 14433 3835 14467
rect 4077 14433 4111 14467
rect 4629 14433 4663 14467
rect 5181 14433 5215 14467
rect 5448 14433 5482 14467
rect 7389 14433 7423 14467
rect 9505 14433 9539 14467
rect 13257 14433 13291 14467
rect 3065 14365 3099 14399
rect 9689 14365 9723 14399
rect 10793 14365 10827 14399
rect 13001 14365 13035 14399
rect 15117 14365 15151 14399
rect 16497 14365 16531 14399
rect 4261 14297 4295 14331
rect 10241 14297 10275 14331
rect 12173 14297 12207 14331
rect 15853 14297 15887 14331
rect 1593 14229 1627 14263
rect 3433 14229 3467 14263
rect 6561 14229 6595 14263
rect 7205 14229 7239 14263
rect 8769 14229 8803 14263
rect 12817 14229 12851 14263
rect 14381 14229 14415 14263
rect 16313 14229 16347 14263
rect 17877 14229 17911 14263
rect 18153 14229 18187 14263
rect 2421 14025 2455 14059
rect 5457 14025 5491 14059
rect 5733 14025 5767 14059
rect 6193 14025 6227 14059
rect 6561 14025 6595 14059
rect 7481 14025 7515 14059
rect 7941 14025 7975 14059
rect 10885 14025 10919 14059
rect 11529 14025 11563 14059
rect 12725 14025 12759 14059
rect 15393 14025 15427 14059
rect 16865 14025 16899 14059
rect 17141 14025 17175 14059
rect 25789 14025 25823 14059
rect 3985 13957 4019 13991
rect 1961 13889 1995 13923
rect 2881 13889 2915 13923
rect 3065 13889 3099 13923
rect 4629 13889 4663 13923
rect 7849 13889 7883 13923
rect 8493 13889 8527 13923
rect 9413 13889 9447 13923
rect 12173 13889 12207 13923
rect 24317 13889 24351 13923
rect 2789 13821 2823 13855
rect 3525 13821 3559 13855
rect 3893 13821 3927 13855
rect 4445 13821 4479 13855
rect 5549 13821 5583 13855
rect 9505 13821 9539 13855
rect 9772 13821 9806 13855
rect 13093 13821 13127 13855
rect 13185 13821 13219 13855
rect 15485 13821 15519 13855
rect 15741 13821 15775 13855
rect 24409 13821 24443 13855
rect 24676 13821 24710 13855
rect 1409 13753 1443 13787
rect 8309 13753 8343 13787
rect 11437 13753 11471 13787
rect 11897 13753 11931 13787
rect 2329 13685 2363 13719
rect 4353 13685 4387 13719
rect 4997 13685 5031 13719
rect 6837 13685 6871 13719
rect 8401 13685 8435 13719
rect 9045 13685 9079 13719
rect 11989 13685 12023 13719
rect 14473 13685 14507 13719
rect 1961 13481 1995 13515
rect 2881 13481 2915 13515
rect 4077 13481 4111 13515
rect 5825 13481 5859 13515
rect 6929 13481 6963 13515
rect 7389 13481 7423 13515
rect 7757 13481 7791 13515
rect 8769 13481 8803 13515
rect 8953 13481 8987 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 10793 13481 10827 13515
rect 11437 13481 11471 13515
rect 12357 13481 12391 13515
rect 12725 13481 12759 13515
rect 13461 13481 13495 13515
rect 15577 13481 15611 13515
rect 2329 13413 2363 13447
rect 7849 13413 7883 13447
rect 12081 13413 12115 13447
rect 16681 13413 16715 13447
rect 24409 13413 24443 13447
rect 2789 13345 2823 13379
rect 3893 13345 3927 13379
rect 4445 13345 4479 13379
rect 5365 13345 5399 13379
rect 6193 13345 6227 13379
rect 7205 13345 7239 13379
rect 9137 13345 9171 13379
rect 11713 13345 11747 13379
rect 12817 13345 12851 13379
rect 15117 13345 15151 13379
rect 15945 13345 15979 13379
rect 1409 13277 1443 13311
rect 2973 13277 3007 13311
rect 4537 13277 4571 13311
rect 4721 13277 4755 13311
rect 5733 13277 5767 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 7941 13277 7975 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 12909 13277 12943 13311
rect 16037 13277 16071 13311
rect 16221 13277 16255 13311
rect 17141 13277 17175 13311
rect 2421 13209 2455 13243
rect 8493 13209 8527 13243
rect 11529 13209 11563 13243
rect 14473 13209 14507 13243
rect 3525 13141 3559 13175
rect 9413 13141 9447 13175
rect 13737 13141 13771 13175
rect 14105 13141 14139 13175
rect 1593 12937 1627 12971
rect 2513 12937 2547 12971
rect 4813 12937 4847 12971
rect 5825 12937 5859 12971
rect 7389 12937 7423 12971
rect 8861 12937 8895 12971
rect 10609 12937 10643 12971
rect 11621 12937 11655 12971
rect 12265 12937 12299 12971
rect 14933 12937 14967 12971
rect 15761 12937 15795 12971
rect 17141 12937 17175 12971
rect 3985 12869 4019 12903
rect 10333 12869 10367 12903
rect 10977 12869 11011 12903
rect 16773 12869 16807 12903
rect 5365 12801 5399 12835
rect 8033 12801 8067 12835
rect 8953 12801 8987 12835
rect 12725 12801 12759 12835
rect 13553 12801 13587 12835
rect 15577 12801 15611 12835
rect 16221 12801 16255 12835
rect 16313 12801 16347 12835
rect 1409 12733 1443 12767
rect 2605 12733 2639 12767
rect 4353 12733 4387 12767
rect 5181 12733 5215 12767
rect 6653 12733 6687 12767
rect 7757 12733 7791 12767
rect 9220 12733 9254 12767
rect 15301 12733 15335 12767
rect 16129 12733 16163 12767
rect 2145 12665 2179 12699
rect 2872 12665 2906 12699
rect 7297 12665 7331 12699
rect 7849 12665 7883 12699
rect 8493 12665 8527 12699
rect 13461 12665 13495 12699
rect 13798 12665 13832 12699
rect 4721 12597 4755 12631
rect 5273 12597 5307 12631
rect 6285 12597 6319 12631
rect 13001 12597 13035 12631
rect 3157 12393 3191 12427
rect 3893 12393 3927 12427
rect 4077 12393 4111 12427
rect 5733 12393 5767 12427
rect 7205 12393 7239 12427
rect 9689 12393 9723 12427
rect 12909 12393 12943 12427
rect 13553 12393 13587 12427
rect 15025 12393 15059 12427
rect 15761 12393 15795 12427
rect 16313 12393 16347 12427
rect 17325 12393 17359 12427
rect 1685 12325 1719 12359
rect 6193 12325 6227 12359
rect 6929 12325 6963 12359
rect 11774 12325 11808 12359
rect 17233 12325 17267 12359
rect 1777 12257 1811 12291
rect 2033 12257 2067 12291
rect 4445 12257 4479 12291
rect 6101 12257 6135 12291
rect 7656 12257 7690 12291
rect 10057 12257 10091 12291
rect 14933 12257 14967 12291
rect 15669 12257 15703 12291
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 6285 12189 6319 12223
rect 7389 12189 7423 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11529 12189 11563 12223
rect 5641 12121 5675 12155
rect 10701 12121 10735 12155
rect 15853 12189 15887 12223
rect 17509 12189 17543 12223
rect 16865 12121 16899 12155
rect 3433 12053 3467 12087
rect 5089 12053 5123 12087
rect 8769 12053 8803 12087
rect 9413 12053 9447 12087
rect 11437 12053 11471 12087
rect 13277 12053 13311 12087
rect 13921 12053 13955 12087
rect 14289 12053 14323 12087
rect 14657 12053 14691 12087
rect 14933 12053 14967 12087
rect 15301 12053 15335 12087
rect 3433 11849 3467 11883
rect 3709 11849 3743 11883
rect 5365 11849 5399 11883
rect 6193 11849 6227 11883
rect 6653 11849 6687 11883
rect 9321 11849 9355 11883
rect 10701 11849 10735 11883
rect 14105 11849 14139 11883
rect 14565 11849 14599 11883
rect 15393 11849 15427 11883
rect 16497 11849 16531 11883
rect 17325 11849 17359 11883
rect 17601 11849 17635 11883
rect 3157 11781 3191 11815
rect 1777 11713 1811 11747
rect 3985 11781 4019 11815
rect 8217 11781 8251 11815
rect 8861 11781 8895 11815
rect 4537 11713 4571 11747
rect 4997 11713 5031 11747
rect 9873 11713 9907 11747
rect 16037 11713 16071 11747
rect 3709 11645 3743 11679
rect 4353 11645 4387 11679
rect 6837 11645 6871 11679
rect 12173 11645 12207 11679
rect 12725 11645 12759 11679
rect 12992 11645 13026 11679
rect 1685 11577 1719 11611
rect 2022 11577 2056 11611
rect 7104 11577 7138 11611
rect 9781 11577 9815 11611
rect 11345 11577 11379 11611
rect 15209 11577 15243 11611
rect 15761 11577 15795 11611
rect 3801 11509 3835 11543
rect 4445 11509 4479 11543
rect 5733 11509 5767 11543
rect 9229 11509 9263 11543
rect 9689 11509 9723 11543
rect 10425 11509 10459 11543
rect 11161 11509 11195 11543
rect 11805 11509 11839 11543
rect 14933 11509 14967 11543
rect 15853 11509 15887 11543
rect 16865 11509 16899 11543
rect 1869 11305 1903 11339
rect 3893 11305 3927 11339
rect 4077 11305 4111 11339
rect 5641 11305 5675 11339
rect 7481 11305 7515 11339
rect 9413 11305 9447 11339
rect 9689 11305 9723 11339
rect 12817 11305 12851 11339
rect 14749 11305 14783 11339
rect 15117 11305 15151 11339
rect 15761 11305 15795 11339
rect 16865 11305 16899 11339
rect 17233 11305 17267 11339
rect 3525 11237 3559 11271
rect 4445 11237 4479 11271
rect 8493 11237 8527 11271
rect 10057 11237 10091 11271
rect 11621 11237 11655 11271
rect 13185 11237 13219 11271
rect 16773 11237 16807 11271
rect 2421 11169 2455 11203
rect 6009 11169 6043 11203
rect 6101 11169 6135 11203
rect 8401 11169 8435 11203
rect 12633 11169 12667 11203
rect 15669 11169 15703 11203
rect 17325 11169 17359 11203
rect 2513 11101 2547 11135
rect 2605 11101 2639 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 6285 11101 6319 11135
rect 8585 11101 8619 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11713 11101 11747 11135
rect 11805 11101 11839 11135
rect 2053 11033 2087 11067
rect 3065 11033 3099 11067
rect 5273 11033 5307 11067
rect 7849 11033 7883 11067
rect 8033 11033 8067 11067
rect 10885 11033 10919 11067
rect 11253 11033 11287 11067
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 15853 11101 15887 11135
rect 17509 11101 17543 11135
rect 15301 11033 15335 11067
rect 6929 10965 6963 10999
rect 12541 10965 12575 10999
rect 12633 10965 12667 10999
rect 14105 10965 14139 10999
rect 16313 10965 16347 10999
rect 1409 10761 1443 10795
rect 2881 10761 2915 10795
rect 5181 10761 5215 10795
rect 6561 10761 6595 10795
rect 7481 10761 7515 10795
rect 10057 10761 10091 10795
rect 12173 10761 12207 10795
rect 13553 10761 13587 10795
rect 15393 10761 15427 10795
rect 16957 10761 16991 10795
rect 7849 10693 7883 10727
rect 9413 10693 9447 10727
rect 1961 10625 1995 10659
rect 5825 10625 5859 10659
rect 7113 10625 7147 10659
rect 10609 10625 10643 10659
rect 11437 10625 11471 10659
rect 11897 10625 11931 10659
rect 13001 10625 13035 10659
rect 13921 10625 13955 10659
rect 14565 10625 14599 10659
rect 16129 10625 16163 10659
rect 17233 10625 17267 10659
rect 2973 10557 3007 10591
rect 3229 10557 3263 10591
rect 4629 10557 4663 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 8033 10557 8067 10591
rect 8300 10557 8334 10591
rect 11161 10557 11195 10591
rect 12817 10557 12851 10591
rect 16037 10557 16071 10591
rect 1869 10489 1903 10523
rect 12909 10489 12943 10523
rect 14473 10489 14507 10523
rect 15025 10489 15059 10523
rect 15945 10489 15979 10523
rect 1777 10421 1811 10455
rect 2513 10421 2547 10455
rect 4353 10421 4387 10455
rect 4997 10421 5031 10455
rect 6285 10421 6319 10455
rect 9781 10421 9815 10455
rect 10793 10421 10827 10455
rect 11253 10421 11287 10455
rect 12449 10421 12483 10455
rect 14013 10421 14047 10455
rect 14381 10421 14415 10455
rect 15577 10421 15611 10455
rect 17601 10421 17635 10455
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 2789 10217 2823 10251
rect 4077 10217 4111 10251
rect 7481 10217 7515 10251
rect 8493 10217 8527 10251
rect 9413 10217 9447 10251
rect 11437 10217 11471 10251
rect 11805 10217 11839 10251
rect 14749 10217 14783 10251
rect 16773 10217 16807 10251
rect 17049 10217 17083 10251
rect 3433 10149 3467 10183
rect 3893 10149 3927 10183
rect 4445 10149 4479 10183
rect 15025 10149 15059 10183
rect 2329 10081 2363 10115
rect 2881 10081 2915 10115
rect 5641 10081 5675 10115
rect 6101 10081 6135 10115
rect 6368 10081 6402 10115
rect 8125 10081 8159 10115
rect 8585 10081 8619 10115
rect 9956 10081 9990 10115
rect 12173 10081 12207 10115
rect 12532 10081 12566 10115
rect 15669 10081 15703 10115
rect 1409 10013 1443 10047
rect 3065 10013 3099 10047
rect 4537 10013 4571 10047
rect 4629 10013 4663 10047
rect 9689 10013 9723 10047
rect 12265 10013 12299 10047
rect 15761 10013 15795 10047
rect 15853 10013 15887 10047
rect 15301 9945 15335 9979
rect 5181 9877 5215 9911
rect 9045 9877 9079 9911
rect 11069 9877 11103 9911
rect 11989 9877 12023 9911
rect 13645 9877 13679 9911
rect 14013 9877 14047 9911
rect 16313 9877 16347 9911
rect 13461 9673 13495 9707
rect 14933 9673 14967 9707
rect 2697 9605 2731 9639
rect 4997 9605 5031 9639
rect 6837 9605 6871 9639
rect 11805 9605 11839 9639
rect 12265 9605 12299 9639
rect 15577 9605 15611 9639
rect 16773 9605 16807 9639
rect 1685 9537 1719 9571
rect 5549 9537 5583 9571
rect 6653 9537 6687 9571
rect 7481 9537 7515 9571
rect 8861 9537 8895 9571
rect 8953 9537 8987 9571
rect 12449 9537 12483 9571
rect 16313 9537 16347 9571
rect 1409 9469 1443 9503
rect 2796 9469 2830 9503
rect 3056 9469 3090 9503
rect 7849 9469 7883 9503
rect 8309 9469 8343 9503
rect 8769 9469 8803 9503
rect 10149 9469 10183 9503
rect 10416 9469 10450 9503
rect 13553 9469 13587 9503
rect 13809 9469 13843 9503
rect 16129 9469 16163 9503
rect 6193 9401 6227 9435
rect 9689 9401 9723 9435
rect 10057 9401 10091 9435
rect 16221 9401 16255 9435
rect 2329 9333 2363 9367
rect 4169 9333 4203 9367
rect 4445 9333 4479 9367
rect 4813 9333 4847 9367
rect 5365 9333 5399 9367
rect 5457 9333 5491 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 8401 9333 8435 9367
rect 11529 9333 11563 9367
rect 13001 9333 13035 9367
rect 15301 9333 15335 9367
rect 15761 9333 15795 9367
rect 17233 9333 17267 9367
rect 17601 9333 17635 9367
rect 2789 9129 2823 9163
rect 3157 9129 3191 9163
rect 3525 9129 3559 9163
rect 4077 9129 4111 9163
rect 7941 9129 7975 9163
rect 9689 9129 9723 9163
rect 10057 9129 10091 9163
rect 12357 9129 12391 9163
rect 12909 9129 12943 9163
rect 16773 9129 16807 9163
rect 1676 9061 1710 9095
rect 3801 9061 3835 9095
rect 4537 9061 4571 9095
rect 9413 9061 9447 9095
rect 10149 9061 10183 9095
rect 13461 9061 13495 9095
rect 13829 9061 13863 9095
rect 14197 9061 14231 9095
rect 1409 8993 1443 9027
rect 4445 8993 4479 9027
rect 5825 8993 5859 9027
rect 6092 8993 6126 9027
rect 8401 8993 8435 9027
rect 10793 8993 10827 9027
rect 12817 8993 12851 9027
rect 15669 8993 15703 9027
rect 4629 8925 4663 8959
rect 5457 8925 5491 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 9045 8925 9079 8959
rect 10241 8925 10275 8959
rect 13093 8925 13127 8959
rect 15117 8925 15151 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 8033 8857 8067 8891
rect 11621 8857 11655 8891
rect 12449 8857 12483 8891
rect 5181 8789 5215 8823
rect 7205 8789 7239 8823
rect 7481 8789 7515 8823
rect 11253 8789 11287 8823
rect 11897 8789 11931 8823
rect 14657 8789 14691 8823
rect 15301 8789 15335 8823
rect 16497 8789 16531 8823
rect 17233 8789 17267 8823
rect 17601 8789 17635 8823
rect 1777 8585 1811 8619
rect 3617 8585 3651 8619
rect 6561 8585 6595 8619
rect 8033 8585 8067 8619
rect 8585 8585 8619 8619
rect 9781 8585 9815 8619
rect 10793 8585 10827 8619
rect 13553 8585 13587 8619
rect 14105 8585 14139 8619
rect 16313 8585 16347 8619
rect 4077 8517 4111 8551
rect 10609 8517 10643 8551
rect 12541 8517 12575 8551
rect 15577 8517 15611 8551
rect 15945 8517 15979 8551
rect 1869 8449 1903 8483
rect 4629 8449 4663 8483
rect 5457 8449 5491 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 9137 8449 9171 8483
rect 11345 8449 11379 8483
rect 13001 8449 13035 8483
rect 13185 8449 13219 8483
rect 14197 8449 14231 8483
rect 16957 8449 16991 8483
rect 2125 8381 2159 8415
rect 3985 8381 4019 8415
rect 4445 8381 4479 8415
rect 5089 8381 5123 8415
rect 8401 8381 8435 8415
rect 8953 8381 8987 8415
rect 10333 8381 10367 8415
rect 11161 8381 11195 8415
rect 11897 8381 11931 8415
rect 16865 8381 16899 8415
rect 17509 8381 17543 8415
rect 5641 8313 5675 8347
rect 6285 8313 6319 8347
rect 7205 8313 7239 8347
rect 11253 8313 11287 8347
rect 12173 8313 12207 8347
rect 14464 8313 14498 8347
rect 16773 8313 16807 8347
rect 17877 8313 17911 8347
rect 3249 8245 3283 8279
rect 4537 8245 4571 8279
rect 6837 8245 6871 8279
rect 9045 8245 9079 8279
rect 10149 8245 10183 8279
rect 12909 8245 12943 8279
rect 16405 8245 16439 8279
rect 2237 8041 2271 8075
rect 2605 8041 2639 8075
rect 3249 8041 3283 8075
rect 3893 8041 3927 8075
rect 4905 8041 4939 8075
rect 5549 8041 5583 8075
rect 7113 8041 7147 8075
rect 7205 8041 7239 8075
rect 8033 8041 8067 8075
rect 8493 8041 8527 8075
rect 9965 8041 9999 8075
rect 10241 8041 10275 8075
rect 13369 8041 13403 8075
rect 13829 8041 13863 8075
rect 15301 8041 15335 8075
rect 16221 8041 16255 8075
rect 17693 8041 17727 8075
rect 16580 7973 16614 8007
rect 18981 7973 19015 8007
rect 2697 7905 2731 7939
rect 5089 7905 5123 7939
rect 8585 7905 8619 7939
rect 9505 7905 9539 7939
rect 10701 7905 10735 7939
rect 10957 7905 10991 7939
rect 13737 7905 13771 7939
rect 18889 7905 18923 7939
rect 2881 7837 2915 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 7297 7837 7331 7871
rect 12541 7837 12575 7871
rect 13921 7837 13955 7871
rect 15853 7837 15887 7871
rect 16313 7837 16347 7871
rect 19073 7837 19107 7871
rect 4813 7769 4847 7803
rect 6653 7769 6687 7803
rect 14565 7769 14599 7803
rect 1685 7701 1719 7735
rect 2053 7701 2087 7735
rect 4261 7701 4295 7735
rect 5181 7701 5215 7735
rect 6285 7701 6319 7735
rect 6745 7701 6779 7735
rect 9137 7701 9171 7735
rect 12081 7701 12115 7735
rect 13185 7701 13219 7735
rect 14841 7701 14875 7735
rect 18061 7701 18095 7735
rect 18521 7701 18555 7735
rect 5181 7497 5215 7531
rect 6285 7497 6319 7531
rect 7849 7497 7883 7531
rect 10793 7497 10827 7531
rect 13001 7497 13035 7531
rect 16957 7497 16991 7531
rect 17417 7497 17451 7531
rect 19073 7497 19107 7531
rect 2513 7429 2547 7463
rect 4721 7429 4755 7463
rect 11805 7429 11839 7463
rect 15485 7429 15519 7463
rect 2053 7361 2087 7395
rect 3525 7361 3559 7395
rect 3617 7361 3651 7395
rect 5825 7361 5859 7395
rect 7389 7361 7423 7395
rect 8677 7361 8711 7395
rect 11345 7361 11379 7395
rect 13093 7361 13127 7395
rect 15117 7361 15151 7395
rect 16037 7361 16071 7395
rect 16129 7361 16163 7395
rect 18613 7361 18647 7395
rect 1869 7293 1903 7327
rect 2973 7293 3007 7327
rect 3433 7293 3467 7327
rect 5549 7293 5583 7327
rect 7205 7293 7239 7327
rect 10425 7293 10459 7327
rect 15945 7293 15979 7327
rect 17785 7293 17819 7327
rect 18429 7293 18463 7327
rect 19441 7293 19475 7327
rect 1961 7225 1995 7259
rect 4997 7225 5031 7259
rect 5641 7225 5675 7259
rect 8585 7225 8619 7259
rect 8944 7225 8978 7259
rect 12173 7225 12207 7259
rect 13360 7225 13394 7259
rect 1501 7157 1535 7191
rect 3065 7157 3099 7191
rect 4353 7157 4387 7191
rect 6561 7157 6595 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 10057 7157 10091 7191
rect 11161 7157 11195 7191
rect 14473 7157 14507 7191
rect 15577 7157 15611 7191
rect 16681 7157 16715 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 3617 6953 3651 6987
rect 4721 6953 4755 6987
rect 6193 6953 6227 6987
rect 6561 6953 6595 6987
rect 8769 6953 8803 6987
rect 13461 6953 13495 6987
rect 13737 6953 13771 6987
rect 18797 6953 18831 6987
rect 1860 6885 1894 6919
rect 3341 6885 3375 6919
rect 7288 6885 7322 6919
rect 16190 6885 16224 6919
rect 1593 6817 1627 6851
rect 4813 6817 4847 6851
rect 5080 6817 5114 6851
rect 7021 6817 7055 6851
rect 9945 6817 9979 6851
rect 12348 6817 12382 6851
rect 17601 6817 17635 6851
rect 17969 6817 18003 6851
rect 18153 6817 18187 6851
rect 9689 6749 9723 6783
rect 12081 6749 12115 6783
rect 15945 6749 15979 6783
rect 19073 6749 19107 6783
rect 11069 6681 11103 6715
rect 19533 6681 19567 6715
rect 2973 6613 3007 6647
rect 4353 6613 4387 6647
rect 6929 6613 6963 6647
rect 8401 6613 8435 6647
rect 9045 6613 9079 6647
rect 9413 6613 9447 6647
rect 11437 6613 11471 6647
rect 11713 6613 11747 6647
rect 14105 6613 14139 6647
rect 14749 6613 14783 6647
rect 15117 6613 15151 6647
rect 15853 6613 15887 6647
rect 17325 6613 17359 6647
rect 18337 6613 18371 6647
rect 19901 6613 19935 6647
rect 3617 6409 3651 6443
rect 4353 6409 4387 6443
rect 6561 6409 6595 6443
rect 7849 6409 7883 6443
rect 10057 6409 10091 6443
rect 12081 6409 12115 6443
rect 15117 6409 15151 6443
rect 16957 6409 16991 6443
rect 17785 6409 17819 6443
rect 19441 6409 19475 6443
rect 5181 6341 5215 6375
rect 6193 6341 6227 6375
rect 10333 6341 10367 6375
rect 1501 6273 1535 6307
rect 3709 6273 3743 6307
rect 5825 6273 5859 6307
rect 7389 6273 7423 6307
rect 8677 6273 8711 6307
rect 15485 6273 15519 6307
rect 18613 6273 18647 6307
rect 7205 6205 7239 6239
rect 11253 6205 11287 6239
rect 12725 6205 12759 6239
rect 14381 6205 14415 6239
rect 15577 6205 15611 6239
rect 15844 6205 15878 6239
rect 18429 6205 18463 6239
rect 19073 6205 19107 6239
rect 1768 6137 1802 6171
rect 5549 6137 5583 6171
rect 8585 6137 8619 6171
rect 8944 6137 8978 6171
rect 12992 6137 13026 6171
rect 17509 6137 17543 6171
rect 18521 6137 18555 6171
rect 19901 6137 19935 6171
rect 2881 6069 2915 6103
rect 3157 6069 3191 6103
rect 4629 6069 4663 6103
rect 4997 6069 5031 6103
rect 5641 6069 5675 6103
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 10793 6069 10827 6103
rect 11161 6069 11195 6103
rect 11437 6069 11471 6103
rect 14105 6069 14139 6103
rect 18061 6069 18095 6103
rect 20269 6069 20303 6103
rect 2053 5865 2087 5899
rect 3709 5865 3743 5899
rect 4905 5865 4939 5899
rect 6929 5865 6963 5899
rect 7389 5865 7423 5899
rect 8585 5865 8619 5899
rect 9321 5865 9355 5899
rect 10057 5865 10091 5899
rect 11253 5865 11287 5899
rect 12817 5865 12851 5899
rect 13277 5865 13311 5899
rect 16221 5865 16255 5899
rect 16773 5865 16807 5899
rect 17325 5865 17359 5899
rect 19349 5865 19383 5899
rect 4261 5797 4295 5831
rect 5448 5797 5482 5831
rect 8953 5797 8987 5831
rect 11713 5797 11747 5831
rect 16129 5797 16163 5831
rect 18337 5797 18371 5831
rect 18705 5797 18739 5831
rect 2605 5729 2639 5763
rect 3249 5729 3283 5763
rect 5181 5729 5215 5763
rect 7757 5729 7791 5763
rect 11621 5729 11655 5763
rect 13369 5729 13403 5763
rect 14289 5729 14323 5763
rect 14657 5729 14691 5763
rect 17693 5729 17727 5763
rect 19257 5729 19291 5763
rect 22477 5729 22511 5763
rect 2697 5661 2731 5695
rect 2881 5661 2915 5695
rect 7297 5661 7331 5695
rect 7849 5661 7883 5695
rect 8033 5661 8067 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 11897 5661 11931 5695
rect 13461 5661 13495 5695
rect 16313 5661 16347 5695
rect 17785 5661 17819 5695
rect 17877 5661 17911 5695
rect 19441 5661 19475 5695
rect 20729 5661 20763 5695
rect 22753 5661 22787 5695
rect 1685 5593 1719 5627
rect 9689 5593 9723 5627
rect 12909 5593 12943 5627
rect 14933 5593 14967 5627
rect 15669 5593 15703 5627
rect 17141 5593 17175 5627
rect 18889 5593 18923 5627
rect 2237 5525 2271 5559
rect 6561 5525 6595 5559
rect 10793 5525 10827 5559
rect 12449 5525 12483 5559
rect 13921 5525 13955 5559
rect 14473 5525 14507 5559
rect 15761 5525 15795 5559
rect 19993 5525 20027 5559
rect 20361 5525 20395 5559
rect 2421 5321 2455 5355
rect 5273 5321 5307 5355
rect 5641 5321 5675 5355
rect 9045 5321 9079 5355
rect 9229 5321 9263 5355
rect 10241 5321 10275 5355
rect 10609 5321 10643 5355
rect 11805 5321 11839 5355
rect 12265 5321 12299 5355
rect 12817 5321 12851 5355
rect 12909 5321 12943 5355
rect 15853 5321 15887 5355
rect 16037 5321 16071 5355
rect 18061 5321 18095 5355
rect 19165 5321 19199 5355
rect 19809 5321 19843 5355
rect 3985 5253 4019 5287
rect 6193 5253 6227 5287
rect 14473 5253 14507 5287
rect 3065 5185 3099 5219
rect 4537 5185 4571 5219
rect 9689 5185 9723 5219
rect 9781 5185 9815 5219
rect 11345 5185 11379 5219
rect 13369 5185 13403 5219
rect 13553 5185 13587 5219
rect 15117 5185 15151 5219
rect 16589 5185 16623 5219
rect 18613 5185 18647 5219
rect 19441 5185 19475 5219
rect 2329 5117 2363 5151
rect 3525 5117 3559 5151
rect 6929 5117 6963 5151
rect 8769 5117 8803 5151
rect 9597 5117 9631 5151
rect 11253 5117 11287 5151
rect 13277 5117 13311 5151
rect 14381 5117 14415 5151
rect 14841 5117 14875 5151
rect 18429 5117 18463 5151
rect 18521 5117 18555 5151
rect 20269 5117 20303 5151
rect 21005 5117 21039 5151
rect 22477 5117 22511 5151
rect 23673 5117 23707 5151
rect 24225 5117 24259 5151
rect 2881 5049 2915 5083
rect 4353 5049 4387 5083
rect 6561 5049 6595 5083
rect 7174 5049 7208 5083
rect 16497 5049 16531 5083
rect 20545 5049 20579 5083
rect 1869 4981 1903 5015
rect 2789 4981 2823 5015
rect 3801 4981 3835 5015
rect 4445 4981 4479 5015
rect 5733 4981 5767 5015
rect 8309 4981 8343 5015
rect 10793 4981 10827 5015
rect 11161 4981 11195 5015
rect 14013 4981 14047 5015
rect 14933 4981 14967 5015
rect 16405 4981 16439 5015
rect 17325 4981 17359 5015
rect 17693 4981 17727 5015
rect 23857 4981 23891 5015
rect 1869 4777 1903 4811
rect 2329 4777 2363 4811
rect 3249 4777 3283 4811
rect 5825 4777 5859 4811
rect 5917 4777 5951 4811
rect 7021 4777 7055 4811
rect 7389 4777 7423 4811
rect 8033 4777 8067 4811
rect 9505 4777 9539 4811
rect 10885 4777 10919 4811
rect 11437 4777 11471 4811
rect 11805 4777 11839 4811
rect 13001 4777 13035 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15025 4777 15059 4811
rect 16957 4777 16991 4811
rect 17417 4777 17451 4811
rect 17785 4777 17819 4811
rect 19165 4777 19199 4811
rect 20085 4777 20119 4811
rect 22109 4777 22143 4811
rect 2973 4709 3007 4743
rect 4353 4709 4387 4743
rect 6929 4709 6963 4743
rect 10057 4709 10091 4743
rect 11345 4709 11379 4743
rect 19625 4709 19659 4743
rect 2237 4641 2271 4675
rect 4087 4641 4121 4675
rect 7481 4641 7515 4675
rect 13553 4641 13587 4675
rect 14749 4641 14783 4675
rect 15844 4641 15878 4675
rect 18153 4641 18187 4675
rect 19349 4641 19383 4675
rect 21189 4641 21223 4675
rect 22293 4641 22327 4675
rect 2421 4573 2455 4607
rect 4813 4573 4847 4607
rect 6101 4573 6135 4607
rect 7665 4573 7699 4607
rect 8585 4573 8619 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 15577 4573 15611 4607
rect 18245 4573 18279 4607
rect 18337 4573 18371 4607
rect 20453 4573 20487 4607
rect 5273 4505 5307 4539
rect 1685 4437 1719 4471
rect 3709 4437 3743 4471
rect 5457 4437 5491 4471
rect 6469 4437 6503 4471
rect 8493 4437 8527 4471
rect 9137 4437 9171 4471
rect 9689 4437 9723 4471
rect 12541 4437 12575 4471
rect 18797 4437 18831 4471
rect 21373 4437 21407 4471
rect 21833 4437 21867 4471
rect 22477 4437 22511 4471
rect 6561 4233 6595 4267
rect 10149 4233 10183 4267
rect 14013 4233 14047 4267
rect 19441 4233 19475 4267
rect 20637 4233 20671 4267
rect 21005 4233 21039 4267
rect 3341 4165 3375 4199
rect 8309 4165 8343 4199
rect 1961 4097 1995 4131
rect 3985 4097 4019 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6285 4097 6319 4131
rect 7849 4097 7883 4131
rect 8585 4097 8619 4131
rect 9321 4097 9355 4131
rect 10701 4097 10735 4131
rect 11345 4097 11379 4131
rect 13001 4097 13035 4131
rect 17785 4097 17819 4131
rect 18613 4097 18647 4131
rect 20269 4097 20303 4131
rect 5641 4029 5675 4063
rect 7665 4029 7699 4063
rect 9137 4029 9171 4063
rect 11161 4029 11195 4063
rect 12817 4029 12851 4063
rect 14289 4029 14323 4063
rect 16497 4029 16531 4063
rect 17509 4029 17543 4063
rect 18429 4029 18463 4063
rect 19993 4029 20027 4063
rect 21189 4029 21223 4063
rect 21741 4029 21775 4063
rect 22293 4029 22327 4063
rect 22845 4029 22879 4063
rect 2228 3961 2262 3995
rect 5549 3961 5583 3995
rect 9229 3961 9263 3995
rect 13737 3961 13771 3995
rect 14534 3961 14568 3995
rect 16313 3961 16347 3995
rect 16773 3961 16807 3995
rect 18521 3961 18555 3995
rect 19073 3961 19107 3995
rect 1869 3893 1903 3927
rect 3709 3893 3743 3927
rect 4169 3893 4203 3927
rect 4721 3893 4755 3927
rect 5181 3893 5215 3927
rect 7021 3893 7055 3927
rect 7205 3893 7239 3927
rect 7573 3893 7607 3927
rect 8769 3893 8803 3927
rect 9781 3893 9815 3927
rect 10793 3893 10827 3927
rect 11253 3893 11287 3927
rect 11805 3893 11839 3927
rect 12173 3893 12207 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 15669 3893 15703 3927
rect 16037 3893 16071 3927
rect 18061 3893 18095 3927
rect 19625 3893 19659 3927
rect 20085 3893 20119 3927
rect 21373 3893 21407 3927
rect 22109 3893 22143 3927
rect 22477 3893 22511 3927
rect 1685 3689 1719 3723
rect 3157 3689 3191 3723
rect 3893 3689 3927 3723
rect 5825 3689 5859 3723
rect 6193 3689 6227 3723
rect 7665 3689 7699 3723
rect 8401 3689 8435 3723
rect 8861 3689 8895 3723
rect 9137 3689 9171 3723
rect 9413 3689 9447 3723
rect 10885 3689 10919 3723
rect 13093 3689 13127 3723
rect 13185 3689 13219 3723
rect 13369 3689 13403 3723
rect 15577 3689 15611 3723
rect 16037 3689 16071 3723
rect 17141 3689 17175 3723
rect 17509 3689 17543 3723
rect 18153 3689 18187 3723
rect 19073 3689 19107 3723
rect 21465 3689 21499 3723
rect 21833 3689 21867 3723
rect 22569 3689 22603 3723
rect 22937 3689 22971 3723
rect 23673 3689 23707 3723
rect 4322 3621 4356 3655
rect 6530 3621 6564 3655
rect 1777 3553 1811 3587
rect 2044 3553 2078 3587
rect 3433 3553 3467 3587
rect 8493 3553 8527 3587
rect 9873 3553 9907 3587
rect 10149 3553 10183 3587
rect 11428 3553 11462 3587
rect 13737 3621 13771 3655
rect 15945 3621 15979 3655
rect 18521 3621 18555 3655
rect 19165 3621 19199 3655
rect 13829 3553 13863 3587
rect 16957 3553 16991 3587
rect 17601 3553 17635 3587
rect 20913 3553 20947 3587
rect 22017 3553 22051 3587
rect 23121 3553 23155 3587
rect 4077 3485 4111 3519
rect 6285 3485 6319 3519
rect 8033 3485 8067 3519
rect 8861 3485 8895 3519
rect 11161 3485 11195 3519
rect 13093 3485 13127 3519
rect 13921 3485 13955 3519
rect 15117 3485 15151 3519
rect 16221 3485 16255 3519
rect 17693 3485 17727 3519
rect 19257 3485 19291 3519
rect 19717 3485 19751 3519
rect 20085 3485 20119 3519
rect 18705 3417 18739 3451
rect 22201 3417 22235 3451
rect 5457 3349 5491 3383
rect 8677 3349 8711 3383
rect 12541 3349 12575 3383
rect 12909 3349 12943 3383
rect 14381 3349 14415 3383
rect 16589 3349 16623 3383
rect 20453 3349 20487 3383
rect 21097 3349 21131 3383
rect 23305 3349 23339 3383
rect 1409 3145 1443 3179
rect 4077 3145 4111 3179
rect 5917 3145 5951 3179
rect 6929 3145 6963 3179
rect 10609 3145 10643 3179
rect 11897 3145 11931 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 15209 3145 15243 3179
rect 15669 3145 15703 3179
rect 17233 3145 17267 3179
rect 18061 3145 18095 3179
rect 19441 3145 19475 3179
rect 20913 3145 20947 3179
rect 22017 3145 22051 3179
rect 23397 3145 23431 3179
rect 2513 3077 2547 3111
rect 6101 3077 6135 3111
rect 8033 3077 8067 3111
rect 8401 3077 8435 3111
rect 10149 3077 10183 3111
rect 15577 3077 15611 3111
rect 19625 3077 19659 3111
rect 22661 3077 22695 3111
rect 2053 3009 2087 3043
rect 3433 3009 3467 3043
rect 3617 3009 3651 3043
rect 4537 3009 4571 3043
rect 1777 2941 1811 2975
rect 2881 2941 2915 2975
rect 3341 2941 3375 2975
rect 4804 2873 4838 2907
rect 7573 3009 7607 3043
rect 11253 3009 11287 3043
rect 11437 3009 11471 3043
rect 16313 3009 16347 3043
rect 16681 3009 16715 3043
rect 18613 3009 18647 3043
rect 20177 3009 20211 3043
rect 21465 3009 21499 3043
rect 6285 2941 6319 2975
rect 7297 2941 7331 2975
rect 8493 2941 8527 2975
rect 8749 2941 8783 2975
rect 12725 2941 12759 2975
rect 12981 2941 13015 2975
rect 16037 2941 16071 2975
rect 18429 2941 18463 2975
rect 20085 2941 20119 2975
rect 21189 2941 21223 2975
rect 22477 2941 22511 2975
rect 23029 2941 23063 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 6561 2873 6595 2907
rect 7389 2873 7423 2907
rect 12173 2873 12207 2907
rect 16129 2873 16163 2907
rect 17509 2873 17543 2907
rect 18521 2873 18555 2907
rect 1869 2805 1903 2839
rect 2973 2805 3007 2839
rect 6101 2805 6135 2839
rect 9873 2805 9907 2839
rect 10793 2805 10827 2839
rect 11161 2805 11195 2839
rect 14105 2805 14139 2839
rect 19073 2805 19107 2839
rect 19993 2805 20027 2839
rect 23857 2805 23891 2839
rect 1685 2601 1719 2635
rect 2053 2601 2087 2635
rect 3525 2601 3559 2635
rect 5273 2601 5307 2635
rect 6285 2601 6319 2635
rect 8125 2601 8159 2635
rect 8585 2601 8619 2635
rect 9137 2601 9171 2635
rect 10793 2601 10827 2635
rect 11345 2601 11379 2635
rect 11437 2601 11471 2635
rect 11989 2601 12023 2635
rect 13461 2601 13495 2635
rect 14013 2601 14047 2635
rect 15485 2601 15519 2635
rect 18061 2601 18095 2635
rect 18797 2601 18831 2635
rect 20821 2601 20855 2635
rect 22293 2601 22327 2635
rect 23397 2601 23431 2635
rect 2881 2533 2915 2567
rect 6745 2533 6779 2567
rect 8493 2533 8527 2567
rect 12357 2533 12391 2567
rect 12633 2533 12667 2567
rect 14381 2533 14415 2567
rect 14933 2533 14967 2567
rect 2789 2465 2823 2499
rect 3801 2465 3835 2499
rect 5641 2465 5675 2499
rect 5733 2465 5767 2499
rect 7021 2465 7055 2499
rect 9873 2465 9907 2499
rect 11805 2465 11839 2499
rect 3065 2397 3099 2431
rect 4997 2397 5031 2431
rect 5917 2397 5951 2431
rect 8033 2397 8067 2431
rect 8769 2397 8803 2431
rect 10517 2397 10551 2431
rect 11621 2397 11655 2431
rect 4445 2329 4479 2363
rect 9597 2329 9631 2363
rect 13369 2465 13403 2499
rect 15853 2465 15887 2499
rect 15945 2465 15979 2499
rect 17049 2465 17083 2499
rect 17601 2465 17635 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21189 2465 21223 2499
rect 21925 2465 21959 2499
rect 22477 2465 22511 2499
rect 23029 2465 23063 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 25697 2465 25731 2499
rect 13645 2397 13679 2431
rect 16037 2397 16071 2431
rect 16497 2397 16531 2431
rect 16957 2397 16991 2431
rect 18889 2397 18923 2431
rect 21373 2397 21407 2431
rect 12633 2329 12667 2363
rect 12909 2329 12943 2363
rect 20085 2329 20119 2363
rect 22661 2329 22695 2363
rect 2421 2261 2455 2295
rect 4721 2261 4755 2295
rect 4997 2261 5031 2295
rect 5181 2261 5215 2295
rect 7205 2261 7239 2295
rect 7665 2261 7699 2295
rect 10057 2261 10091 2295
rect 10977 2261 11011 2295
rect 11805 2261 11839 2295
rect 13001 2261 13035 2295
rect 15209 2261 15243 2295
rect 17233 2261 17267 2295
rect 18337 2261 18371 2295
rect 19717 2261 19751 2295
rect 24225 2261 24259 2295
rect 25329 2261 25363 2295
<< metal1 >>
rect 4890 26460 4896 26512
rect 4948 26500 4954 26512
rect 12618 26500 12624 26512
rect 4948 26472 12624 26500
rect 4948 26460 4954 26472
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 3970 26324 3976 26376
rect 4028 26364 4034 26376
rect 4028 26336 8064 26364
rect 4028 26324 4034 26336
rect 8036 26296 8064 26336
rect 13722 26296 13728 26308
rect 8036 26268 13728 26296
rect 13722 26256 13728 26268
rect 13780 26256 13786 26308
rect 2406 25984 2412 26036
rect 2464 26024 2470 26036
rect 9674 26024 9680 26036
rect 2464 25996 9680 26024
rect 2464 25984 2470 25996
rect 9674 25984 9680 25996
rect 9732 25984 9738 26036
rect 7466 25916 7472 25968
rect 7524 25956 7530 25968
rect 12434 25956 12440 25968
rect 7524 25928 12440 25956
rect 7524 25916 7530 25928
rect 12434 25916 12440 25928
rect 12492 25916 12498 25968
rect 3234 25848 3240 25900
rect 3292 25888 3298 25900
rect 12526 25888 12532 25900
rect 3292 25860 12532 25888
rect 3292 25848 3298 25860
rect 12526 25848 12532 25860
rect 12584 25848 12590 25900
rect 3970 25780 3976 25832
rect 4028 25820 4034 25832
rect 11238 25820 11244 25832
rect 4028 25792 11244 25820
rect 4028 25780 4034 25792
rect 11238 25780 11244 25792
rect 11296 25780 11302 25832
rect 3050 25712 3056 25764
rect 3108 25752 3114 25764
rect 5350 25752 5356 25764
rect 3108 25724 5356 25752
rect 3108 25712 3114 25724
rect 5350 25712 5356 25724
rect 5408 25712 5414 25764
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 11054 25684 11060 25696
rect 4120 25656 11060 25684
rect 4120 25644 4126 25656
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 4120 25452 9965 25480
rect 4120 25440 4126 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 11054 25480 11060 25492
rect 11015 25452 11060 25480
rect 9953 25443 10011 25449
rect 11054 25440 11060 25452
rect 11112 25440 11118 25492
rect 2041 25415 2099 25421
rect 2041 25381 2053 25415
rect 2087 25412 2099 25415
rect 7466 25412 7472 25424
rect 2087 25384 7472 25412
rect 2087 25381 2099 25384
rect 2041 25375 2099 25381
rect 7466 25372 7472 25384
rect 7524 25372 7530 25424
rect 1765 25347 1823 25353
rect 1765 25313 1777 25347
rect 1811 25344 1823 25347
rect 2406 25344 2412 25356
rect 1811 25316 2412 25344
rect 1811 25313 1823 25316
rect 1765 25307 1823 25313
rect 2406 25304 2412 25316
rect 2464 25304 2470 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4154 25344 4160 25356
rect 4111 25316 4160 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4154 25304 4160 25316
rect 4212 25304 4218 25356
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25344 5227 25347
rect 6822 25344 6828 25356
rect 5215 25316 6828 25344
rect 5215 25313 5227 25316
rect 5169 25307 5227 25313
rect 6822 25304 6828 25316
rect 6880 25304 6886 25356
rect 7558 25344 7564 25356
rect 7519 25316 7564 25344
rect 7558 25304 7564 25316
rect 7616 25304 7622 25356
rect 7653 25347 7711 25353
rect 7653 25313 7665 25347
rect 7699 25344 7711 25347
rect 7834 25344 7840 25356
rect 7699 25316 7840 25344
rect 7699 25313 7711 25316
rect 7653 25307 7711 25313
rect 7834 25304 7840 25316
rect 7892 25304 7898 25356
rect 9769 25347 9827 25353
rect 9769 25313 9781 25347
rect 9815 25344 9827 25347
rect 10594 25344 10600 25356
rect 9815 25316 10600 25344
rect 9815 25313 9827 25316
rect 9769 25307 9827 25313
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 10873 25347 10931 25353
rect 10873 25313 10885 25347
rect 10919 25313 10931 25347
rect 10873 25307 10931 25313
rect 1854 25236 1860 25288
rect 1912 25276 1918 25288
rect 7745 25279 7803 25285
rect 1912 25248 7328 25276
rect 1912 25236 1918 25248
rect 1578 25168 1584 25220
rect 1636 25208 1642 25220
rect 1673 25211 1731 25217
rect 1673 25208 1685 25211
rect 1636 25180 1685 25208
rect 1636 25168 1642 25180
rect 1673 25177 1685 25180
rect 1719 25208 1731 25211
rect 7193 25211 7251 25217
rect 7193 25208 7205 25211
rect 1719 25180 7205 25208
rect 1719 25177 1731 25180
rect 1673 25171 1731 25177
rect 7193 25177 7205 25180
rect 7239 25177 7251 25211
rect 7300 25208 7328 25248
rect 7745 25245 7757 25279
rect 7791 25276 7803 25279
rect 8386 25276 8392 25288
rect 7791 25248 8392 25276
rect 7791 25245 7803 25248
rect 7745 25239 7803 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 10888 25208 10916 25307
rect 12526 25304 12532 25356
rect 12584 25344 12590 25356
rect 12621 25347 12679 25353
rect 12621 25344 12633 25347
rect 12584 25316 12633 25344
rect 12584 25304 12590 25316
rect 12621 25313 12633 25316
rect 12667 25344 12679 25347
rect 13354 25344 13360 25356
rect 12667 25316 13360 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 13354 25304 13360 25316
rect 13412 25304 13418 25356
rect 13630 25304 13636 25356
rect 13688 25344 13694 25356
rect 13725 25347 13783 25353
rect 13725 25344 13737 25347
rect 13688 25316 13737 25344
rect 13688 25304 13694 25316
rect 13725 25313 13737 25316
rect 13771 25313 13783 25347
rect 15470 25344 15476 25356
rect 15431 25316 15476 25344
rect 13725 25307 13783 25313
rect 15470 25304 15476 25316
rect 15528 25304 15534 25356
rect 11425 25211 11483 25217
rect 11425 25208 11437 25211
rect 7300 25180 11437 25208
rect 7193 25171 7251 25177
rect 11425 25177 11437 25180
rect 11471 25177 11483 25211
rect 11425 25171 11483 25177
rect 13909 25211 13967 25217
rect 13909 25177 13921 25211
rect 13955 25208 13967 25211
rect 24762 25208 24768 25220
rect 13955 25180 24768 25208
rect 13955 25177 13967 25180
rect 13909 25171 13967 25177
rect 24762 25168 24768 25180
rect 24820 25168 24826 25220
rect 2774 25100 2780 25152
rect 2832 25140 2838 25152
rect 4249 25143 4307 25149
rect 4249 25140 4261 25143
rect 2832 25112 4261 25140
rect 2832 25100 2838 25112
rect 4249 25109 4261 25112
rect 4295 25109 4307 25143
rect 5350 25140 5356 25152
rect 5311 25112 5356 25140
rect 4249 25103 4307 25109
rect 5350 25100 5356 25112
rect 5408 25100 5414 25152
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 5721 25143 5779 25149
rect 5721 25140 5733 25143
rect 5592 25112 5733 25140
rect 5592 25100 5598 25112
rect 5721 25109 5733 25112
rect 5767 25109 5779 25143
rect 5721 25103 5779 25109
rect 6733 25143 6791 25149
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 7834 25140 7840 25152
rect 6779 25112 7840 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 12805 25143 12863 25149
rect 12805 25140 12817 25143
rect 8352 25112 12817 25140
rect 8352 25100 8358 25112
rect 12805 25109 12817 25112
rect 12851 25109 12863 25143
rect 13538 25140 13544 25152
rect 13499 25112 13544 25140
rect 12805 25103 12863 25109
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 15657 25143 15715 25149
rect 15657 25109 15669 25143
rect 15703 25140 15715 25143
rect 26510 25140 26516 25152
rect 15703 25112 26516 25140
rect 15703 25109 15715 25112
rect 15657 25103 15715 25109
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2406 24936 2412 24948
rect 2367 24908 2412 24936
rect 2406 24896 2412 24908
rect 2464 24896 2470 24948
rect 2958 24896 2964 24948
rect 3016 24936 3022 24948
rect 5350 24936 5356 24948
rect 3016 24908 5356 24936
rect 3016 24896 3022 24908
rect 5350 24896 5356 24908
rect 5408 24896 5414 24948
rect 5534 24896 5540 24948
rect 5592 24936 5598 24948
rect 7009 24939 7067 24945
rect 7009 24936 7021 24939
rect 5592 24908 7021 24936
rect 5592 24896 5598 24908
rect 7009 24905 7021 24908
rect 7055 24905 7067 24939
rect 7009 24899 7067 24905
rect 7558 24896 7564 24948
rect 7616 24896 7622 24948
rect 10594 24936 10600 24948
rect 10555 24908 10600 24936
rect 10594 24896 10600 24908
rect 10652 24896 10658 24948
rect 12618 24936 12624 24948
rect 12579 24908 12624 24936
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 13354 24936 13360 24948
rect 13315 24908 13360 24936
rect 13354 24896 13360 24908
rect 13412 24896 13418 24948
rect 13722 24936 13728 24948
rect 13683 24908 13728 24936
rect 13722 24896 13728 24908
rect 13780 24896 13786 24948
rect 15470 24896 15476 24948
rect 15528 24936 15534 24948
rect 16025 24939 16083 24945
rect 16025 24936 16037 24939
rect 15528 24908 16037 24936
rect 15528 24896 15534 24908
rect 16025 24905 16037 24908
rect 16071 24905 16083 24939
rect 16025 24899 16083 24905
rect 5460 24840 5856 24868
rect 1854 24800 1860 24812
rect 1815 24772 1860 24800
rect 1854 24760 1860 24772
rect 1912 24760 1918 24812
rect 4706 24800 4712 24812
rect 4619 24772 4712 24800
rect 4706 24760 4712 24772
rect 4764 24800 4770 24812
rect 5460 24800 5488 24840
rect 4764 24772 5488 24800
rect 4764 24760 4770 24772
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 5828 24809 5856 24840
rect 6914 24828 6920 24880
rect 6972 24868 6978 24880
rect 7576 24868 7604 24896
rect 8021 24871 8079 24877
rect 8021 24868 8033 24871
rect 6972 24840 8033 24868
rect 6972 24828 6978 24840
rect 8021 24837 8033 24840
rect 8067 24837 8079 24871
rect 8021 24831 8079 24837
rect 5629 24803 5687 24809
rect 5629 24800 5641 24803
rect 5592 24772 5641 24800
rect 5592 24760 5598 24772
rect 5629 24769 5641 24772
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 1578 24732 1584 24744
rect 1539 24704 1584 24732
rect 1578 24692 1584 24704
rect 1636 24692 1642 24744
rect 2869 24735 2927 24741
rect 2869 24701 2881 24735
rect 2915 24732 2927 24735
rect 5828 24732 5856 24763
rect 7190 24760 7196 24812
rect 7248 24800 7254 24812
rect 7561 24803 7619 24809
rect 7561 24800 7573 24803
rect 7248 24772 7573 24800
rect 7248 24760 7254 24772
rect 7561 24769 7573 24772
rect 7607 24769 7619 24803
rect 10612 24800 10640 24896
rect 11241 24803 11299 24809
rect 11241 24800 11253 24803
rect 10612 24772 11253 24800
rect 7561 24763 7619 24769
rect 11241 24769 11253 24772
rect 11287 24769 11299 24803
rect 15488 24800 15516 24896
rect 11241 24763 11299 24769
rect 14200 24772 15516 24800
rect 14200 24744 14228 24772
rect 6270 24732 6276 24744
rect 2915 24704 3740 24732
rect 5828 24704 6276 24732
rect 2915 24701 2927 24704
rect 2869 24695 2927 24701
rect 3145 24667 3203 24673
rect 3145 24633 3157 24667
rect 3191 24664 3203 24667
rect 3510 24664 3516 24676
rect 3191 24636 3516 24664
rect 3191 24633 3203 24636
rect 3145 24627 3203 24633
rect 3510 24624 3516 24636
rect 3568 24624 3574 24676
rect 3712 24605 3740 24704
rect 6270 24692 6276 24704
rect 6328 24692 6334 24744
rect 6641 24735 6699 24741
rect 6641 24701 6653 24735
rect 6687 24732 6699 24735
rect 8570 24732 8576 24744
rect 6687 24704 7512 24732
rect 8531 24704 8576 24732
rect 6687 24701 6699 24704
rect 6641 24695 6699 24701
rect 4154 24664 4160 24676
rect 4067 24636 4160 24664
rect 4154 24624 4160 24636
rect 4212 24664 4218 24676
rect 4614 24664 4620 24676
rect 4212 24636 4620 24664
rect 4212 24624 4218 24636
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 7484 24673 7512 24704
rect 8570 24692 8576 24704
rect 8628 24732 8634 24744
rect 9125 24735 9183 24741
rect 9125 24732 9137 24735
rect 8628 24704 9137 24732
rect 8628 24692 8634 24704
rect 9125 24701 9137 24704
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 9858 24732 9864 24744
rect 9723 24704 9864 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9858 24692 9864 24704
rect 9916 24732 9922 24744
rect 10229 24735 10287 24741
rect 10229 24732 10241 24735
rect 9916 24704 10241 24732
rect 9916 24692 9922 24704
rect 10229 24701 10241 24704
rect 10275 24701 10287 24735
rect 10229 24695 10287 24701
rect 11057 24735 11115 24741
rect 11057 24701 11069 24735
rect 11103 24732 11115 24735
rect 11103 24704 11928 24732
rect 11103 24701 11115 24704
rect 11057 24695 11115 24701
rect 5077 24667 5135 24673
rect 5077 24633 5089 24667
rect 5123 24664 5135 24667
rect 7469 24667 7527 24673
rect 5123 24636 5580 24664
rect 5123 24633 5135 24636
rect 5077 24627 5135 24633
rect 5552 24608 5580 24636
rect 7469 24633 7481 24667
rect 7515 24664 7527 24667
rect 8846 24664 8852 24676
rect 7515 24636 8852 24664
rect 7515 24633 7527 24636
rect 7469 24627 7527 24633
rect 8846 24624 8852 24636
rect 8904 24624 8910 24676
rect 3697 24599 3755 24605
rect 3697 24565 3709 24599
rect 3743 24596 3755 24599
rect 4522 24596 4528 24608
rect 3743 24568 4528 24596
rect 3743 24565 3755 24568
rect 3697 24559 3755 24565
rect 4522 24556 4528 24568
rect 4580 24556 4586 24608
rect 5166 24596 5172 24608
rect 5127 24568 5172 24596
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 5534 24596 5540 24608
rect 5495 24568 5540 24596
rect 5534 24556 5540 24568
rect 5592 24556 5598 24608
rect 6273 24599 6331 24605
rect 6273 24565 6285 24599
rect 6319 24596 6331 24599
rect 7377 24599 7435 24605
rect 7377 24596 7389 24599
rect 6319 24568 7389 24596
rect 6319 24565 6331 24568
rect 6273 24559 6331 24565
rect 7377 24565 7389 24568
rect 7423 24596 7435 24599
rect 7558 24596 7564 24608
rect 7423 24568 7564 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 7558 24556 7564 24568
rect 7616 24556 7622 24608
rect 8386 24596 8392 24608
rect 8347 24568 8392 24596
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 8754 24596 8760 24608
rect 8715 24568 8760 24596
rect 8754 24556 8760 24568
rect 8812 24556 8818 24608
rect 9858 24596 9864 24608
rect 9819 24568 9864 24596
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 11900 24605 11928 24704
rect 12158 24692 12164 24744
rect 12216 24732 12222 24744
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 12216 24704 12449 24732
rect 12216 24692 12222 24704
rect 12437 24701 12449 24704
rect 12483 24732 12495 24735
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12483 24704 13001 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 12989 24701 13001 24704
rect 13035 24701 13047 24735
rect 13538 24732 13544 24744
rect 13499 24704 13544 24732
rect 12989 24695 13047 24701
rect 13538 24692 13544 24704
rect 13596 24692 13602 24744
rect 14182 24692 14188 24744
rect 14240 24692 14246 24744
rect 15473 24735 15531 24741
rect 15473 24701 15485 24735
rect 15519 24732 15531 24735
rect 16853 24735 16911 24741
rect 15519 24704 15553 24732
rect 15519 24701 15531 24704
rect 15473 24695 15531 24701
rect 16853 24701 16865 24735
rect 16899 24732 16911 24735
rect 16899 24704 17540 24732
rect 16899 24701 16911 24704
rect 16853 24695 16911 24701
rect 15381 24667 15439 24673
rect 15381 24633 15393 24667
rect 15427 24664 15439 24667
rect 15488 24664 15516 24695
rect 15930 24664 15936 24676
rect 15427 24636 15936 24664
rect 15427 24633 15439 24636
rect 15381 24627 15439 24633
rect 15930 24624 15936 24636
rect 15988 24624 15994 24676
rect 11885 24599 11943 24605
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 12066 24596 12072 24608
rect 11931 24568 12072 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 12066 24556 12072 24568
rect 12124 24556 12130 24608
rect 13630 24556 13636 24608
rect 13688 24596 13694 24608
rect 14090 24596 14096 24608
rect 13688 24568 14096 24596
rect 13688 24556 13694 24568
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 15654 24596 15660 24608
rect 15615 24568 15660 24596
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 17034 24596 17040 24608
rect 16995 24568 17040 24596
rect 17034 24556 17040 24568
rect 17092 24556 17098 24608
rect 17512 24605 17540 24704
rect 17497 24599 17555 24605
rect 17497 24565 17509 24599
rect 17543 24596 17555 24599
rect 17770 24596 17776 24608
rect 17543 24568 17776 24596
rect 17543 24565 17555 24568
rect 17497 24559 17555 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 11238 24352 11244 24404
rect 11296 24392 11302 24404
rect 12253 24395 12311 24401
rect 12253 24392 12265 24395
rect 11296 24364 12265 24392
rect 11296 24352 11302 24364
rect 12253 24361 12265 24364
rect 12299 24361 12311 24395
rect 12253 24355 12311 24361
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16206 24392 16212 24404
rect 15519 24364 16212 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 17681 24395 17739 24401
rect 17681 24361 17693 24395
rect 17727 24392 17739 24395
rect 18506 24392 18512 24404
rect 17727 24364 18512 24392
rect 17727 24361 17739 24364
rect 17681 24355 17739 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 18782 24392 18788 24404
rect 18743 24364 18788 24392
rect 18782 24352 18788 24364
rect 18840 24352 18846 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19978 24392 19984 24404
rect 19935 24364 19984 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22002 24392 22008 24404
rect 21131 24364 22008 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 22186 24392 22192 24404
rect 22147 24364 22192 24392
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 4893 24327 4951 24333
rect 4893 24293 4905 24327
rect 4939 24324 4951 24327
rect 4982 24324 4988 24336
rect 4939 24296 4988 24324
rect 4939 24293 4951 24296
rect 4893 24287 4951 24293
rect 4982 24284 4988 24296
rect 5040 24284 5046 24336
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24225 1731 24259
rect 1946 24256 1952 24268
rect 1907 24228 1952 24256
rect 1673 24219 1731 24225
rect 1688 24188 1716 24219
rect 1946 24216 1952 24228
rect 2004 24216 2010 24268
rect 5258 24256 5264 24268
rect 5000 24228 5264 24256
rect 1688 24160 2544 24188
rect 2516 24061 2544 24160
rect 2866 24148 2872 24200
rect 2924 24188 2930 24200
rect 2961 24191 3019 24197
rect 2961 24188 2973 24191
rect 2924 24160 2973 24188
rect 2924 24148 2930 24160
rect 2961 24157 2973 24160
rect 3007 24157 3019 24191
rect 2961 24151 3019 24157
rect 4430 24148 4436 24200
rect 4488 24188 4494 24200
rect 5000 24197 5028 24228
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 7190 24265 7196 24268
rect 6825 24259 6883 24265
rect 6825 24225 6837 24259
rect 6871 24256 6883 24259
rect 7184 24256 7196 24265
rect 6871 24228 7196 24256
rect 6871 24225 6883 24228
rect 6825 24219 6883 24225
rect 7184 24219 7196 24228
rect 7190 24216 7196 24219
rect 7248 24216 7254 24268
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 10117 24259 10175 24265
rect 10117 24256 10129 24259
rect 10008 24228 10129 24256
rect 10008 24216 10014 24228
rect 10117 24225 10129 24228
rect 10163 24225 10175 24259
rect 10117 24219 10175 24225
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 12069 24259 12127 24265
rect 12069 24256 12081 24259
rect 11112 24228 12081 24256
rect 11112 24216 11118 24228
rect 12069 24225 12081 24228
rect 12115 24225 12127 24259
rect 12069 24219 12127 24225
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 13541 24259 13599 24265
rect 13541 24256 13553 24259
rect 13504 24228 13553 24256
rect 13504 24216 13510 24228
rect 13541 24225 13553 24228
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 13817 24259 13875 24265
rect 13817 24225 13829 24259
rect 13863 24256 13875 24259
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 13863 24228 15301 24256
rect 13863 24225 13875 24228
rect 13817 24219 13875 24225
rect 15289 24225 15301 24228
rect 15335 24256 15347 24259
rect 15562 24256 15568 24268
rect 15335 24228 15568 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15562 24216 15568 24228
rect 15620 24216 15626 24268
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24256 16451 24259
rect 16666 24256 16672 24268
rect 16439 24228 16672 24256
rect 16439 24225 16451 24228
rect 16393 24219 16451 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 18138 24216 18144 24268
rect 18196 24256 18202 24268
rect 18601 24259 18659 24265
rect 18601 24256 18613 24259
rect 18196 24228 18613 24256
rect 18196 24216 18202 24228
rect 18601 24225 18613 24228
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 20070 24256 20076 24268
rect 19751 24228 20076 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 20070 24216 20076 24228
rect 20128 24216 20134 24268
rect 20898 24256 20904 24268
rect 20859 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 22002 24256 22008 24268
rect 21963 24228 22008 24256
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4488 24160 4997 24188
rect 4488 24148 4494 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5077 24151 5135 24157
rect 6917 24191 6975 24197
rect 6917 24157 6929 24191
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 4525 24123 4583 24129
rect 4525 24120 4537 24123
rect 3476 24092 4537 24120
rect 3476 24080 3482 24092
rect 4525 24089 4537 24092
rect 4571 24089 4583 24123
rect 5092 24120 5120 24151
rect 5442 24120 5448 24132
rect 4525 24083 4583 24089
rect 5000 24092 5448 24120
rect 2501 24055 2559 24061
rect 2501 24021 2513 24055
rect 2547 24052 2559 24055
rect 3326 24052 3332 24064
rect 2547 24024 3332 24052
rect 2547 24021 2559 24024
rect 2501 24015 2559 24021
rect 3326 24012 3332 24024
rect 3384 24012 3390 24064
rect 4338 24052 4344 24064
rect 4299 24024 4344 24052
rect 4338 24012 4344 24024
rect 4396 24052 4402 24064
rect 5000 24052 5028 24092
rect 5442 24080 5448 24092
rect 5500 24080 5506 24132
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 6932 24120 6960 24151
rect 6696 24092 6960 24120
rect 6696 24080 6702 24092
rect 4396 24024 5028 24052
rect 5629 24055 5687 24061
rect 4396 24012 4402 24024
rect 5629 24021 5641 24055
rect 5675 24052 5687 24055
rect 6822 24052 6828 24064
rect 5675 24024 6828 24052
rect 5675 24021 5687 24024
rect 5629 24015 5687 24021
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 6932 24052 6960 24092
rect 7852 24092 8616 24120
rect 7282 24052 7288 24064
rect 6932 24024 7288 24052
rect 7282 24012 7288 24024
rect 7340 24052 7346 24064
rect 7852 24052 7880 24092
rect 8588 24064 8616 24092
rect 8294 24052 8300 24064
rect 7340 24024 7880 24052
rect 8255 24024 8300 24052
rect 7340 24012 7346 24024
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 8570 24052 8576 24064
rect 8531 24024 8576 24052
rect 8570 24012 8576 24024
rect 8628 24012 8634 24064
rect 9122 24052 9128 24064
rect 9035 24024 9128 24052
rect 9122 24012 9128 24024
rect 9180 24052 9186 24064
rect 9493 24055 9551 24061
rect 9493 24052 9505 24055
rect 9180 24024 9505 24052
rect 9180 24012 9186 24024
rect 9493 24021 9505 24024
rect 9539 24052 9551 24055
rect 9876 24052 9904 24151
rect 16577 24123 16635 24129
rect 16577 24089 16589 24123
rect 16623 24120 16635 24123
rect 17862 24120 17868 24132
rect 16623 24092 17868 24120
rect 16623 24089 16635 24092
rect 16577 24083 16635 24089
rect 17862 24080 17868 24092
rect 17920 24080 17926 24132
rect 10134 24052 10140 24064
rect 9539 24024 10140 24052
rect 9539 24021 9551 24024
rect 9493 24015 9551 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 11238 24052 11244 24064
rect 11199 24024 11244 24052
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 11609 24055 11667 24061
rect 11609 24021 11621 24055
rect 11655 24052 11667 24055
rect 11698 24052 11704 24064
rect 11655 24024 11704 24052
rect 11655 24021 11667 24024
rect 11609 24015 11667 24021
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 12710 24052 12716 24064
rect 12671 24024 12716 24052
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 13998 24012 14004 24064
rect 14056 24052 14062 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 14056 24024 14289 24052
rect 14056 24012 14062 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2406 23848 2412 23860
rect 2367 23820 2412 23848
rect 2406 23808 2412 23820
rect 2464 23808 2470 23860
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 4065 23851 4123 23857
rect 4065 23817 4077 23851
rect 4111 23848 4123 23851
rect 4890 23848 4896 23860
rect 4111 23820 4896 23848
rect 4111 23817 4123 23820
rect 4065 23811 4123 23817
rect 4890 23808 4896 23820
rect 4948 23808 4954 23860
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 5905 23851 5963 23857
rect 5905 23848 5917 23851
rect 5500 23820 5917 23848
rect 5500 23808 5506 23820
rect 5905 23817 5917 23820
rect 5951 23817 5963 23851
rect 6270 23848 6276 23860
rect 6231 23820 6276 23848
rect 5905 23811 5963 23817
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 6638 23848 6644 23860
rect 6599 23820 6644 23848
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12437 23851 12495 23857
rect 12437 23848 12449 23851
rect 12124 23820 12449 23848
rect 12124 23808 12130 23820
rect 12437 23817 12449 23820
rect 12483 23817 12495 23851
rect 12437 23811 12495 23817
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 15657 23851 15715 23857
rect 15657 23848 15669 23851
rect 15620 23820 15669 23848
rect 15620 23808 15626 23820
rect 15657 23817 15669 23820
rect 15703 23817 15715 23851
rect 15657 23811 15715 23817
rect 16393 23851 16451 23857
rect 16393 23817 16405 23851
rect 16439 23848 16451 23851
rect 16758 23848 16764 23860
rect 16439 23820 16764 23848
rect 16439 23817 16451 23820
rect 16393 23811 16451 23817
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19058 23848 19064 23860
rect 18279 23820 19064 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 19518 23848 19524 23860
rect 19383 23820 19524 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23382 23848 23388 23860
rect 22695 23820 23388 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 25314 23848 25320 23860
rect 23891 23820 25320 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 1581 23647 1639 23653
rect 1581 23613 1593 23647
rect 1627 23644 1639 23647
rect 2406 23644 2412 23656
rect 1627 23616 2412 23644
rect 1627 23613 1639 23616
rect 1581 23607 1639 23613
rect 2406 23604 2412 23616
rect 2464 23604 2470 23656
rect 2884 23644 2912 23808
rect 4430 23780 4436 23792
rect 4391 23752 4436 23780
rect 4430 23740 4436 23752
rect 4488 23740 4494 23792
rect 3510 23712 3516 23724
rect 3471 23684 3516 23712
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 5534 23672 5540 23724
rect 5592 23712 5598 23724
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 5592 23684 6837 23712
rect 5592 23672 5598 23684
rect 6825 23681 6837 23684
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7760 23684 7972 23712
rect 7760 23656 7788 23684
rect 3329 23647 3387 23653
rect 3329 23644 3341 23647
rect 2884 23616 3341 23644
rect 3329 23613 3341 23616
rect 3375 23613 3387 23647
rect 3329 23607 3387 23613
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3476 23616 3521 23644
rect 3476 23604 3482 23616
rect 4154 23604 4160 23656
rect 4212 23644 4218 23656
rect 4525 23647 4583 23653
rect 4525 23644 4537 23647
rect 4212 23616 4537 23644
rect 4212 23604 4218 23616
rect 4525 23613 4537 23616
rect 4571 23613 4583 23647
rect 7742 23644 7748 23656
rect 7703 23616 7748 23644
rect 4525 23607 4583 23613
rect 7742 23604 7748 23616
rect 7800 23604 7806 23656
rect 7837 23647 7895 23653
rect 7837 23613 7849 23647
rect 7883 23613 7895 23647
rect 7944 23644 7972 23684
rect 12710 23672 12716 23724
rect 12768 23712 12774 23724
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 12768 23684 12909 23712
rect 12768 23672 12774 23684
rect 12897 23681 12909 23684
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13722 23712 13728 23724
rect 13127 23684 13728 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 8093 23647 8151 23653
rect 8093 23644 8105 23647
rect 7944 23616 8105 23644
rect 7837 23607 7895 23613
rect 8093 23613 8105 23616
rect 8139 23613 8151 23647
rect 10134 23644 10140 23656
rect 10047 23616 10140 23644
rect 8093 23607 8151 23613
rect 1854 23576 1860 23588
rect 1815 23548 1860 23576
rect 1854 23536 1860 23548
rect 1912 23536 1918 23588
rect 4706 23536 4712 23588
rect 4764 23585 4770 23588
rect 4764 23579 4828 23585
rect 4764 23545 4782 23579
rect 4816 23545 4828 23579
rect 4764 23539 4828 23545
rect 4764 23536 4770 23539
rect 7190 23536 7196 23588
rect 7248 23576 7254 23588
rect 7377 23579 7435 23585
rect 7377 23576 7389 23579
rect 7248 23548 7389 23576
rect 7248 23536 7254 23548
rect 7377 23545 7389 23548
rect 7423 23576 7435 23579
rect 7852 23576 7880 23607
rect 10134 23604 10140 23616
rect 10192 23644 10198 23656
rect 11698 23644 11704 23656
rect 10192 23616 11704 23644
rect 10192 23604 10198 23616
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 11882 23644 11888 23656
rect 11795 23616 11888 23644
rect 11882 23604 11888 23616
rect 11940 23644 11946 23656
rect 13096 23644 13124 23675
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13998 23712 14004 23724
rect 13959 23684 14004 23712
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 20898 23712 20904 23724
rect 20859 23684 20904 23712
rect 20898 23672 20904 23684
rect 20956 23672 20962 23724
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 11940 23616 13124 23644
rect 16040 23616 16221 23644
rect 11940 23604 11946 23616
rect 8570 23576 8576 23588
rect 7423 23548 7788 23576
rect 7852 23548 8576 23576
rect 7423 23545 7435 23548
rect 7377 23539 7435 23545
rect 2682 23468 2688 23520
rect 2740 23508 2746 23520
rect 2961 23511 3019 23517
rect 2961 23508 2973 23511
rect 2740 23480 2973 23508
rect 2740 23468 2746 23480
rect 2961 23477 2973 23480
rect 3007 23477 3019 23511
rect 7760 23508 7788 23548
rect 8570 23536 8576 23548
rect 8628 23536 8634 23588
rect 9585 23579 9643 23585
rect 9585 23545 9597 23579
rect 9631 23576 9643 23579
rect 10382 23579 10440 23585
rect 10382 23576 10394 23579
rect 9631 23548 10394 23576
rect 9631 23545 9643 23548
rect 9585 23539 9643 23545
rect 10382 23545 10394 23548
rect 10428 23576 10440 23579
rect 10778 23576 10784 23588
rect 10428 23548 10784 23576
rect 10428 23545 10440 23548
rect 10382 23539 10440 23545
rect 10778 23536 10784 23548
rect 10836 23536 10842 23588
rect 12066 23536 12072 23588
rect 12124 23576 12130 23588
rect 13446 23576 13452 23588
rect 12124 23548 13452 23576
rect 12124 23536 12130 23548
rect 13446 23536 13452 23548
rect 13504 23536 13510 23588
rect 14246 23579 14304 23585
rect 14246 23576 14258 23579
rect 14016 23548 14258 23576
rect 14016 23520 14044 23548
rect 14246 23545 14258 23548
rect 14292 23545 14304 23579
rect 14246 23539 14304 23545
rect 16040 23520 16068 23616
rect 16209 23613 16221 23616
rect 16255 23613 16267 23647
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 16209 23607 16267 23613
rect 18046 23604 18052 23616
rect 18104 23644 18110 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18104 23616 18613 23644
rect 18104 23604 18110 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18601 23607 18659 23613
rect 19058 23604 19064 23656
rect 19116 23644 19122 23656
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 19116 23616 19165 23644
rect 19116 23604 19122 23616
rect 19153 23613 19165 23616
rect 19199 23644 19211 23647
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19199 23616 19717 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 20254 23644 20260 23656
rect 20215 23616 20260 23644
rect 19705 23607 19763 23613
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 21082 23604 21088 23656
rect 21140 23644 21146 23656
rect 21361 23647 21419 23653
rect 21361 23644 21373 23647
rect 21140 23616 21373 23644
rect 21140 23604 21146 23616
rect 21361 23613 21373 23616
rect 21407 23613 21419 23647
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 21361 23607 21419 23613
rect 22462 23604 22468 23616
rect 22520 23644 22526 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22520 23616 23029 23644
rect 22520 23604 22526 23616
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23532 23616 23673 23644
rect 23532 23604 23538 23616
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 18138 23536 18144 23588
rect 18196 23576 18202 23588
rect 18969 23579 19027 23585
rect 18969 23576 18981 23579
rect 18196 23548 18981 23576
rect 18196 23536 18202 23548
rect 18969 23545 18981 23548
rect 19015 23545 19027 23579
rect 18969 23539 19027 23545
rect 8202 23508 8208 23520
rect 7760 23480 8208 23508
rect 2961 23471 3019 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 9217 23511 9275 23517
rect 9217 23508 9229 23511
rect 8444 23480 9229 23508
rect 8444 23468 8450 23480
rect 9217 23477 9229 23480
rect 9263 23477 9275 23511
rect 9950 23508 9956 23520
rect 9911 23480 9956 23508
rect 9217 23471 9275 23477
rect 9950 23468 9956 23480
rect 10008 23508 10014 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 10008 23480 11529 23508
rect 10008 23468 10014 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 12253 23511 12311 23517
rect 12253 23477 12265 23511
rect 12299 23508 12311 23511
rect 12805 23511 12863 23517
rect 12805 23508 12817 23511
rect 12299 23480 12817 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 12805 23477 12817 23480
rect 12851 23508 12863 23511
rect 12894 23508 12900 23520
rect 12851 23480 12900 23508
rect 12851 23477 12863 23480
rect 12805 23471 12863 23477
rect 12894 23468 12900 23480
rect 12952 23468 12958 23520
rect 13909 23511 13967 23517
rect 13909 23477 13921 23511
rect 13955 23508 13967 23511
rect 13998 23508 14004 23520
rect 13955 23480 14004 23508
rect 13955 23477 13967 23480
rect 13909 23471 13967 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15378 23508 15384 23520
rect 15339 23480 15384 23508
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 16022 23508 16028 23520
rect 15983 23480 16028 23508
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 16666 23468 16672 23520
rect 16724 23508 16730 23520
rect 16761 23511 16819 23517
rect 16761 23508 16773 23511
rect 16724 23480 16773 23508
rect 16724 23468 16730 23480
rect 16761 23477 16773 23480
rect 16807 23477 16819 23511
rect 17494 23508 17500 23520
rect 17455 23480 17500 23508
rect 16761 23471 16819 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 20070 23508 20076 23520
rect 20031 23480 20076 23508
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 22002 23508 22008 23520
rect 21963 23480 22008 23508
rect 22002 23468 22008 23480
rect 22060 23468 22066 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 3418 23304 3424 23316
rect 3379 23276 3424 23304
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 8665 23307 8723 23313
rect 8665 23304 8677 23307
rect 8352 23276 8677 23304
rect 8352 23264 8358 23276
rect 8665 23273 8677 23276
rect 8711 23273 8723 23307
rect 9122 23304 9128 23316
rect 9083 23276 9128 23304
rect 8665 23267 8723 23273
rect 9122 23264 9128 23276
rect 9180 23264 9186 23316
rect 10778 23304 10784 23316
rect 10739 23276 10784 23304
rect 10778 23264 10784 23276
rect 10836 23304 10842 23316
rect 12621 23307 12679 23313
rect 12621 23304 12633 23307
rect 10836 23276 12633 23304
rect 10836 23264 10842 23276
rect 12621 23273 12633 23276
rect 12667 23273 12679 23307
rect 12621 23267 12679 23273
rect 12710 23264 12716 23316
rect 12768 23304 12774 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 12768 23276 13461 23304
rect 12768 23264 12774 23276
rect 13449 23273 13461 23276
rect 13495 23273 13507 23307
rect 13449 23267 13507 23273
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 14090 23304 14096 23316
rect 13780 23276 14096 23304
rect 13780 23264 13786 23276
rect 14090 23264 14096 23276
rect 14148 23304 14154 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 14148 23276 14473 23304
rect 14148 23264 14154 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 19337 23307 19395 23313
rect 19337 23273 19349 23307
rect 19383 23304 19395 23307
rect 20622 23304 20628 23316
rect 19383 23276 20628 23304
rect 19383 23273 19395 23276
rect 19337 23267 19395 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 2041 23239 2099 23245
rect 2041 23205 2053 23239
rect 2087 23236 2099 23239
rect 3234 23236 3240 23248
rect 2087 23208 3240 23236
rect 2087 23205 2099 23208
rect 2041 23199 2099 23205
rect 3234 23196 3240 23208
rect 3292 23196 3298 23248
rect 11508 23239 11566 23245
rect 11508 23205 11520 23239
rect 11554 23236 11566 23239
rect 11882 23236 11888 23248
rect 11554 23208 11888 23236
rect 11554 23205 11566 23208
rect 11508 23199 11566 23205
rect 11882 23196 11888 23208
rect 11940 23196 11946 23248
rect 13817 23239 13875 23245
rect 13817 23205 13829 23239
rect 13863 23236 13875 23239
rect 13906 23236 13912 23248
rect 13863 23208 13912 23236
rect 13863 23205 13875 23208
rect 13817 23199 13875 23205
rect 13906 23196 13912 23208
rect 13964 23196 13970 23248
rect 16577 23239 16635 23245
rect 16577 23205 16589 23239
rect 16623 23236 16635 23239
rect 17494 23236 17500 23248
rect 16623 23208 17500 23236
rect 16623 23205 16635 23208
rect 16577 23199 16635 23205
rect 17494 23196 17500 23208
rect 17552 23196 17558 23248
rect 22649 23239 22707 23245
rect 22649 23205 22661 23239
rect 22695 23236 22707 23239
rect 23382 23236 23388 23248
rect 22695 23208 23388 23236
rect 22695 23205 22707 23208
rect 22649 23199 22707 23205
rect 23382 23196 23388 23208
rect 23440 23196 23446 23248
rect 1762 23168 1768 23180
rect 1675 23140 1768 23168
rect 1762 23128 1768 23140
rect 1820 23168 1826 23180
rect 2682 23168 2688 23180
rect 1820 23140 2688 23168
rect 1820 23128 1826 23140
rect 2682 23128 2688 23140
rect 2740 23128 2746 23180
rect 4338 23177 4344 23180
rect 4332 23168 4344 23177
rect 4299 23140 4344 23168
rect 4332 23131 4344 23140
rect 4338 23128 4344 23131
rect 4396 23128 4402 23180
rect 7282 23168 7288 23180
rect 7243 23140 7288 23168
rect 7282 23128 7288 23140
rect 7340 23128 7346 23180
rect 7374 23128 7380 23180
rect 7432 23168 7438 23180
rect 7541 23171 7599 23177
rect 7541 23168 7553 23171
rect 7432 23140 7553 23168
rect 7432 23128 7438 23140
rect 7541 23137 7553 23140
rect 7587 23168 7599 23171
rect 8386 23168 8392 23180
rect 7587 23140 8392 23168
rect 7587 23137 7599 23140
rect 7541 23131 7599 23137
rect 8386 23128 8392 23140
rect 8444 23128 8450 23180
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23168 10103 23171
rect 10318 23168 10324 23180
rect 10091 23140 10324 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23168 11299 23171
rect 11790 23168 11796 23180
rect 11287 23140 11796 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 15102 23168 15108 23180
rect 13924 23140 15108 23168
rect 4062 23100 4068 23112
rect 3896 23072 4068 23100
rect 3896 22976 3924 23072
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 6270 23100 6276 23112
rect 6231 23072 6276 23100
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 10134 23100 10140 23112
rect 9539 23072 10140 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 9306 22992 9312 23044
rect 9364 23032 9370 23044
rect 9950 23032 9956 23044
rect 9364 23004 9956 23032
rect 9364 22992 9370 23004
rect 9950 22992 9956 23004
rect 10008 23032 10014 23044
rect 10244 23032 10272 23063
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 13924 23109 13952 23140
rect 15102 23128 15108 23140
rect 15160 23128 15166 23180
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 16298 23168 16304 23180
rect 16259 23140 16304 23168
rect 16298 23128 16304 23140
rect 16356 23128 16362 23180
rect 17862 23168 17868 23180
rect 17823 23140 17868 23168
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 19150 23168 19156 23180
rect 18187 23140 19156 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 19150 23128 19156 23140
rect 19208 23128 19214 23180
rect 22370 23168 22376 23180
rect 22331 23140 22376 23168
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 13909 23103 13967 23109
rect 13909 23100 13921 23103
rect 13596 23072 13921 23100
rect 13596 23060 13602 23072
rect 13909 23069 13921 23072
rect 13955 23069 13967 23103
rect 14090 23100 14096 23112
rect 14003 23072 14096 23100
rect 13909 23063 13967 23069
rect 14090 23060 14096 23072
rect 14148 23100 14154 23112
rect 15378 23100 15384 23112
rect 14148 23072 15384 23100
rect 14148 23060 14154 23072
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 10008 23004 10272 23032
rect 10008 22992 10014 23004
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 2406 22924 2412 22976
rect 2464 22964 2470 22976
rect 2501 22967 2559 22973
rect 2501 22964 2513 22967
rect 2464 22936 2513 22964
rect 2464 22924 2470 22936
rect 2501 22933 2513 22936
rect 2547 22933 2559 22967
rect 2501 22927 2559 22933
rect 3053 22967 3111 22973
rect 3053 22933 3065 22967
rect 3099 22964 3111 22967
rect 3510 22964 3516 22976
rect 3099 22936 3516 22964
rect 3099 22933 3111 22936
rect 3053 22927 3111 22933
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 3878 22964 3884 22976
rect 3839 22936 3884 22964
rect 3878 22924 3884 22936
rect 3936 22924 3942 22976
rect 5442 22964 5448 22976
rect 5403 22936 5448 22964
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 9490 22924 9496 22976
rect 9548 22964 9554 22976
rect 9677 22967 9735 22973
rect 9677 22964 9689 22967
rect 9548 22936 9689 22964
rect 9548 22924 9554 22936
rect 9677 22933 9689 22936
rect 9723 22933 9735 22967
rect 12894 22964 12900 22976
rect 12855 22936 12900 22964
rect 9677 22927 9735 22933
rect 12894 22924 12900 22936
rect 12952 22924 12958 22976
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 13265 22967 13323 22973
rect 13265 22964 13277 22967
rect 13136 22936 13277 22964
rect 13136 22924 13142 22936
rect 13265 22933 13277 22936
rect 13311 22933 13323 22967
rect 20254 22964 20260 22976
rect 20215 22936 20260 22964
rect 13265 22927 13323 22933
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 21361 22967 21419 22973
rect 21361 22964 21373 22967
rect 21140 22936 21373 22964
rect 21140 22924 21146 22936
rect 21361 22933 21373 22936
rect 21407 22933 21419 22967
rect 21361 22927 21419 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1673 22763 1731 22769
rect 1673 22729 1685 22763
rect 1719 22760 1731 22763
rect 1762 22760 1768 22772
rect 1719 22732 1768 22760
rect 1719 22729 1731 22732
rect 1673 22723 1731 22729
rect 1762 22720 1768 22732
rect 1820 22720 1826 22772
rect 2133 22763 2191 22769
rect 2133 22729 2145 22763
rect 2179 22760 2191 22763
rect 5534 22760 5540 22772
rect 2179 22732 5540 22760
rect 2179 22729 2191 22732
rect 2133 22723 2191 22729
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 5629 22763 5687 22769
rect 5629 22729 5641 22763
rect 5675 22760 5687 22763
rect 5997 22763 6055 22769
rect 5997 22760 6009 22763
rect 5675 22732 6009 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 5997 22729 6009 22732
rect 6043 22760 6055 22763
rect 6638 22760 6644 22772
rect 6043 22732 6644 22760
rect 6043 22729 6055 22732
rect 5997 22723 6055 22729
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 7374 22760 7380 22772
rect 7335 22732 7380 22760
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 7834 22760 7840 22772
rect 7795 22732 7840 22760
rect 7834 22720 7840 22732
rect 7892 22720 7898 22772
rect 8846 22760 8852 22772
rect 8807 22732 8852 22760
rect 8846 22720 8852 22732
rect 8904 22720 8910 22772
rect 9306 22760 9312 22772
rect 9267 22732 9312 22760
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 9950 22760 9956 22772
rect 9732 22732 9956 22760
rect 9732 22720 9738 22732
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 10781 22763 10839 22769
rect 10781 22760 10793 22763
rect 10192 22732 10793 22760
rect 10192 22720 10198 22732
rect 10781 22729 10793 22732
rect 10827 22729 10839 22763
rect 11882 22760 11888 22772
rect 11843 22732 11888 22760
rect 10781 22723 10839 22729
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 12158 22760 12164 22772
rect 12119 22732 12164 22760
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 13449 22763 13507 22769
rect 13449 22729 13461 22763
rect 13495 22760 13507 22763
rect 13538 22760 13544 22772
rect 13495 22732 13544 22760
rect 13495 22729 13507 22732
rect 13449 22723 13507 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 13872 22732 14933 22760
rect 13872 22720 13878 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 14921 22723 14979 22729
rect 15289 22763 15347 22769
rect 15289 22729 15301 22763
rect 15335 22760 15347 22763
rect 15378 22760 15384 22772
rect 15335 22732 15384 22760
rect 15335 22729 15347 22732
rect 15289 22723 15347 22729
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 19150 22760 19156 22772
rect 19111 22732 19156 22760
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 22370 22760 22376 22772
rect 22331 22732 22376 22760
rect 22370 22720 22376 22732
rect 22428 22720 22434 22772
rect 2406 22584 2412 22636
rect 2464 22624 2470 22636
rect 2593 22627 2651 22633
rect 2593 22624 2605 22627
rect 2464 22596 2605 22624
rect 2464 22584 2470 22596
rect 2593 22593 2605 22596
rect 2639 22593 2651 22627
rect 2593 22587 2651 22593
rect 2777 22627 2835 22633
rect 2777 22593 2789 22627
rect 2823 22624 2835 22627
rect 3234 22624 3240 22636
rect 2823 22596 3240 22624
rect 2823 22593 2835 22596
rect 2777 22587 2835 22593
rect 2041 22559 2099 22565
rect 2041 22525 2053 22559
rect 2087 22556 2099 22559
rect 2792 22556 2820 22587
rect 3234 22584 3240 22596
rect 3292 22584 3298 22636
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3568 22596 3801 22624
rect 3568 22584 3574 22596
rect 3789 22593 3801 22596
rect 3835 22624 3847 22627
rect 6825 22627 6883 22633
rect 3835 22596 4016 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 2087 22528 2820 22556
rect 2087 22525 2099 22528
rect 2041 22519 2099 22525
rect 3418 22516 3424 22568
rect 3476 22556 3482 22568
rect 3878 22556 3884 22568
rect 3476 22528 3884 22556
rect 3476 22516 3482 22528
rect 3878 22516 3884 22528
rect 3936 22516 3942 22568
rect 3988 22556 4016 22596
rect 6825 22593 6837 22627
rect 6871 22624 6883 22627
rect 6914 22624 6920 22636
rect 6871 22596 6920 22624
rect 6871 22593 6883 22596
rect 6825 22587 6883 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7745 22627 7803 22633
rect 7745 22593 7757 22627
rect 7791 22624 7803 22627
rect 8202 22624 8208 22636
rect 7791 22596 8208 22624
rect 7791 22593 7803 22596
rect 7745 22587 7803 22593
rect 8202 22584 8208 22596
rect 8260 22624 8266 22636
rect 8297 22627 8355 22633
rect 8297 22624 8309 22627
rect 8260 22596 8309 22624
rect 8260 22584 8266 22596
rect 8297 22593 8309 22596
rect 8343 22593 8355 22627
rect 8297 22587 8355 22593
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22624 8539 22627
rect 8864 22624 8892 22720
rect 10229 22695 10287 22701
rect 10229 22661 10241 22695
rect 10275 22692 10287 22695
rect 10318 22692 10324 22704
rect 10275 22664 10324 22692
rect 10275 22661 10287 22664
rect 10229 22655 10287 22661
rect 10318 22652 10324 22664
rect 10376 22652 10382 22704
rect 11054 22692 11060 22704
rect 10612 22664 11060 22692
rect 8527 22596 8892 22624
rect 9677 22627 9735 22633
rect 8527 22593 8539 22596
rect 8481 22587 8539 22593
rect 9677 22593 9689 22627
rect 9723 22624 9735 22627
rect 10612 22624 10640 22664
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 12618 22692 12624 22704
rect 12579 22664 12624 22692
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 9723 22596 10640 22624
rect 10689 22627 10747 22633
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11238 22624 11244 22636
rect 10735 22596 11244 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 11238 22584 11244 22596
rect 11296 22584 11302 22636
rect 11333 22627 11391 22633
rect 11333 22593 11345 22627
rect 11379 22593 11391 22627
rect 11333 22587 11391 22593
rect 4148 22559 4206 22565
rect 4148 22556 4160 22559
rect 3988 22528 4160 22556
rect 4148 22525 4160 22528
rect 4194 22556 4206 22559
rect 5442 22556 5448 22568
rect 4194 22528 5448 22556
rect 4194 22525 4206 22528
rect 4148 22519 4206 22525
rect 5442 22516 5448 22528
rect 5500 22516 5506 22568
rect 9401 22559 9459 22565
rect 9401 22525 9413 22559
rect 9447 22556 9459 22559
rect 9490 22556 9496 22568
rect 9447 22528 9496 22556
rect 9447 22525 9459 22528
rect 9401 22519 9459 22525
rect 9490 22516 9496 22528
rect 9548 22516 9554 22568
rect 10778 22516 10784 22568
rect 10836 22556 10842 22568
rect 11348 22556 11376 22587
rect 11698 22584 11704 22636
rect 11756 22624 11762 22636
rect 16022 22624 16028 22636
rect 11756 22596 13584 22624
rect 15983 22596 16028 22624
rect 11756 22584 11762 22596
rect 10836 22528 11376 22556
rect 10836 22516 10842 22528
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 13556 22565 13584 22596
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 12216 22528 12449 22556
rect 12216 22516 12222 22528
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 13541 22559 13599 22565
rect 13541 22525 13553 22559
rect 13587 22556 13599 22559
rect 13808 22559 13866 22565
rect 13587 22528 13676 22556
rect 13587 22525 13599 22528
rect 13541 22519 13599 22525
rect 1394 22448 1400 22500
rect 1452 22488 1458 22500
rect 2501 22491 2559 22497
rect 2501 22488 2513 22491
rect 1452 22460 2513 22488
rect 1452 22448 1458 22460
rect 2501 22457 2513 22460
rect 2547 22488 2559 22491
rect 3145 22491 3203 22497
rect 3145 22488 3157 22491
rect 2547 22460 3157 22488
rect 2547 22457 2559 22460
rect 2501 22451 2559 22457
rect 3145 22457 3157 22460
rect 3191 22457 3203 22491
rect 3145 22451 3203 22457
rect 13081 22491 13139 22497
rect 13081 22457 13093 22491
rect 13127 22488 13139 22491
rect 13648 22488 13676 22528
rect 13808 22525 13820 22559
rect 13854 22556 13866 22559
rect 14090 22556 14096 22568
rect 13854 22528 14096 22556
rect 13854 22525 13866 22528
rect 13808 22519 13866 22525
rect 14090 22516 14096 22528
rect 14148 22516 14154 22568
rect 15746 22556 15752 22568
rect 15659 22528 15752 22556
rect 15746 22516 15752 22528
rect 15804 22556 15810 22568
rect 16485 22559 16543 22565
rect 16485 22556 16497 22559
rect 15804 22528 16497 22556
rect 15804 22516 15810 22528
rect 16485 22525 16497 22528
rect 16531 22525 16543 22559
rect 16485 22519 16543 22525
rect 13722 22488 13728 22500
rect 13127 22460 13584 22488
rect 13648 22460 13728 22488
rect 13127 22457 13139 22460
rect 13081 22451 13139 22457
rect 5258 22420 5264 22432
rect 5219 22392 5264 22420
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 8202 22420 8208 22432
rect 8163 22392 8208 22420
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 10870 22380 10876 22432
rect 10928 22420 10934 22432
rect 11149 22423 11207 22429
rect 11149 22420 11161 22423
rect 10928 22392 11161 22420
rect 10928 22380 10934 22392
rect 11149 22389 11161 22392
rect 11195 22389 11207 22423
rect 13556 22420 13584 22460
rect 13722 22448 13728 22460
rect 13780 22448 13786 22500
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 17862 22488 17868 22500
rect 15344 22460 17868 22488
rect 15344 22448 15350 22460
rect 17862 22448 17868 22460
rect 17920 22488 17926 22500
rect 18233 22491 18291 22497
rect 18233 22488 18245 22491
rect 17920 22460 18245 22488
rect 17920 22448 17926 22460
rect 18233 22457 18245 22460
rect 18279 22457 18291 22491
rect 18233 22451 18291 22457
rect 13906 22420 13912 22432
rect 13556 22392 13912 22420
rect 11149 22383 11207 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 16022 22380 16028 22432
rect 16080 22420 16086 22432
rect 16298 22420 16304 22432
rect 16080 22392 16304 22420
rect 16080 22380 16086 22392
rect 16298 22380 16304 22392
rect 16356 22420 16362 22432
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16356 22392 16865 22420
rect 16356 22380 16362 22392
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 4338 22216 4344 22228
rect 4299 22188 4344 22216
rect 4338 22176 4344 22188
rect 4396 22176 4402 22228
rect 9125 22219 9183 22225
rect 9125 22185 9137 22219
rect 9171 22216 9183 22219
rect 9490 22216 9496 22228
rect 9171 22188 9496 22216
rect 9171 22185 9183 22188
rect 9125 22179 9183 22185
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 13354 22176 13360 22228
rect 13412 22216 13418 22228
rect 13722 22216 13728 22228
rect 13412 22188 13728 22216
rect 13412 22176 13418 22188
rect 13722 22176 13728 22188
rect 13780 22216 13786 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 13780 22188 14657 22216
rect 13780 22176 13786 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 14645 22179 14703 22185
rect 2777 22151 2835 22157
rect 2777 22117 2789 22151
rect 2823 22148 2835 22151
rect 2866 22148 2872 22160
rect 2823 22120 2872 22148
rect 2823 22117 2835 22120
rect 2777 22111 2835 22117
rect 2866 22108 2872 22120
rect 2924 22108 2930 22160
rect 3050 22108 3056 22160
rect 3108 22108 3114 22160
rect 5068 22151 5126 22157
rect 5068 22117 5080 22151
rect 5114 22148 5126 22151
rect 5258 22148 5264 22160
rect 5114 22120 5264 22148
rect 5114 22117 5126 22120
rect 5068 22111 5126 22117
rect 5258 22108 5264 22120
rect 5316 22108 5322 22160
rect 6270 22148 6276 22160
rect 5552 22120 6276 22148
rect 3068 22080 3096 22108
rect 2884 22052 3096 22080
rect 2498 21972 2504 22024
rect 2556 22012 2562 22024
rect 2884 22021 2912 22052
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 5552 22080 5580 22120
rect 6270 22108 6276 22120
rect 6328 22108 6334 22160
rect 7006 22148 7012 22160
rect 6967 22120 7012 22148
rect 7006 22108 7012 22120
rect 7064 22108 7070 22160
rect 8389 22151 8447 22157
rect 8389 22148 8401 22151
rect 8220 22120 8401 22148
rect 4212 22052 5580 22080
rect 4212 22040 4218 22052
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7466 22080 7472 22092
rect 7156 22052 7472 22080
rect 7156 22040 7162 22052
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 7742 22040 7748 22092
rect 7800 22080 7806 22092
rect 8220 22080 8248 22120
rect 8389 22117 8401 22120
rect 8435 22117 8447 22151
rect 14001 22151 14059 22157
rect 14001 22148 14013 22151
rect 8389 22111 8447 22117
rect 13832 22120 14013 22148
rect 7800 22052 8248 22080
rect 7800 22040 7806 22052
rect 9858 22040 9864 22092
rect 9916 22080 9922 22092
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 9916 22052 10057 22080
rect 9916 22040 9922 22052
rect 10045 22049 10057 22052
rect 10091 22049 10103 22083
rect 10045 22043 10103 22049
rect 11422 22040 11428 22092
rect 11480 22080 11486 22092
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 11480 22052 11713 22080
rect 11480 22040 11486 22052
rect 11701 22049 11713 22052
rect 11747 22049 11759 22083
rect 12526 22080 12532 22092
rect 12487 22052 12532 22080
rect 11701 22043 11759 22049
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13722 22080 13728 22092
rect 13587 22052 13728 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2556 21984 2881 22012
rect 2556 21972 2562 21984
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 3050 22012 3056 22024
rect 3011 21984 3056 22012
rect 2869 21975 2927 21981
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 3418 21972 3424 22024
rect 3476 22012 3482 22024
rect 3513 22015 3571 22021
rect 3513 22012 3525 22015
rect 3476 21984 3525 22012
rect 3476 21972 3482 21984
rect 3513 21981 3525 21984
rect 3559 22012 3571 22015
rect 4709 22015 4767 22021
rect 4709 22012 4721 22015
rect 3559 21984 4721 22012
rect 3559 21981 3571 21984
rect 3513 21975 3571 21981
rect 4709 21981 4721 21984
rect 4755 22012 4767 22015
rect 4798 22012 4804 22024
rect 4755 21984 4804 22012
rect 4755 21981 4767 21984
rect 4709 21975 4767 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 21981 8539 22015
rect 8481 21975 8539 21981
rect 1673 21947 1731 21953
rect 1673 21913 1685 21947
rect 1719 21944 1731 21947
rect 1854 21944 1860 21956
rect 1719 21916 1860 21944
rect 1719 21913 1731 21916
rect 1673 21907 1731 21913
rect 1854 21904 1860 21916
rect 1912 21904 1918 21956
rect 2409 21947 2467 21953
rect 2409 21913 2421 21947
rect 2455 21944 2467 21947
rect 3789 21947 3847 21953
rect 3789 21944 3801 21947
rect 2455 21916 3801 21944
rect 2455 21913 2467 21916
rect 2409 21907 2467 21913
rect 3789 21913 3801 21916
rect 3835 21944 3847 21947
rect 4246 21944 4252 21956
rect 3835 21916 4252 21944
rect 3835 21913 3847 21916
rect 3789 21907 3847 21913
rect 4246 21904 4252 21916
rect 4304 21904 4310 21956
rect 7282 21904 7288 21956
rect 7340 21944 7346 21956
rect 7837 21947 7895 21953
rect 7837 21944 7849 21947
rect 7340 21916 7849 21944
rect 7340 21904 7346 21916
rect 7837 21913 7849 21916
rect 7883 21944 7895 21947
rect 8202 21944 8208 21956
rect 7883 21916 8208 21944
rect 7883 21913 7895 21916
rect 7837 21907 7895 21913
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 8496 21944 8524 21975
rect 8570 21972 8576 22024
rect 8628 22012 8634 22024
rect 10134 22012 10140 22024
rect 8628 21984 8673 22012
rect 10095 21984 10140 22012
rect 8628 21972 8634 21984
rect 10134 21972 10140 21984
rect 10192 21972 10198 22024
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 11790 22012 11796 22024
rect 11751 21984 11796 22012
rect 10229 21975 10287 21981
rect 8754 21944 8760 21956
rect 8496 21916 8760 21944
rect 8754 21904 8760 21916
rect 8812 21944 8818 21956
rect 9677 21947 9735 21953
rect 9677 21944 9689 21947
rect 8812 21916 9689 21944
rect 8812 21904 8818 21916
rect 9677 21913 9689 21916
rect 9723 21913 9735 21947
rect 9677 21907 9735 21913
rect 1946 21876 1952 21888
rect 1907 21848 1952 21876
rect 1946 21836 1952 21848
rect 2004 21836 2010 21888
rect 6178 21876 6184 21888
rect 6139 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 6546 21876 6552 21888
rect 6507 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21876 6610 21888
rect 6822 21876 6828 21888
rect 6604 21848 6828 21876
rect 6604 21836 6610 21848
rect 6822 21836 6828 21848
rect 6880 21836 6886 21888
rect 7561 21879 7619 21885
rect 7561 21845 7573 21879
rect 7607 21876 7619 21879
rect 7742 21876 7748 21888
rect 7607 21848 7748 21876
rect 7607 21845 7619 21848
rect 7561 21839 7619 21845
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 8018 21876 8024 21888
rect 7979 21848 8024 21876
rect 8018 21836 8024 21848
rect 8076 21836 8082 21888
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 9493 21879 9551 21885
rect 9493 21876 9505 21879
rect 8444 21848 9505 21876
rect 8444 21836 8450 21848
rect 9493 21845 9505 21848
rect 9539 21876 9551 21879
rect 10244 21876 10272 21975
rect 11790 21972 11796 21984
rect 11848 21972 11854 22024
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 13173 22015 13231 22021
rect 11940 21984 11985 22012
rect 11940 21972 11946 21984
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13446 22012 13452 22024
rect 13219 21984 13452 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 13446 21972 13452 21984
rect 13504 22012 13510 22024
rect 13832 22012 13860 22120
rect 14001 22117 14013 22120
rect 14047 22117 14059 22151
rect 14001 22111 14059 22117
rect 14660 22080 14688 22179
rect 15562 22089 15568 22092
rect 15289 22083 15347 22089
rect 15289 22080 15301 22083
rect 14660 22052 15301 22080
rect 15289 22049 15301 22052
rect 15335 22049 15347 22083
rect 15556 22080 15568 22089
rect 15523 22052 15568 22080
rect 15289 22043 15347 22049
rect 15556 22043 15568 22052
rect 15562 22040 15568 22043
rect 15620 22040 15626 22092
rect 14090 22012 14096 22024
rect 13504 21984 13860 22012
rect 14051 21984 14096 22012
rect 13504 21972 13510 21984
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14323 21984 14504 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 11238 21944 11244 21956
rect 11199 21916 11244 21944
rect 11238 21904 11244 21916
rect 11296 21904 11302 21956
rect 13998 21904 14004 21956
rect 14056 21944 14062 21956
rect 14476 21944 14504 21984
rect 14056 21916 14504 21944
rect 14056 21904 14062 21916
rect 10870 21876 10876 21888
rect 9539 21848 10272 21876
rect 10831 21848 10876 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 11330 21876 11336 21888
rect 11291 21848 11336 21876
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 13630 21876 13636 21888
rect 13591 21848 13636 21876
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 14476 21876 14504 21916
rect 16669 21879 16727 21885
rect 16669 21876 16681 21879
rect 14476 21848 16681 21876
rect 16669 21845 16681 21848
rect 16715 21845 16727 21879
rect 16669 21839 16727 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1394 21672 1400 21684
rect 1355 21644 1400 21672
rect 1394 21632 1400 21644
rect 1452 21632 1458 21684
rect 2498 21672 2504 21684
rect 2459 21644 2504 21672
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 3050 21632 3056 21684
rect 3108 21672 3114 21684
rect 3237 21675 3295 21681
rect 3237 21672 3249 21675
rect 3108 21644 3249 21672
rect 3108 21632 3114 21644
rect 3237 21641 3249 21644
rect 3283 21672 3295 21675
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 3283 21644 4905 21672
rect 3283 21641 3295 21644
rect 3237 21635 3295 21641
rect 4893 21641 4905 21644
rect 4939 21672 4951 21675
rect 5258 21672 5264 21684
rect 4939 21644 5264 21672
rect 4939 21641 4951 21644
rect 4893 21635 4951 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 8478 21672 8484 21684
rect 8067 21644 8484 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8478 21632 8484 21644
rect 8536 21672 8542 21684
rect 9490 21672 9496 21684
rect 8536 21644 9496 21672
rect 8536 21632 8542 21644
rect 9490 21632 9496 21644
rect 9548 21632 9554 21684
rect 9950 21632 9956 21684
rect 10008 21672 10014 21684
rect 10321 21675 10379 21681
rect 10321 21672 10333 21675
rect 10008 21644 10333 21672
rect 10008 21632 10014 21644
rect 10321 21641 10333 21644
rect 10367 21641 10379 21675
rect 10321 21635 10379 21641
rect 11698 21632 11704 21684
rect 11756 21672 11762 21684
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 11756 21644 11897 21672
rect 11756 21632 11762 21644
rect 11885 21641 11897 21644
rect 11931 21641 11943 21675
rect 11885 21635 11943 21641
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 12216 21644 12633 21672
rect 12216 21632 12222 21644
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 13265 21675 13323 21681
rect 13265 21641 13277 21675
rect 13311 21672 13323 21675
rect 13998 21672 14004 21684
rect 13311 21644 14004 21672
rect 13311 21641 13323 21644
rect 13265 21635 13323 21641
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 14148 21644 15945 21672
rect 14148 21632 14154 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 3697 21607 3755 21613
rect 3697 21573 3709 21607
rect 3743 21604 3755 21607
rect 6178 21604 6184 21616
rect 3743 21576 6184 21604
rect 3743 21573 3755 21576
rect 3697 21567 3755 21573
rect 1854 21496 1860 21548
rect 1912 21536 1918 21548
rect 1949 21539 2007 21545
rect 1949 21536 1961 21539
rect 1912 21508 1961 21536
rect 1912 21496 1918 21508
rect 1949 21505 1961 21508
rect 1995 21505 2007 21539
rect 4246 21536 4252 21548
rect 4207 21508 4252 21536
rect 1949 21499 2007 21505
rect 1670 21428 1676 21480
rect 1728 21468 1734 21480
rect 1765 21471 1823 21477
rect 1765 21468 1777 21471
rect 1728 21440 1777 21468
rect 1728 21428 1734 21440
rect 1765 21437 1777 21440
rect 1811 21437 1823 21471
rect 1964 21468 1992 21499
rect 4246 21496 4252 21508
rect 4304 21496 4310 21548
rect 4448 21545 4476 21576
rect 6178 21564 6184 21576
rect 6236 21564 6242 21616
rect 10226 21604 10232 21616
rect 10187 21576 10232 21604
rect 10226 21564 10232 21576
rect 10284 21564 10290 21616
rect 15105 21607 15163 21613
rect 15105 21573 15117 21607
rect 15151 21604 15163 21607
rect 15151 21576 15516 21604
rect 15151 21573 15163 21576
rect 15105 21567 15163 21573
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 4614 21496 4620 21548
rect 4672 21536 4678 21548
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 4672 21508 5549 21536
rect 4672 21496 4678 21508
rect 5537 21505 5549 21508
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 6914 21496 6920 21548
rect 6972 21536 6978 21548
rect 7009 21539 7067 21545
rect 7009 21536 7021 21539
rect 6972 21508 7021 21536
rect 6972 21496 6978 21508
rect 7009 21505 7021 21508
rect 7055 21505 7067 21539
rect 7009 21499 7067 21505
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21536 11023 21539
rect 11238 21536 11244 21548
rect 11011 21508 11244 21536
rect 11011 21505 11023 21508
rect 10965 21499 11023 21505
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 13078 21536 13084 21548
rect 12084 21508 13084 21536
rect 2406 21468 2412 21480
rect 1964 21440 2412 21468
rect 1765 21431 1823 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 4154 21468 4160 21480
rect 4115 21440 4160 21468
rect 4154 21428 4160 21440
rect 4212 21428 4218 21480
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5442 21468 5448 21480
rect 5399 21440 5448 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5442 21428 5448 21440
rect 5500 21468 5506 21480
rect 6089 21471 6147 21477
rect 6089 21468 6101 21471
rect 5500 21440 6101 21468
rect 5500 21428 5506 21440
rect 6089 21437 6101 21440
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6687 21440 6837 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 6825 21437 6837 21440
rect 6871 21468 6883 21471
rect 8018 21468 8024 21480
rect 6871 21440 8024 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 8113 21471 8171 21477
rect 8113 21437 8125 21471
rect 8159 21468 8171 21471
rect 8202 21468 8208 21480
rect 8159 21440 8208 21468
rect 8159 21437 8171 21440
rect 8113 21431 8171 21437
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 8386 21477 8392 21480
rect 8380 21468 8392 21477
rect 8312 21440 8392 21468
rect 1486 21360 1492 21412
rect 1544 21400 1550 21412
rect 2498 21400 2504 21412
rect 1544 21372 2504 21400
rect 1544 21360 1550 21372
rect 2498 21360 2504 21372
rect 2556 21360 2562 21412
rect 3326 21360 3332 21412
rect 3384 21400 3390 21412
rect 7653 21403 7711 21409
rect 3384 21372 3832 21400
rect 3384 21360 3390 21372
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 1857 21335 1915 21341
rect 1857 21332 1869 21335
rect 1452 21304 1869 21332
rect 1452 21292 1458 21304
rect 1857 21301 1869 21304
rect 1903 21332 1915 21335
rect 1946 21332 1952 21344
rect 1903 21304 1952 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 2866 21332 2872 21344
rect 2779 21304 2872 21332
rect 2866 21292 2872 21304
rect 2924 21332 2930 21344
rect 3694 21332 3700 21344
rect 2924 21304 3700 21332
rect 2924 21292 2930 21304
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 3804 21341 3832 21372
rect 7653 21369 7665 21403
rect 7699 21400 7711 21403
rect 7926 21400 7932 21412
rect 7699 21372 7932 21400
rect 7699 21369 7711 21372
rect 7653 21363 7711 21369
rect 7926 21360 7932 21372
rect 7984 21400 7990 21412
rect 8312 21400 8340 21440
rect 8380 21431 8392 21440
rect 8386 21428 8392 21431
rect 8444 21428 8450 21480
rect 10781 21471 10839 21477
rect 10781 21437 10793 21471
rect 10827 21468 10839 21471
rect 11330 21468 11336 21480
rect 10827 21440 11336 21468
rect 10827 21437 10839 21440
rect 10781 21431 10839 21437
rect 11330 21428 11336 21440
rect 11388 21428 11394 21480
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 12084 21477 12112 21508
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 13354 21496 13360 21548
rect 13412 21536 13418 21548
rect 13722 21536 13728 21548
rect 13412 21508 13728 21536
rect 13412 21496 13418 21508
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 15488 21545 15516 21576
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 15562 21536 15568 21548
rect 15519 21508 15568 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 15562 21496 15568 21508
rect 15620 21536 15626 21548
rect 16577 21539 16635 21545
rect 16577 21536 16589 21539
rect 15620 21508 16589 21536
rect 15620 21496 15626 21508
rect 16577 21505 16589 21508
rect 16623 21536 16635 21539
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16623 21508 16957 21536
rect 16623 21505 16635 21508
rect 16577 21499 16635 21505
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11664 21440 12081 21468
rect 11664 21428 11670 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 12069 21431 12127 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21468 12495 21471
rect 12526 21468 12532 21480
rect 12483 21440 12532 21468
rect 12483 21437 12495 21440
rect 12437 21431 12495 21437
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 16666 21468 16672 21480
rect 13740 21440 16672 21468
rect 7984 21372 8340 21400
rect 7984 21360 7990 21372
rect 12158 21360 12164 21412
rect 12216 21400 12222 21412
rect 13740 21400 13768 21440
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 13970 21403 14028 21409
rect 13970 21400 13982 21403
rect 12216 21372 13768 21400
rect 13832 21372 13982 21400
rect 12216 21360 12222 21372
rect 13832 21344 13860 21372
rect 13970 21369 13982 21372
rect 14016 21369 14028 21403
rect 13970 21363 14028 21369
rect 3789 21335 3847 21341
rect 3789 21301 3801 21335
rect 3835 21301 3847 21335
rect 3789 21295 3847 21301
rect 4798 21292 4804 21344
rect 4856 21332 4862 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 4856 21304 5273 21332
rect 4856 21292 4862 21304
rect 5261 21301 5273 21304
rect 5307 21332 5319 21335
rect 6546 21332 6552 21344
rect 5307 21304 6552 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 9950 21332 9956 21344
rect 9907 21304 9956 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10686 21332 10692 21344
rect 10647 21304 10692 21332
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 11422 21332 11428 21344
rect 11383 21304 11428 21332
rect 11422 21292 11428 21304
rect 11480 21292 11486 21344
rect 11790 21332 11796 21344
rect 11751 21304 11796 21332
rect 11790 21292 11796 21304
rect 11848 21292 11854 21344
rect 13633 21335 13691 21341
rect 13633 21301 13645 21335
rect 13679 21332 13691 21335
rect 13814 21332 13820 21344
rect 13679 21304 13820 21332
rect 13679 21301 13691 21304
rect 13633 21295 13691 21301
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 15749 21335 15807 21341
rect 15749 21332 15761 21335
rect 15712 21304 15761 21332
rect 15712 21292 15718 21304
rect 15749 21301 15761 21304
rect 15795 21332 15807 21335
rect 15930 21332 15936 21344
rect 15795 21304 15936 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 15930 21292 15936 21304
rect 15988 21332 15994 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 15988 21304 16313 21332
rect 15988 21292 15994 21304
rect 16301 21301 16313 21304
rect 16347 21301 16359 21335
rect 16301 21295 16359 21301
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 16448 21304 16493 21332
rect 16448 21292 16454 21304
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1397 21131 1455 21137
rect 1397 21097 1409 21131
rect 1443 21128 1455 21131
rect 1670 21128 1676 21140
rect 1443 21100 1676 21128
rect 1443 21097 1455 21100
rect 1397 21091 1455 21097
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 3881 21131 3939 21137
rect 3881 21097 3893 21131
rect 3927 21128 3939 21131
rect 4154 21128 4160 21140
rect 3927 21100 4160 21128
rect 3927 21097 3939 21100
rect 3881 21091 3939 21097
rect 4154 21088 4160 21100
rect 4212 21088 4218 21140
rect 4890 21128 4896 21140
rect 4851 21100 4896 21128
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 8386 21128 8392 21140
rect 8347 21100 8392 21128
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 8754 21128 8760 21140
rect 8715 21100 8760 21128
rect 8754 21088 8760 21100
rect 8812 21088 8818 21140
rect 9125 21131 9183 21137
rect 9125 21097 9137 21131
rect 9171 21128 9183 21131
rect 9674 21128 9680 21140
rect 9171 21100 9680 21128
rect 9171 21097 9183 21100
rect 9125 21091 9183 21097
rect 9674 21088 9680 21100
rect 9732 21128 9738 21140
rect 10686 21128 10692 21140
rect 9732 21100 10692 21128
rect 9732 21088 9738 21100
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 11054 21128 11060 21140
rect 10967 21100 11060 21128
rect 11054 21088 11060 21100
rect 11112 21128 11118 21140
rect 11112 21100 11192 21128
rect 11112 21088 11118 21100
rect 4341 21063 4399 21069
rect 4341 21029 4353 21063
rect 4387 21060 4399 21063
rect 4430 21060 4436 21072
rect 4387 21032 4436 21060
rect 4387 21029 4399 21032
rect 4341 21023 4399 21029
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 1765 20995 1823 21001
rect 1765 20992 1777 20995
rect 1544 20964 1777 20992
rect 1544 20952 1550 20964
rect 1765 20961 1777 20964
rect 1811 20961 1823 20995
rect 1765 20955 1823 20961
rect 4065 20995 4123 21001
rect 4065 20961 4077 20995
rect 4111 20992 4123 20995
rect 4908 20992 4936 21088
rect 5905 21063 5963 21069
rect 5905 21029 5917 21063
rect 5951 21060 5963 21063
rect 5994 21060 6000 21072
rect 5951 21032 6000 21060
rect 5951 21029 5963 21032
rect 5905 21023 5963 21029
rect 5994 21020 6000 21032
rect 6052 21020 6058 21072
rect 7190 21020 7196 21072
rect 7248 21069 7254 21072
rect 7248 21063 7312 21069
rect 7248 21029 7266 21063
rect 7300 21029 7312 21063
rect 7248 21023 7312 21029
rect 7248 21020 7254 21023
rect 9490 21020 9496 21072
rect 9548 21060 9554 21072
rect 9858 21060 9864 21072
rect 9548 21032 9864 21060
rect 9548 21020 9554 21032
rect 9858 21020 9864 21032
rect 9916 21069 9922 21072
rect 9916 21063 9980 21069
rect 9916 21029 9934 21063
rect 9968 21029 9980 21063
rect 11164 21060 11192 21100
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 11701 21131 11759 21137
rect 11701 21128 11713 21131
rect 11388 21100 11713 21128
rect 11388 21088 11394 21100
rect 11701 21097 11713 21100
rect 11747 21097 11759 21131
rect 12066 21128 12072 21140
rect 12027 21100 12072 21128
rect 11701 21091 11759 21097
rect 12066 21088 12072 21100
rect 12124 21088 12130 21140
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 13504 21100 13645 21128
rect 13504 21088 13510 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 14645 21131 14703 21137
rect 14645 21128 14657 21131
rect 13780 21100 14657 21128
rect 13780 21088 13786 21100
rect 14645 21097 14657 21100
rect 14691 21128 14703 21131
rect 15013 21131 15071 21137
rect 15013 21128 15025 21131
rect 14691 21100 15025 21128
rect 14691 21097 14703 21100
rect 14645 21091 14703 21097
rect 15013 21097 15025 21100
rect 15059 21128 15071 21131
rect 15378 21128 15384 21140
rect 15059 21100 15384 21128
rect 15059 21097 15071 21100
rect 15013 21091 15071 21097
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 11425 21063 11483 21069
rect 11425 21060 11437 21063
rect 11164 21032 11437 21060
rect 9916 21023 9980 21029
rect 11425 21029 11437 21032
rect 11471 21060 11483 21063
rect 11882 21060 11888 21072
rect 11471 21032 11888 21060
rect 11471 21029 11483 21032
rect 11425 21023 11483 21029
rect 9916 21020 9922 21023
rect 11882 21020 11888 21032
rect 11940 21020 11946 21072
rect 13541 21063 13599 21069
rect 13541 21029 13553 21063
rect 13587 21060 13599 21063
rect 14090 21060 14096 21072
rect 13587 21032 14096 21060
rect 13587 21029 13599 21032
rect 13541 21023 13599 21029
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 4111 20964 4936 20992
rect 4111 20961 4123 20964
rect 4065 20955 4123 20961
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5592 20964 5825 20992
rect 5592 20952 5598 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 5813 20955 5871 20961
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20992 6975 20995
rect 7098 20992 7104 21004
rect 6963 20964 7104 20992
rect 6963 20961 6975 20964
rect 6917 20955 6975 20961
rect 7098 20952 7104 20964
rect 7156 20952 7162 21004
rect 9398 20992 9404 21004
rect 9359 20964 9404 20992
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 10226 20992 10232 21004
rect 9723 20964 10232 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 14001 20995 14059 21001
rect 12492 20964 12537 20992
rect 12492 20952 12498 20964
rect 14001 20961 14013 20995
rect 14047 20992 14059 20995
rect 14047 20964 14596 20992
rect 14047 20961 14059 20964
rect 14001 20955 14059 20961
rect 14568 20936 14596 20964
rect 1854 20924 1860 20936
rect 1815 20896 1860 20924
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20893 2007 20927
rect 6086 20924 6092 20936
rect 6047 20896 6092 20924
rect 1949 20887 2007 20893
rect 1964 20788 1992 20887
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 2777 20859 2835 20865
rect 2777 20856 2789 20859
rect 2240 20828 2789 20856
rect 2038 20788 2044 20800
rect 1964 20760 2044 20788
rect 2038 20748 2044 20760
rect 2096 20788 2102 20800
rect 2240 20788 2268 20828
rect 2777 20825 2789 20828
rect 2823 20825 2835 20859
rect 2777 20819 2835 20825
rect 2096 20760 2268 20788
rect 2501 20791 2559 20797
rect 2096 20748 2102 20760
rect 2501 20757 2513 20791
rect 2547 20788 2559 20791
rect 2590 20788 2596 20800
rect 2547 20760 2596 20788
rect 2547 20757 2559 20760
rect 2501 20751 2559 20757
rect 2590 20748 2596 20760
rect 2648 20748 2654 20800
rect 3510 20788 3516 20800
rect 3471 20760 3516 20788
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 5261 20791 5319 20797
rect 5261 20757 5273 20791
rect 5307 20788 5319 20791
rect 5442 20788 5448 20800
rect 5307 20760 5448 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 6546 20788 6552 20800
rect 6459 20760 6552 20788
rect 6546 20748 6552 20760
rect 6604 20788 6610 20800
rect 6822 20788 6828 20800
rect 6604 20760 6828 20788
rect 6604 20748 6610 20760
rect 6822 20748 6828 20760
rect 6880 20788 6886 20800
rect 7024 20788 7052 20887
rect 8202 20816 8208 20868
rect 8260 20856 8266 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 8260 20828 9229 20856
rect 8260 20816 8266 20828
rect 9217 20825 9229 20828
rect 9263 20856 9275 20859
rect 9490 20856 9496 20868
rect 9263 20828 9496 20856
rect 9263 20825 9275 20828
rect 9217 20819 9275 20825
rect 9490 20816 9496 20828
rect 9548 20816 9554 20868
rect 8220 20788 8248 20816
rect 6880 20760 8248 20788
rect 12544 20788 12572 20887
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 13814 20924 13820 20936
rect 12676 20896 13820 20924
rect 12676 20884 12682 20896
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 14292 20856 14320 20887
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14608 20896 15301 20924
rect 14608 20884 14614 20896
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 16298 20924 16304 20936
rect 16259 20896 16304 20924
rect 15289 20887 15347 20893
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 15562 20856 15568 20868
rect 14292 20828 15568 20856
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 13170 20788 13176 20800
rect 12544 20760 13176 20788
rect 6880 20748 6886 20760
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 14734 20748 14740 20800
rect 14792 20788 14798 20800
rect 15933 20791 15991 20797
rect 15933 20788 15945 20791
rect 14792 20760 15945 20788
rect 14792 20748 14798 20760
rect 15933 20757 15945 20760
rect 15979 20788 15991 20791
rect 16390 20788 16396 20800
rect 15979 20760 16396 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16390 20748 16396 20760
rect 16448 20748 16454 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2498 20544 2504 20596
rect 2556 20584 2562 20596
rect 3234 20584 3240 20596
rect 2556 20556 3240 20584
rect 2556 20544 2562 20556
rect 3234 20544 3240 20556
rect 3292 20544 3298 20596
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 6273 20587 6331 20593
rect 6273 20584 6285 20587
rect 6144 20556 6285 20584
rect 6144 20544 6150 20556
rect 6273 20553 6285 20556
rect 6319 20584 6331 20587
rect 6641 20587 6699 20593
rect 6641 20584 6653 20587
rect 6319 20556 6653 20584
rect 6319 20553 6331 20556
rect 6273 20547 6331 20553
rect 6641 20553 6653 20556
rect 6687 20584 6699 20587
rect 7190 20584 7196 20596
rect 6687 20556 7196 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7190 20544 7196 20556
rect 7248 20584 7254 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7248 20556 8217 20584
rect 7248 20544 7254 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 9214 20584 9220 20596
rect 9175 20556 9220 20584
rect 8205 20547 8263 20553
rect 9214 20544 9220 20556
rect 9272 20544 9278 20596
rect 9769 20587 9827 20593
rect 9769 20553 9781 20587
rect 9815 20584 9827 20587
rect 9858 20584 9864 20596
rect 9815 20556 9864 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 12161 20587 12219 20593
rect 12161 20553 12173 20587
rect 12207 20584 12219 20587
rect 12618 20584 12624 20596
rect 12207 20556 12624 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 13814 20584 13820 20596
rect 13775 20556 13820 20584
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 14090 20584 14096 20596
rect 14051 20556 14096 20584
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14550 20584 14556 20596
rect 14511 20556 14556 20584
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 15562 20584 15568 20596
rect 15243 20556 15568 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 16025 20587 16083 20593
rect 16025 20553 16037 20587
rect 16071 20584 16083 20587
rect 16114 20584 16120 20596
rect 16071 20556 16120 20584
rect 16071 20553 16083 20556
rect 16025 20547 16083 20553
rect 16114 20544 16120 20556
rect 16172 20544 16178 20596
rect 8573 20519 8631 20525
rect 8573 20485 8585 20519
rect 8619 20516 8631 20519
rect 8754 20516 8760 20528
rect 8619 20488 8760 20516
rect 8619 20485 8631 20488
rect 8573 20479 8631 20485
rect 8754 20476 8760 20488
rect 8812 20516 8818 20528
rect 9398 20516 9404 20528
rect 8812 20488 9404 20516
rect 8812 20476 8818 20488
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 15378 20476 15384 20528
rect 15436 20516 15442 20528
rect 15473 20519 15531 20525
rect 15473 20516 15485 20519
rect 15436 20488 15485 20516
rect 15436 20476 15442 20488
rect 15473 20485 15485 20488
rect 15519 20485 15531 20519
rect 15473 20479 15531 20485
rect 1854 20448 1860 20460
rect 1596 20420 1860 20448
rect 1596 20256 1624 20420
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 3050 20448 3056 20460
rect 2731 20420 3056 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 3050 20408 3056 20420
rect 3108 20408 3114 20460
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 4154 20448 4160 20460
rect 3568 20420 4160 20448
rect 3568 20408 3574 20420
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 4709 20451 4767 20457
rect 4709 20417 4721 20451
rect 4755 20448 4767 20451
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 4755 20420 5825 20448
rect 4755 20417 4767 20420
rect 4709 20411 4767 20417
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 5859 20420 6960 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 4062 20380 4068 20392
rect 4023 20352 4068 20380
rect 4062 20340 4068 20352
rect 4120 20380 4126 20392
rect 4338 20380 4344 20392
rect 4120 20352 4344 20380
rect 4120 20340 4126 20352
rect 4338 20340 4344 20352
rect 4396 20340 4402 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5000 20352 5641 20380
rect 1946 20272 1952 20324
rect 2004 20312 2010 20324
rect 2501 20315 2559 20321
rect 2501 20312 2513 20315
rect 2004 20284 2513 20312
rect 2004 20272 2010 20284
rect 2501 20281 2513 20284
rect 2547 20281 2559 20315
rect 2501 20275 2559 20281
rect 3513 20315 3571 20321
rect 3513 20281 3525 20315
rect 3559 20312 3571 20315
rect 3559 20284 4016 20312
rect 3559 20281 3571 20284
rect 3513 20275 3571 20281
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 2041 20247 2099 20253
rect 2041 20244 2053 20247
rect 1820 20216 2053 20244
rect 1820 20204 1826 20216
rect 2041 20213 2053 20216
rect 2087 20213 2099 20247
rect 2041 20207 2099 20213
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 2590 20244 2596 20256
rect 2455 20216 2596 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 3050 20244 3056 20256
rect 3011 20216 3056 20244
rect 3050 20204 3056 20216
rect 3108 20204 3114 20256
rect 3602 20244 3608 20256
rect 3563 20216 3608 20244
rect 3602 20204 3608 20216
rect 3660 20204 3666 20256
rect 3988 20253 4016 20284
rect 3973 20247 4031 20253
rect 3973 20213 3985 20247
rect 4019 20244 4031 20247
rect 4246 20244 4252 20256
rect 4019 20216 4252 20244
rect 4019 20213 4031 20216
rect 3973 20207 4031 20213
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4430 20204 4436 20256
rect 4488 20244 4494 20256
rect 5000 20253 5028 20352
rect 5629 20349 5641 20352
rect 5675 20380 5687 20383
rect 6822 20380 6828 20392
rect 5675 20352 6684 20380
rect 6783 20352 6828 20380
rect 5675 20349 5687 20352
rect 5629 20343 5687 20349
rect 5442 20272 5448 20324
rect 5500 20312 5506 20324
rect 5537 20315 5595 20321
rect 5537 20312 5549 20315
rect 5500 20284 5549 20312
rect 5500 20272 5506 20284
rect 5537 20281 5549 20284
rect 5583 20312 5595 20315
rect 6086 20312 6092 20324
rect 5583 20284 6092 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 6086 20272 6092 20284
rect 6144 20272 6150 20324
rect 6656 20312 6684 20352
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 6932 20380 6960 20420
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 11756 20420 12449 20448
rect 11756 20408 11762 20420
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 14642 20448 14648 20460
rect 14603 20420 14648 20448
rect 12437 20411 12495 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 7098 20389 7104 20392
rect 7092 20380 7104 20389
rect 6932 20352 7104 20380
rect 7092 20343 7104 20352
rect 7098 20340 7104 20343
rect 7156 20340 7162 20392
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8956 20352 9045 20380
rect 7282 20312 7288 20324
rect 6656 20284 7288 20312
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 8956 20256 8984 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20380 10195 20383
rect 10226 20380 10232 20392
rect 10183 20352 10232 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 10226 20340 10232 20352
rect 10284 20380 10290 20392
rect 11716 20380 11744 20408
rect 15838 20380 15844 20392
rect 10284 20352 11744 20380
rect 15751 20352 15844 20380
rect 10284 20340 10290 20352
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16393 20383 16451 20389
rect 16393 20380 16405 20383
rect 15896 20352 16405 20380
rect 15896 20340 15902 20352
rect 16393 20349 16405 20352
rect 16439 20349 16451 20383
rect 16393 20343 16451 20349
rect 10404 20315 10462 20321
rect 10404 20281 10416 20315
rect 10450 20312 10462 20315
rect 11054 20312 11060 20324
rect 10450 20284 11060 20312
rect 10450 20281 10462 20284
rect 10404 20275 10462 20281
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 12704 20315 12762 20321
rect 12704 20281 12716 20315
rect 12750 20312 12762 20315
rect 13078 20312 13084 20324
rect 12750 20284 13084 20312
rect 12750 20281 12762 20284
rect 12704 20275 12762 20281
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 4985 20247 5043 20253
rect 4985 20244 4997 20247
rect 4488 20216 4997 20244
rect 4488 20204 4494 20216
rect 4985 20213 4997 20216
rect 5031 20213 5043 20247
rect 5166 20244 5172 20256
rect 5127 20216 5172 20244
rect 4985 20207 5043 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 8938 20244 8944 20256
rect 8899 20216 8944 20244
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11388 20216 11529 20244
rect 11388 20204 11394 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14182 20244 14188 20256
rect 13872 20216 14188 20244
rect 13872 20204 13878 20216
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2041 20043 2099 20049
rect 2041 20040 2053 20043
rect 2004 20012 2053 20040
rect 2004 20000 2010 20012
rect 2041 20009 2053 20012
rect 2087 20009 2099 20043
rect 2041 20003 2099 20009
rect 2682 20000 2688 20052
rect 2740 20040 2746 20052
rect 2869 20043 2927 20049
rect 2869 20040 2881 20043
rect 2740 20012 2881 20040
rect 2740 20000 2746 20012
rect 2869 20009 2881 20012
rect 2915 20009 2927 20043
rect 2869 20003 2927 20009
rect 3697 20043 3755 20049
rect 3697 20009 3709 20043
rect 3743 20040 3755 20043
rect 4062 20040 4068 20052
rect 3743 20012 4068 20040
rect 3743 20009 3755 20012
rect 3697 20003 3755 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 5813 20043 5871 20049
rect 5813 20009 5825 20043
rect 5859 20040 5871 20043
rect 5994 20040 6000 20052
rect 5859 20012 6000 20040
rect 5859 20009 5871 20012
rect 5813 20003 5871 20009
rect 5994 20000 6000 20012
rect 6052 20040 6058 20052
rect 6733 20043 6791 20049
rect 6733 20040 6745 20043
rect 6052 20012 6745 20040
rect 6052 20000 6058 20012
rect 6733 20009 6745 20012
rect 6779 20009 6791 20043
rect 6733 20003 6791 20009
rect 7193 20043 7251 20049
rect 7193 20009 7205 20043
rect 7239 20040 7251 20043
rect 7374 20040 7380 20052
rect 7239 20012 7380 20040
rect 7239 20009 7251 20012
rect 7193 20003 7251 20009
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 7926 20040 7932 20052
rect 7887 20012 7932 20040
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 9674 20040 9680 20052
rect 9635 20012 9680 20040
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10781 20043 10839 20049
rect 10781 20009 10793 20043
rect 10827 20040 10839 20043
rect 11054 20040 11060 20052
rect 10827 20012 11060 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 3878 19932 3884 19984
rect 3936 19972 3942 19984
rect 4154 19972 4160 19984
rect 3936 19944 4160 19972
rect 3936 19932 3942 19944
rect 4154 19932 4160 19944
rect 4212 19972 4218 19984
rect 4310 19975 4368 19981
rect 4310 19972 4322 19975
rect 4212 19944 4322 19972
rect 4212 19932 4218 19944
rect 4310 19941 4322 19944
rect 4356 19941 4368 19975
rect 4310 19935 4368 19941
rect 5166 19932 5172 19984
rect 5224 19972 5230 19984
rect 5534 19972 5540 19984
rect 5224 19944 5540 19972
rect 5224 19932 5230 19944
rect 5534 19932 5540 19944
rect 5592 19972 5598 19984
rect 6089 19975 6147 19981
rect 6089 19972 6101 19975
rect 5592 19944 6101 19972
rect 5592 19932 5598 19944
rect 6089 19941 6101 19944
rect 6135 19941 6147 19975
rect 6546 19972 6552 19984
rect 6507 19944 6552 19972
rect 6089 19935 6147 19941
rect 6546 19932 6552 19944
rect 6604 19932 6610 19984
rect 10137 19975 10195 19981
rect 10137 19941 10149 19975
rect 10183 19972 10195 19975
rect 10318 19972 10324 19984
rect 10183 19944 10324 19972
rect 10183 19941 10195 19944
rect 10137 19935 10195 19941
rect 10318 19932 10324 19944
rect 10376 19932 10382 19984
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3786 19904 3792 19916
rect 2823 19876 3792 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19904 7159 19907
rect 7650 19904 7656 19916
rect 7147 19876 7656 19904
rect 7147 19873 7159 19876
rect 7101 19867 7159 19873
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19904 8355 19907
rect 8386 19904 8392 19916
rect 8343 19876 8392 19904
rect 8343 19873 8355 19876
rect 8297 19867 8355 19873
rect 8386 19864 8392 19876
rect 8444 19904 8450 19916
rect 8849 19907 8907 19913
rect 8849 19904 8861 19907
rect 8444 19876 8861 19904
rect 8444 19864 8450 19876
rect 8849 19873 8861 19876
rect 8895 19873 8907 19907
rect 8849 19867 8907 19873
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10045 19907 10103 19913
rect 10045 19904 10057 19907
rect 9732 19876 10057 19904
rect 9732 19864 9738 19876
rect 10045 19873 10057 19876
rect 10091 19873 10103 19907
rect 10045 19867 10103 19873
rect 3050 19836 3056 19848
rect 2963 19808 3056 19836
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 4062 19836 4068 19848
rect 4023 19808 4068 19836
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 7285 19839 7343 19845
rect 7285 19836 7297 19839
rect 7248 19808 7297 19836
rect 7248 19796 7254 19808
rect 7285 19805 7297 19808
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10321 19839 10379 19845
rect 10321 19836 10333 19839
rect 10192 19808 10333 19836
rect 10192 19796 10198 19808
rect 10321 19805 10333 19808
rect 10367 19836 10379 19839
rect 10796 19836 10824 20003
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 13170 20000 13176 20052
rect 13228 20040 13234 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 13228 20012 13461 20040
rect 13228 20000 13234 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13814 20040 13820 20052
rect 13775 20012 13820 20040
rect 13449 20003 13507 20009
rect 13814 20000 13820 20012
rect 13872 20040 13878 20052
rect 13872 20012 14320 20040
rect 13872 20000 13878 20012
rect 14292 19984 14320 20012
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14608 20012 14933 20040
rect 14608 20000 14614 20012
rect 14921 20009 14933 20012
rect 14967 20040 14979 20043
rect 15378 20040 15384 20052
rect 14967 20012 15384 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 11698 19972 11704 19984
rect 11256 19944 11704 19972
rect 11256 19913 11284 19944
rect 11698 19932 11704 19944
rect 11756 19932 11762 19984
rect 12434 19932 12440 19984
rect 12492 19972 12498 19984
rect 13265 19975 13323 19981
rect 13265 19972 13277 19975
rect 12492 19944 13277 19972
rect 12492 19932 12498 19944
rect 13265 19941 13277 19944
rect 13311 19941 13323 19975
rect 13265 19935 13323 19941
rect 14274 19932 14280 19984
rect 14332 19932 14338 19984
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 11497 19907 11555 19913
rect 11497 19904 11509 19907
rect 11388 19876 11509 19904
rect 11388 19864 11394 19876
rect 11497 19873 11509 19876
rect 11543 19873 11555 19907
rect 11497 19867 11555 19873
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 15194 19904 15200 19916
rect 14148 19876 15200 19904
rect 14148 19864 14154 19876
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 15304 19913 15332 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15545 19907 15603 19913
rect 15545 19904 15557 19907
rect 15436 19876 15557 19904
rect 15436 19864 15442 19876
rect 15545 19873 15557 19876
rect 15591 19873 15603 19907
rect 15545 19867 15603 19873
rect 13906 19836 13912 19848
rect 10367 19808 10824 19836
rect 13867 19808 13912 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 13906 19796 13912 19808
rect 13964 19796 13970 19848
rect 14001 19839 14059 19845
rect 14001 19805 14013 19839
rect 14047 19805 14059 19839
rect 14001 19799 14059 19805
rect 3068 19768 3096 19796
rect 3970 19768 3976 19780
rect 3068 19740 3976 19768
rect 3970 19728 3976 19740
rect 4028 19728 4034 19780
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 8481 19771 8539 19777
rect 8481 19768 8493 19771
rect 5408 19740 8493 19768
rect 5408 19728 5414 19740
rect 8481 19737 8493 19740
rect 8527 19737 8539 19771
rect 8481 19731 8539 19737
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 10870 19768 10876 19780
rect 10744 19740 10876 19768
rect 10744 19728 10750 19740
rect 10870 19728 10876 19740
rect 10928 19768 10934 19780
rect 12621 19771 12679 19777
rect 10928 19740 11284 19768
rect 10928 19728 10934 19740
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 1581 19703 1639 19709
rect 1581 19700 1593 19703
rect 1544 19672 1593 19700
rect 1544 19660 1550 19672
rect 1581 19669 1593 19672
rect 1627 19669 1639 19703
rect 1581 19663 1639 19669
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 2409 19703 2467 19709
rect 2409 19700 2421 19703
rect 2188 19672 2421 19700
rect 2188 19660 2194 19672
rect 2409 19669 2421 19672
rect 2455 19669 2467 19703
rect 2409 19663 2467 19669
rect 5166 19660 5172 19712
rect 5224 19700 5230 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5224 19672 5457 19700
rect 5224 19660 5230 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 9398 19700 9404 19712
rect 9359 19672 9404 19700
rect 5445 19663 5503 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 11146 19700 11152 19712
rect 11107 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11256 19700 11284 19740
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 12989 19771 13047 19777
rect 12989 19768 13001 19771
rect 12667 19740 13001 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 12989 19737 13001 19740
rect 13035 19768 13047 19771
rect 13078 19768 13084 19780
rect 13035 19740 13084 19768
rect 13035 19737 13047 19740
rect 12989 19731 13047 19737
rect 13078 19728 13084 19740
rect 13136 19768 13142 19780
rect 14016 19768 14044 19799
rect 13136 19740 14044 19768
rect 13136 19728 13142 19740
rect 14458 19700 14464 19712
rect 11256 19672 14464 19700
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 3786 19496 3792 19508
rect 3747 19468 3792 19496
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 7190 19496 7196 19508
rect 6319 19468 7196 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 7650 19496 7656 19508
rect 7423 19468 7656 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 10965 19499 11023 19505
rect 10965 19465 10977 19499
rect 11011 19496 11023 19499
rect 11330 19496 11336 19508
rect 11011 19468 11336 19496
rect 11011 19465 11023 19468
rect 10965 19459 11023 19465
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12492 19468 12537 19496
rect 12492 19456 12498 19468
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 15528 19468 16681 19496
rect 15528 19456 15534 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 1302 19388 1308 19440
rect 1360 19428 1366 19440
rect 1578 19428 1584 19440
rect 1360 19400 1584 19428
rect 1360 19388 1366 19400
rect 1578 19388 1584 19400
rect 1636 19388 1642 19440
rect 3050 19388 3056 19440
rect 3108 19428 3114 19440
rect 4062 19428 4068 19440
rect 3108 19400 4068 19428
rect 3108 19388 3114 19400
rect 4062 19388 4068 19400
rect 4120 19388 4126 19440
rect 13906 19428 13912 19440
rect 13819 19400 13912 19428
rect 13906 19388 13912 19400
rect 13964 19428 13970 19440
rect 14366 19428 14372 19440
rect 13964 19400 14372 19428
rect 13964 19388 13970 19400
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 3234 19360 3240 19372
rect 2700 19332 3240 19360
rect 2700 19304 2728 19332
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 4080 19360 4108 19388
rect 3384 19332 3429 19360
rect 4080 19332 4200 19360
rect 3384 19320 3390 19332
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1578 19292 1584 19304
rect 1443 19264 1584 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2682 19252 2688 19304
rect 2740 19252 2746 19304
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19292 3111 19295
rect 3602 19292 3608 19304
rect 3099 19264 3608 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 3602 19252 3608 19264
rect 3660 19292 3666 19304
rect 4062 19292 4068 19304
rect 3660 19264 4068 19292
rect 3660 19252 3666 19264
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4172 19292 4200 19332
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6144 19332 6837 19360
rect 6144 19320 6150 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 7374 19360 7380 19372
rect 6825 19323 6883 19329
rect 6932 19332 7380 19360
rect 4249 19295 4307 19301
rect 4249 19292 4261 19295
rect 4172 19264 4261 19292
rect 4249 19261 4261 19264
rect 4295 19292 4307 19295
rect 6546 19292 6552 19304
rect 4295 19264 6552 19292
rect 4295 19261 4307 19264
rect 4249 19255 4307 19261
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6932 19292 6960 19332
rect 7374 19320 7380 19332
rect 7432 19360 7438 19372
rect 7834 19360 7840 19372
rect 7432 19332 7840 19360
rect 7432 19320 7438 19332
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 7926 19320 7932 19372
rect 7984 19360 7990 19372
rect 8389 19363 8447 19369
rect 8389 19360 8401 19363
rect 7984 19332 8401 19360
rect 7984 19320 7990 19332
rect 8389 19329 8401 19332
rect 8435 19329 8447 19363
rect 8389 19323 8447 19329
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9953 19363 10011 19369
rect 9953 19360 9965 19363
rect 9456 19332 9965 19360
rect 9456 19320 9462 19332
rect 9953 19329 9965 19332
rect 9999 19360 10011 19363
rect 10962 19360 10968 19372
rect 9999 19332 10968 19360
rect 9999 19329 10011 19332
rect 9953 19323 10011 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 13078 19360 13084 19372
rect 13039 19332 13084 19360
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 14274 19360 14280 19372
rect 13740 19332 14280 19360
rect 6687 19264 6960 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7558 19292 7564 19304
rect 7340 19264 7564 19292
rect 7340 19252 7346 19264
rect 7558 19252 7564 19264
rect 7616 19292 7622 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7616 19264 7665 19292
rect 7616 19252 7622 19264
rect 7653 19261 7665 19264
rect 7699 19292 7711 19295
rect 8297 19295 8355 19301
rect 8297 19292 8309 19295
rect 7699 19264 8309 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 8297 19261 8309 19264
rect 8343 19261 8355 19295
rect 8297 19255 8355 19261
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 9674 19292 9680 19304
rect 8987 19264 9680 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 10376 19264 10425 19292
rect 10376 19252 10382 19264
rect 10413 19261 10425 19264
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 11057 19295 11115 19301
rect 11057 19261 11069 19295
rect 11103 19292 11115 19295
rect 11146 19292 11152 19304
rect 11103 19264 11152 19292
rect 11103 19261 11115 19264
rect 11057 19255 11115 19261
rect 11146 19252 11152 19264
rect 11204 19292 11210 19304
rect 11204 19264 11560 19292
rect 11204 19252 11210 19264
rect 1670 19224 1676 19236
rect 1631 19196 1676 19224
rect 1670 19184 1676 19196
rect 1728 19184 1734 19236
rect 2501 19227 2559 19233
rect 2501 19193 2513 19227
rect 2547 19224 2559 19227
rect 2700 19224 2728 19252
rect 2547 19196 2728 19224
rect 4516 19227 4574 19233
rect 2547 19193 2559 19196
rect 2501 19187 2559 19193
rect 4516 19193 4528 19227
rect 4562 19224 4574 19227
rect 5166 19224 5172 19236
rect 4562 19196 5172 19224
rect 4562 19193 4574 19196
rect 4516 19187 4574 19193
rect 5166 19184 5172 19196
rect 5224 19184 5230 19236
rect 9861 19227 9919 19233
rect 9861 19224 9873 19227
rect 9232 19196 9873 19224
rect 9232 19168 9260 19196
rect 9861 19193 9873 19196
rect 9907 19193 9919 19227
rect 11330 19224 11336 19236
rect 11291 19196 11336 19224
rect 9861 19187 9919 19193
rect 11330 19184 11336 19196
rect 11388 19184 11394 19236
rect 11532 19224 11560 19264
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12216 19264 12909 19292
rect 12216 19252 12222 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13740 19292 13768 19332
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 14642 19360 14648 19372
rect 14603 19332 14648 19360
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 15838 19360 15844 19372
rect 15799 19332 15844 19360
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 15562 19292 15568 19304
rect 13587 19264 13768 19292
rect 15523 19264 15568 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 15562 19252 15568 19264
rect 15620 19292 15626 19304
rect 16301 19295 16359 19301
rect 16301 19292 16313 19295
rect 15620 19264 16313 19292
rect 15620 19252 15626 19264
rect 16301 19261 16313 19264
rect 16347 19261 16359 19295
rect 16301 19255 16359 19261
rect 13630 19224 13636 19236
rect 11532 19196 13636 19224
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 14369 19227 14427 19233
rect 14369 19224 14381 19227
rect 14240 19196 14381 19224
rect 14240 19184 14246 19196
rect 14369 19193 14381 19196
rect 14415 19224 14427 19227
rect 15013 19227 15071 19233
rect 15013 19224 15025 19227
rect 14415 19196 15025 19224
rect 14415 19193 14427 19196
rect 14369 19187 14427 19193
rect 15013 19193 15025 19196
rect 15059 19193 15071 19227
rect 15013 19187 15071 19193
rect 2682 19156 2688 19168
rect 2643 19128 2688 19156
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3510 19156 3516 19168
rect 3191 19128 3516 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 3602 19116 3608 19168
rect 3660 19156 3666 19168
rect 3970 19156 3976 19168
rect 3660 19128 3976 19156
rect 3660 19116 3666 19128
rect 3970 19116 3976 19128
rect 4028 19156 4034 19168
rect 4065 19159 4123 19165
rect 4065 19156 4077 19159
rect 4028 19128 4077 19156
rect 4028 19116 4034 19128
rect 4065 19125 4077 19128
rect 4111 19125 4123 19159
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 4065 19119 4123 19125
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7800 19128 7849 19156
rect 7800 19116 7806 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 8202 19156 8208 19168
rect 8163 19128 8208 19156
rect 7837 19119 7895 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 9364 19128 9413 19156
rect 9364 19116 9370 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 9490 19116 9496 19168
rect 9548 19156 9554 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9548 19128 9781 19156
rect 9548 19116 9554 19128
rect 9769 19125 9781 19128
rect 9815 19125 9827 19159
rect 11882 19156 11888 19168
rect 11843 19128 11888 19156
rect 9769 19119 9827 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12158 19156 12164 19168
rect 12119 19128 12164 19156
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 12802 19156 12808 19168
rect 12763 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13998 19156 14004 19168
rect 13959 19128 14004 19156
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 15378 19156 15384 19168
rect 15339 19128 15384 19156
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 3142 18952 3148 18964
rect 2832 18924 3148 18952
rect 2832 18912 2838 18924
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 3878 18952 3884 18964
rect 3839 18924 3884 18952
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 4246 18952 4252 18964
rect 4207 18924 4252 18952
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 4706 18952 4712 18964
rect 4667 18924 4712 18952
rect 4706 18912 4712 18924
rect 4764 18952 4770 18964
rect 5629 18955 5687 18961
rect 5629 18952 5641 18955
rect 4764 18924 5641 18952
rect 4764 18912 4770 18924
rect 5629 18921 5641 18924
rect 5675 18921 5687 18955
rect 5629 18915 5687 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7837 18955 7895 18961
rect 7837 18952 7849 18955
rect 7064 18924 7849 18952
rect 7064 18912 7070 18924
rect 7837 18921 7849 18924
rect 7883 18952 7895 18955
rect 8202 18952 8208 18964
rect 7883 18924 8208 18952
rect 7883 18921 7895 18924
rect 7837 18915 7895 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 8352 18924 8493 18952
rect 8352 18912 8358 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 9674 18952 9680 18964
rect 9635 18924 9680 18952
rect 8481 18915 8539 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 10134 18952 10140 18964
rect 10095 18924 10140 18952
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 12897 18955 12955 18961
rect 12897 18921 12909 18955
rect 12943 18952 12955 18955
rect 13078 18952 13084 18964
rect 12943 18924 13084 18952
rect 12943 18921 12955 18924
rect 12897 18915 12955 18921
rect 13078 18912 13084 18924
rect 13136 18952 13142 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 13136 18924 13461 18952
rect 13136 18912 13142 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 13630 18952 13636 18964
rect 13591 18924 13636 18952
rect 13449 18915 13507 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 14093 18955 14151 18961
rect 14093 18952 14105 18955
rect 13780 18924 14105 18952
rect 13780 18912 13786 18924
rect 14093 18921 14105 18924
rect 14139 18952 14151 18955
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 14139 18924 15301 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 15289 18921 15301 18924
rect 15335 18921 15347 18955
rect 15289 18915 15347 18921
rect 2317 18887 2375 18893
rect 2317 18853 2329 18887
rect 2363 18884 2375 18887
rect 2363 18856 3096 18884
rect 2363 18853 2375 18856
rect 2317 18847 2375 18853
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 3068 18757 3096 18856
rect 4522 18776 4528 18828
rect 4580 18816 4586 18828
rect 4617 18819 4675 18825
rect 4617 18816 4629 18819
rect 4580 18788 4629 18816
rect 4580 18776 4586 18788
rect 4617 18785 4629 18788
rect 4663 18785 4675 18819
rect 5626 18816 5632 18828
rect 4617 18779 4675 18785
rect 4816 18788 5632 18816
rect 4816 18760 4844 18788
rect 5626 18776 5632 18788
rect 5684 18816 5690 18828
rect 6069 18819 6127 18825
rect 6069 18816 6081 18819
rect 5684 18788 6081 18816
rect 5684 18776 5690 18788
rect 6069 18785 6081 18788
rect 6115 18785 6127 18819
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 6069 18779 6127 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10962 18825 10968 18828
rect 10945 18819 10968 18825
rect 10945 18816 10957 18819
rect 10376 18788 10957 18816
rect 10376 18776 10382 18788
rect 10945 18785 10957 18788
rect 11020 18816 11026 18828
rect 13998 18816 14004 18828
rect 11020 18788 11093 18816
rect 13959 18788 14004 18816
rect 10945 18779 10968 18785
rect 10962 18776 10968 18779
rect 11020 18776 11026 18788
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3878 18748 3884 18760
rect 3099 18720 3884 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18717 5871 18751
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 5813 18711 5871 18717
rect 7208 18720 8585 18748
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 3510 18680 3516 18692
rect 2455 18652 3516 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 3510 18640 3516 18652
rect 3568 18640 3574 18692
rect 1673 18615 1731 18621
rect 1673 18581 1685 18615
rect 1719 18612 1731 18615
rect 1946 18612 1952 18624
rect 1719 18584 1952 18612
rect 1719 18581 1731 18584
rect 1673 18575 1731 18581
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3384 18584 3433 18612
rect 3384 18572 3390 18584
rect 3421 18581 3433 18584
rect 3467 18612 3479 18615
rect 5166 18612 5172 18624
rect 3467 18584 5172 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 5166 18572 5172 18584
rect 5224 18612 5230 18624
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 5224 18584 5273 18612
rect 5224 18572 5230 18584
rect 5261 18581 5273 18584
rect 5307 18581 5319 18615
rect 5828 18612 5856 18711
rect 7208 18624 7236 18720
rect 8573 18717 8585 18720
rect 8619 18748 8631 18751
rect 9398 18748 9404 18760
rect 8619 18720 9404 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 12529 18751 12587 18757
rect 12529 18717 12541 18751
rect 12575 18748 12587 18751
rect 12802 18748 12808 18760
rect 12575 18720 12808 18748
rect 12575 18717 12587 18720
rect 12529 18711 12587 18717
rect 6546 18612 6552 18624
rect 5828 18584 6552 18612
rect 5261 18575 5319 18581
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 7190 18612 7196 18624
rect 7151 18584 7196 18612
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 7561 18615 7619 18621
rect 7561 18581 7573 18615
rect 7607 18612 7619 18615
rect 7834 18612 7840 18624
rect 7607 18584 7840 18612
rect 7607 18581 7619 18584
rect 7561 18575 7619 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 8294 18612 8300 18624
rect 8067 18584 8300 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 9030 18612 9036 18624
rect 8991 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9398 18612 9404 18624
rect 9359 18584 9404 18612
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 10704 18612 10732 18711
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 14090 18708 14096 18760
rect 14148 18748 14154 18760
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 14148 18720 14197 18748
rect 14148 18708 14154 18720
rect 14185 18717 14197 18720
rect 14231 18717 14243 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 14185 18711 14243 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16482 18748 16488 18760
rect 15979 18720 16488 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 14642 18640 14648 18692
rect 14700 18680 14706 18692
rect 14737 18683 14795 18689
rect 14737 18680 14749 18683
rect 14700 18652 14749 18680
rect 14700 18640 14706 18652
rect 14737 18649 14749 18652
rect 14783 18680 14795 18683
rect 15948 18680 15976 18711
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 14783 18652 15976 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 10870 18612 10876 18624
rect 10643 18584 10876 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 12066 18612 12072 18624
rect 12027 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1394 18408 1400 18420
rect 1355 18380 1400 18408
rect 1394 18368 1400 18380
rect 1452 18368 1458 18420
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4246 18408 4252 18420
rect 4028 18380 4252 18408
rect 4028 18368 4034 18380
rect 4246 18368 4252 18380
rect 4304 18408 4310 18420
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 4304 18380 4445 18408
rect 4304 18368 4310 18380
rect 4433 18377 4445 18380
rect 4479 18377 4491 18411
rect 4798 18408 4804 18420
rect 4759 18380 4804 18408
rect 4433 18371 4491 18377
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 5074 18408 5080 18420
rect 5035 18380 5080 18408
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5442 18408 5448 18420
rect 5403 18380 5448 18408
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 7285 18411 7343 18417
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 9030 18408 9036 18420
rect 7331 18380 9036 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10778 18408 10784 18420
rect 10739 18380 10784 18408
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11112 18380 11376 18408
rect 11112 18368 11118 18380
rect 4816 18340 4844 18368
rect 5813 18343 5871 18349
rect 5813 18340 5825 18343
rect 4816 18312 5825 18340
rect 5813 18309 5825 18312
rect 5859 18309 5871 18343
rect 5813 18303 5871 18309
rect 8202 18300 8208 18352
rect 8260 18340 8266 18352
rect 8297 18343 8355 18349
rect 8297 18340 8309 18343
rect 8260 18312 8309 18340
rect 8260 18300 8266 18312
rect 8297 18309 8309 18312
rect 8343 18309 8355 18343
rect 8297 18303 8355 18309
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 8665 18343 8723 18349
rect 8665 18340 8677 18343
rect 8444 18312 8677 18340
rect 8444 18300 8450 18312
rect 8665 18309 8677 18312
rect 8711 18309 8723 18343
rect 8665 18303 8723 18309
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9861 18343 9919 18349
rect 9861 18340 9873 18343
rect 8895 18312 9873 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 9861 18309 9873 18312
rect 9907 18340 9919 18343
rect 11348 18340 11376 18380
rect 11422 18368 11428 18420
rect 11480 18408 11486 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 11480 18380 12173 18408
rect 11480 18368 11486 18380
rect 12161 18377 12173 18380
rect 12207 18408 12219 18411
rect 12526 18408 12532 18420
rect 12207 18380 12532 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12526 18368 12532 18380
rect 12584 18408 12590 18420
rect 13725 18411 13783 18417
rect 12584 18380 12940 18408
rect 12584 18368 12590 18380
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 9907 18312 11284 18340
rect 11348 18312 11805 18340
rect 9907 18309 9919 18312
rect 9861 18303 9919 18309
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 3050 18272 3056 18284
rect 2832 18244 3056 18272
rect 2832 18232 2838 18244
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7742 18272 7748 18284
rect 6687 18244 7748 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 7834 18232 7840 18284
rect 7892 18272 7898 18284
rect 7892 18244 7937 18272
rect 7892 18232 7898 18244
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9309 18275 9367 18281
rect 9309 18272 9321 18275
rect 9088 18244 9321 18272
rect 9088 18232 9094 18244
rect 9309 18241 9321 18244
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 10318 18272 10324 18284
rect 9539 18244 10324 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 11256 18281 11284 18312
rect 11793 18309 11805 18312
rect 11839 18340 11851 18343
rect 11839 18312 12204 18340
rect 11839 18309 11851 18312
rect 11793 18303 11851 18309
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 12066 18272 12072 18284
rect 11471 18244 12072 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 1394 18164 1400 18216
rect 1452 18204 1458 18216
rect 1854 18204 1860 18216
rect 1452 18176 1860 18204
rect 1452 18164 1458 18176
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 5261 18207 5319 18213
rect 5261 18204 5273 18207
rect 5132 18176 5273 18204
rect 5132 18164 5138 18176
rect 5261 18173 5273 18176
rect 5307 18173 5319 18207
rect 7190 18204 7196 18216
rect 7103 18176 7196 18204
rect 5261 18167 5319 18173
rect 7190 18164 7196 18176
rect 7248 18204 7254 18216
rect 7650 18204 7656 18216
rect 7248 18176 7656 18204
rect 7248 18164 7254 18176
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18204 10747 18207
rect 11440 18204 11468 18235
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 10735 18176 11468 18204
rect 12176 18204 12204 18312
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 12492 18312 12537 18340
rect 12492 18300 12498 18312
rect 12912 18281 12940 18380
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 14090 18408 14096 18420
rect 13771 18380 14096 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 14090 18368 14096 18380
rect 14148 18408 14154 18420
rect 15378 18408 15384 18420
rect 14148 18380 15384 18408
rect 14148 18368 14154 18380
rect 15378 18368 15384 18380
rect 15436 18408 15442 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 15436 18380 15761 18408
rect 15436 18368 15442 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 15749 18371 15807 18377
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14323 18244 14504 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 12986 18204 12992 18216
rect 12176 18176 12992 18204
rect 10735 18173 10747 18176
rect 10689 18167 10747 18173
rect 12986 18164 12992 18176
rect 13044 18204 13050 18216
rect 13096 18204 13124 18235
rect 13044 18176 13124 18204
rect 14369 18207 14427 18213
rect 13044 18164 13050 18176
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 14476 18204 14504 18244
rect 14642 18213 14648 18216
rect 14636 18204 14648 18213
rect 14476 18176 14648 18204
rect 14369 18167 14427 18173
rect 14636 18167 14648 18176
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 1946 18136 1952 18148
rect 1811 18108 1952 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 1946 18096 1952 18108
rect 2004 18096 2010 18148
rect 2958 18136 2964 18148
rect 2871 18108 2964 18136
rect 2958 18096 2964 18108
rect 3016 18136 3022 18148
rect 3298 18139 3356 18145
rect 3298 18136 3310 18139
rect 3016 18108 3310 18136
rect 3016 18096 3022 18108
rect 3298 18105 3310 18108
rect 3344 18105 3356 18139
rect 3298 18099 3356 18105
rect 4522 18096 4528 18148
rect 4580 18136 4586 18148
rect 6181 18139 6239 18145
rect 6181 18136 6193 18139
rect 4580 18108 6193 18136
rect 4580 18096 4586 18108
rect 6181 18105 6193 18108
rect 6227 18105 6239 18139
rect 14384 18136 14412 18167
rect 14642 18164 14648 18167
rect 14700 18164 14706 18216
rect 15746 18164 15752 18216
rect 15804 18204 15810 18216
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 15804 18176 16773 18204
rect 15804 18164 15810 18176
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 14550 18136 14556 18148
rect 14384 18108 14556 18136
rect 6181 18099 6239 18105
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 15654 18096 15660 18148
rect 15712 18136 15718 18148
rect 16025 18139 16083 18145
rect 16025 18136 16037 18139
rect 15712 18108 16037 18136
rect 15712 18096 15718 18108
rect 16025 18105 16037 18108
rect 16071 18105 16083 18139
rect 16025 18099 16083 18105
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2498 18068 2504 18080
rect 2280 18040 2504 18068
rect 2280 18028 2286 18040
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7248 18040 7665 18068
rect 7248 18028 7254 18040
rect 7653 18037 7665 18040
rect 7699 18037 7711 18071
rect 7653 18031 7711 18037
rect 9217 18071 9275 18077
rect 9217 18037 9229 18071
rect 9263 18068 9275 18071
rect 9398 18068 9404 18080
rect 9263 18040 9404 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11330 18068 11336 18080
rect 11195 18040 11336 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 14826 18068 14832 18080
rect 14700 18040 14832 18068
rect 14700 18028 14706 18040
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 16482 18068 16488 18080
rect 16443 18040 16488 18068
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 2866 17864 2872 17876
rect 2455 17836 2872 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 2866 17824 2872 17836
rect 2924 17864 2930 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 2924 17836 3433 17864
rect 2924 17824 2930 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3568 17836 3801 17864
rect 3568 17824 3574 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 3789 17827 3847 17833
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4249 17867 4307 17873
rect 4249 17864 4261 17867
rect 4212 17836 4261 17864
rect 4212 17824 4218 17836
rect 4249 17833 4261 17836
rect 4295 17833 4307 17867
rect 4249 17827 4307 17833
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 4522 17864 4528 17876
rect 4479 17836 4528 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 5905 17867 5963 17873
rect 5905 17833 5917 17867
rect 5951 17864 5963 17867
rect 6546 17864 6552 17876
rect 5951 17836 6552 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6546 17824 6552 17836
rect 6604 17824 6610 17876
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 8757 17867 8815 17873
rect 8757 17864 8769 17867
rect 7892 17836 8769 17864
rect 7892 17824 7898 17836
rect 8757 17833 8769 17836
rect 8803 17833 8815 17867
rect 8757 17827 8815 17833
rect 1394 17756 1400 17808
rect 1452 17796 1458 17808
rect 2777 17799 2835 17805
rect 2777 17796 2789 17799
rect 1452 17768 2789 17796
rect 1452 17756 1458 17768
rect 2777 17765 2789 17768
rect 2823 17796 2835 17799
rect 4062 17796 4068 17808
rect 2823 17768 4068 17796
rect 2823 17765 2835 17768
rect 2777 17759 2835 17765
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 8772 17796 8800 17827
rect 10962 17824 10968 17876
rect 11020 17864 11026 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 11020 17836 11069 17864
rect 11020 17824 11026 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 13722 17864 13728 17876
rect 13683 17836 13728 17864
rect 11057 17827 11115 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 13998 17864 14004 17876
rect 13959 17836 14004 17864
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14182 17864 14188 17876
rect 14143 17836 14188 17864
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 9922 17799 9980 17805
rect 9922 17796 9934 17799
rect 8772 17768 9934 17796
rect 9922 17765 9934 17768
rect 9968 17765 9980 17799
rect 9922 17759 9980 17765
rect 2866 17728 2872 17740
rect 2779 17700 2872 17728
rect 2866 17688 2872 17700
rect 2924 17728 2930 17740
rect 2924 17700 4476 17728
rect 2924 17688 2930 17700
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 1673 17595 1731 17601
rect 1673 17561 1685 17595
rect 1719 17592 1731 17595
rect 1854 17592 1860 17604
rect 1719 17564 1860 17592
rect 1719 17561 1731 17564
rect 1673 17555 1731 17561
rect 1854 17552 1860 17564
rect 1912 17592 1918 17604
rect 2498 17592 2504 17604
rect 1912 17564 2504 17592
rect 1912 17552 1918 17564
rect 2498 17552 2504 17564
rect 2556 17552 2562 17604
rect 4448 17592 4476 17700
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4764 17700 4813 17728
rect 4764 17688 4770 17700
rect 4801 17697 4813 17700
rect 4847 17728 4859 17731
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 4847 17700 5457 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17728 6055 17731
rect 6086 17728 6092 17740
rect 6043 17700 6092 17728
rect 6043 17697 6055 17700
rect 5997 17691 6055 17697
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 7650 17737 7656 17740
rect 7644 17728 7656 17737
rect 7611 17700 7656 17728
rect 7644 17691 7656 17700
rect 7650 17688 7656 17691
rect 7708 17688 7714 17740
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9640 17700 9689 17728
rect 9640 17688 9646 17700
rect 9677 17697 9689 17700
rect 9723 17728 9735 17731
rect 10778 17728 10784 17740
rect 9723 17700 10784 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12233 17731 12291 17737
rect 12233 17728 12245 17731
rect 12124 17700 12245 17728
rect 12124 17688 12130 17700
rect 12233 17697 12245 17700
rect 12279 17697 12291 17731
rect 14660 17728 14688 17827
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 16632 17836 16681 17864
rect 16632 17824 16638 17836
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 14826 17728 14832 17740
rect 14660 17700 14832 17728
rect 12233 17691 12291 17697
rect 14826 17688 14832 17700
rect 14884 17728 14890 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14884 17700 15301 17728
rect 14884 17688 14890 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 15556 17731 15614 17737
rect 15556 17697 15568 17731
rect 15602 17728 15614 17731
rect 15838 17728 15844 17740
rect 15602 17700 15844 17728
rect 15602 17697 15614 17700
rect 15556 17691 15614 17697
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 4890 17660 4896 17672
rect 4851 17632 4896 17660
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 5074 17660 5080 17672
rect 5035 17632 5080 17660
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 6178 17660 6184 17672
rect 6139 17632 6184 17660
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 6604 17632 6929 17660
rect 6604 17620 6610 17632
rect 6917 17629 6929 17632
rect 6963 17660 6975 17663
rect 7374 17660 7380 17672
rect 6963 17632 7380 17660
rect 6963 17629 6975 17632
rect 6917 17623 6975 17629
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 10928 17632 11989 17660
rect 10928 17620 10934 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 6270 17592 6276 17604
rect 4448 17564 6276 17592
rect 6270 17552 6276 17564
rect 6328 17552 6334 17604
rect 2038 17524 2044 17536
rect 1951 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17524 2102 17536
rect 2682 17524 2688 17536
rect 2096 17496 2688 17524
rect 2096 17484 2102 17496
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 7190 17524 7196 17536
rect 7151 17496 7196 17524
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 9122 17524 9128 17536
rect 9083 17496 9128 17524
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 9398 17524 9404 17536
rect 9359 17496 9404 17524
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 11330 17524 11336 17536
rect 11291 17496 11336 17524
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11885 17527 11943 17533
rect 11885 17493 11897 17527
rect 11931 17524 11943 17527
rect 11992 17524 12020 17623
rect 12158 17524 12164 17536
rect 11931 17496 12164 17524
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12894 17484 12900 17536
rect 12952 17524 12958 17536
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 12952 17496 13369 17524
rect 12952 17484 12958 17496
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1452 17292 1593 17320
rect 1452 17280 1458 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2774 17320 2780 17332
rect 1581 17283 1639 17289
rect 2148 17292 2780 17320
rect 2148 17193 2176 17292
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3513 17323 3571 17329
rect 3513 17320 3525 17323
rect 3108 17292 3525 17320
rect 3108 17280 3114 17292
rect 3513 17289 3525 17292
rect 3559 17320 3571 17323
rect 3789 17323 3847 17329
rect 3789 17320 3801 17323
rect 3559 17292 3801 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3789 17289 3801 17292
rect 3835 17289 3847 17323
rect 4246 17320 4252 17332
rect 4207 17292 4252 17320
rect 3789 17283 3847 17289
rect 4246 17280 4252 17292
rect 4304 17280 4310 17332
rect 4706 17320 4712 17332
rect 4667 17292 4712 17320
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5132 17292 5733 17320
rect 5132 17280 5138 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 5721 17283 5779 17289
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7892 17292 7941 17320
rect 7892 17280 7898 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 7929 17283 7987 17289
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 9398 17320 9404 17332
rect 8159 17292 9404 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 4264 17184 4292 17280
rect 5350 17212 5356 17264
rect 5408 17252 5414 17264
rect 7009 17255 7067 17261
rect 7009 17252 7021 17255
rect 5408 17224 7021 17252
rect 5408 17212 5414 17224
rect 7009 17221 7021 17224
rect 7055 17221 7067 17255
rect 7009 17215 7067 17221
rect 5258 17184 5264 17196
rect 4264 17156 5264 17184
rect 2133 17147 2191 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 7944 17184 7972 17283
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 11330 17320 11336 17332
rect 9907 17292 11336 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 9214 17252 9220 17264
rect 8680 17224 9220 17252
rect 8680 17193 8708 17224
rect 9214 17212 9220 17224
rect 9272 17252 9278 17264
rect 9677 17255 9735 17261
rect 9677 17252 9689 17255
rect 9272 17224 9689 17252
rect 9272 17212 9278 17224
rect 9677 17221 9689 17224
rect 9723 17221 9735 17255
rect 9677 17215 9735 17221
rect 9950 17212 9956 17264
rect 10008 17252 10014 17264
rect 11146 17252 11152 17264
rect 10008 17224 11152 17252
rect 10008 17212 10014 17224
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 12894 17212 12900 17264
rect 12952 17252 12958 17264
rect 13909 17255 13967 17261
rect 13909 17252 13921 17255
rect 12952 17224 13921 17252
rect 12952 17212 12958 17224
rect 13909 17221 13921 17224
rect 13955 17221 13967 17255
rect 13909 17215 13967 17221
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 7944 17156 8677 17184
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9180 17156 9413 17184
rect 9180 17144 9186 17156
rect 9401 17153 9413 17156
rect 9447 17184 9459 17187
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 9447 17156 10517 17184
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 10505 17153 10517 17156
rect 10551 17184 10563 17187
rect 10962 17184 10968 17196
rect 10551 17156 10968 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17184 13050 17196
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13044 17156 13461 17184
rect 13044 17144 13050 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13924 17184 13952 17215
rect 16850 17184 16856 17196
rect 13924 17156 14228 17184
rect 16811 17156 16856 17184
rect 13449 17147 13507 17153
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 2389 17119 2447 17125
rect 2389 17116 2401 17119
rect 2280 17088 2401 17116
rect 2280 17076 2286 17088
rect 2389 17085 2401 17088
rect 2435 17085 2447 17119
rect 2389 17079 2447 17085
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 4798 17116 4804 17128
rect 4304 17088 4804 17116
rect 4304 17076 4310 17088
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 842 17008 848 17060
rect 900 17048 906 17060
rect 2041 17051 2099 17057
rect 2041 17048 2053 17051
rect 900 17020 2053 17048
rect 900 17008 906 17020
rect 2041 17017 2053 17020
rect 2087 17048 2099 17051
rect 2866 17048 2872 17060
rect 2087 17020 2872 17048
rect 2087 17017 2099 17020
rect 2041 17011 2099 17017
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 5169 17051 5227 17057
rect 5169 17048 5181 17051
rect 4632 17020 5181 17048
rect 4632 16992 4660 17020
rect 5169 17017 5181 17020
rect 5215 17017 5227 17051
rect 5169 17011 5227 17017
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 6549 17051 6607 17057
rect 6549 17048 6561 17051
rect 5592 17020 6561 17048
rect 5592 17008 5598 17020
rect 6549 17017 6561 17020
rect 6595 17048 6607 17051
rect 6840 17048 6868 17079
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8352 17088 8493 17116
rect 8352 17076 8358 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8846 17116 8852 17128
rect 8619 17088 8852 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8846 17076 8852 17088
rect 8904 17116 8910 17128
rect 9306 17116 9312 17128
rect 8904 17088 9312 17116
rect 8904 17076 8910 17088
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9858 17116 9864 17128
rect 9416 17088 9864 17116
rect 9416 17060 9444 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17116 12311 17119
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12299 17088 12817 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12805 17085 12817 17088
rect 12851 17116 12863 17119
rect 13170 17116 13176 17128
rect 12851 17088 13176 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 13630 17116 13636 17128
rect 13228 17088 13636 17116
rect 13228 17076 13234 17088
rect 13630 17076 13636 17088
rect 13688 17076 13694 17128
rect 14090 17116 14096 17128
rect 14051 17088 14096 17116
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14200 17116 14228 17156
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 14349 17119 14407 17125
rect 14349 17116 14361 17119
rect 14200 17088 14361 17116
rect 14349 17085 14361 17088
rect 14395 17085 14407 17119
rect 14349 17079 14407 17085
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 16761 17119 16819 17125
rect 16761 17116 16773 17119
rect 16724 17088 16773 17116
rect 16724 17076 16730 17088
rect 16761 17085 16773 17088
rect 16807 17085 16819 17119
rect 16761 17079 16819 17085
rect 6595 17020 6868 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 9398 17008 9404 17060
rect 9456 17008 9462 17060
rect 9950 17008 9956 17060
rect 10008 17048 10014 17060
rect 10229 17051 10287 17057
rect 10229 17048 10241 17051
rect 10008 17020 10241 17048
rect 10008 17008 10014 17020
rect 10229 17017 10241 17020
rect 10275 17048 10287 17051
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 10275 17020 10885 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 10873 17017 10885 17020
rect 10919 17017 10931 17051
rect 11790 17048 11796 17060
rect 11751 17020 11796 17048
rect 10873 17011 10931 17017
rect 11790 17008 11796 17020
rect 11848 17048 11854 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 11848 17020 12909 17048
rect 11848 17008 11854 17020
rect 12897 17017 12909 17020
rect 12943 17048 12955 17051
rect 16209 17051 16267 17057
rect 16209 17048 16221 17051
rect 12943 17020 16221 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 16209 17017 16221 17020
rect 16255 17048 16267 17051
rect 16255 17020 16712 17048
rect 16255 17017 16267 17020
rect 16209 17011 16267 17017
rect 4614 16980 4620 16992
rect 4575 16952 4620 16980
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 5077 16983 5135 16989
rect 5077 16980 5089 16983
rect 4856 16952 5089 16980
rect 4856 16940 4862 16952
rect 5077 16949 5089 16952
rect 5123 16949 5135 16983
rect 6086 16980 6092 16992
rect 6047 16952 6092 16980
rect 5077 16943 5135 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7377 16983 7435 16989
rect 7377 16980 7389 16983
rect 6972 16952 7389 16980
rect 6972 16940 6978 16952
rect 7377 16949 7389 16952
rect 7423 16980 7435 16983
rect 7650 16980 7656 16992
rect 7423 16952 7656 16980
rect 7423 16949 7435 16952
rect 7377 16943 7435 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 9916 16952 10333 16980
rect 9916 16940 9922 16952
rect 10321 16949 10333 16952
rect 10367 16980 10379 16983
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10367 16952 11253 16980
rect 10367 16949 10379 16952
rect 10321 16943 10379 16949
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 15470 16980 15476 16992
rect 12492 16952 12537 16980
rect 15431 16952 15476 16980
rect 12492 16940 12498 16952
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 15838 16980 15844 16992
rect 15799 16952 15844 16980
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 16574 16980 16580 16992
rect 16347 16952 16580 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16684 16989 16712 17020
rect 16669 16983 16727 16989
rect 16669 16949 16681 16983
rect 16715 16980 16727 16983
rect 16758 16980 16764 16992
rect 16715 16952 16764 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 2222 16776 2228 16788
rect 2183 16748 2228 16776
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 3050 16776 3056 16788
rect 2455 16748 3056 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 3050 16736 3056 16748
rect 3108 16776 3114 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 3108 16748 3433 16776
rect 3108 16736 3114 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 3421 16739 3479 16745
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16776 4123 16779
rect 4798 16776 4804 16788
rect 4111 16748 4804 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 4948 16748 5089 16776
rect 4948 16736 4954 16748
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 6181 16779 6239 16785
rect 6181 16745 6193 16779
rect 6227 16776 6239 16779
rect 6546 16776 6552 16788
rect 6227 16748 6552 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 6917 16779 6975 16785
rect 6917 16745 6929 16779
rect 6963 16776 6975 16779
rect 7006 16776 7012 16788
rect 6963 16748 7012 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 7742 16776 7748 16788
rect 7703 16748 7748 16776
rect 7742 16736 7748 16748
rect 7800 16776 7806 16788
rect 8202 16776 8208 16788
rect 7800 16748 8208 16776
rect 7800 16736 7806 16748
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8352 16748 9137 16776
rect 8352 16736 8358 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9861 16779 9919 16785
rect 9861 16745 9873 16779
rect 9907 16776 9919 16779
rect 9950 16776 9956 16788
rect 9907 16748 9956 16776
rect 9907 16745 9919 16748
rect 9861 16739 9919 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10836 16748 10885 16776
rect 10836 16736 10842 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 11238 16776 11244 16788
rect 11199 16748 11244 16776
rect 10873 16739 10931 16745
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 12066 16776 12072 16788
rect 12027 16748 12072 16776
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12250 16776 12256 16788
rect 12211 16748 12256 16776
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 12526 16776 12532 16788
rect 12400 16748 12532 16776
rect 12400 16736 12406 16748
rect 12526 16736 12532 16748
rect 12584 16776 12590 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 12584 16748 12725 16776
rect 12584 16736 12590 16748
rect 12713 16745 12725 16748
rect 12759 16745 12771 16779
rect 12713 16739 12771 16745
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14884 16748 15025 16776
rect 14884 16736 14890 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 15746 16776 15752 16788
rect 15335 16748 15752 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 2240 16708 2268 16736
rect 2682 16708 2688 16720
rect 2240 16680 2688 16708
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 2777 16711 2835 16717
rect 2777 16677 2789 16711
rect 2823 16708 2835 16711
rect 3326 16708 3332 16720
rect 2823 16680 3332 16708
rect 2823 16677 2835 16680
rect 2777 16671 2835 16677
rect 3326 16668 3332 16680
rect 3384 16668 3390 16720
rect 3881 16711 3939 16717
rect 3881 16677 3893 16711
rect 3927 16708 3939 16711
rect 4908 16708 4936 16736
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 3927 16680 4936 16708
rect 5000 16680 5549 16708
rect 3927 16677 3939 16680
rect 3881 16671 3939 16677
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 2280 16612 2881 16640
rect 2280 16600 2286 16612
rect 2869 16609 2881 16612
rect 2915 16609 2927 16643
rect 2869 16603 2927 16609
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 5000 16640 5028 16680
rect 5537 16677 5549 16680
rect 5583 16708 5595 16711
rect 5626 16708 5632 16720
rect 5583 16680 5632 16708
rect 5583 16677 5595 16680
rect 5537 16671 5595 16677
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 8846 16708 8852 16720
rect 8807 16680 8852 16708
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 10042 16708 10048 16720
rect 9732 16680 10048 16708
rect 9732 16668 9738 16680
rect 10042 16668 10048 16680
rect 10100 16668 10106 16720
rect 12621 16711 12679 16717
rect 12621 16708 12633 16711
rect 12544 16680 12633 16708
rect 12544 16652 12572 16680
rect 12621 16677 12633 16680
rect 12667 16677 12679 16711
rect 12621 16671 12679 16677
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16708 15715 16711
rect 15930 16708 15936 16720
rect 15703 16680 15936 16708
rect 15703 16677 15715 16680
rect 15657 16671 15715 16677
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 16390 16668 16396 16720
rect 16448 16708 16454 16720
rect 17037 16711 17095 16717
rect 17037 16708 17049 16711
rect 16448 16680 17049 16708
rect 16448 16668 16454 16680
rect 17037 16677 17049 16680
rect 17083 16677 17095 16711
rect 17037 16671 17095 16677
rect 4856 16612 5028 16640
rect 4856 16600 4862 16612
rect 5166 16600 5172 16652
rect 5224 16640 5230 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 5224 16612 5457 16640
rect 5224 16600 5230 16612
rect 5445 16609 5457 16612
rect 5491 16609 5503 16643
rect 10226 16640 10232 16652
rect 10139 16612 10232 16640
rect 5445 16603 5503 16609
rect 10226 16600 10232 16612
rect 10284 16640 10290 16652
rect 11330 16640 11336 16652
rect 10284 16612 11336 16640
rect 10284 16600 10290 16612
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15528 16612 16313 16640
rect 15528 16600 15534 16612
rect 16301 16609 16313 16612
rect 16347 16640 16359 16643
rect 16850 16640 16856 16652
rect 16347 16612 16856 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3053 16575 3111 16581
rect 3053 16572 3065 16575
rect 3016 16544 3065 16572
rect 3016 16532 3022 16544
rect 3053 16541 3065 16544
rect 3099 16572 3111 16575
rect 3694 16572 3700 16584
rect 3099 16544 3700 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 7834 16572 7840 16584
rect 7795 16544 7840 16572
rect 5629 16535 5687 16541
rect 5258 16464 5264 16516
rect 5316 16504 5322 16516
rect 5644 16504 5672 16535
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 8018 16572 8024 16584
rect 7979 16544 8024 16572
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 10100 16544 10333 16572
rect 10100 16532 10106 16544
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16541 10563 16575
rect 12802 16572 12808 16584
rect 12763 16544 12808 16572
rect 10505 16535 10563 16541
rect 7374 16504 7380 16516
rect 5316 16476 5672 16504
rect 7335 16476 7380 16504
rect 5316 16464 5322 16476
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 9950 16504 9956 16516
rect 9272 16476 9956 16504
rect 9272 16464 9278 16476
rect 9950 16464 9956 16476
rect 10008 16504 10014 16516
rect 10520 16504 10548 16535
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 15933 16575 15991 16581
rect 15933 16572 15945 16575
rect 15896 16544 15945 16572
rect 15896 16532 15902 16544
rect 15933 16541 15945 16544
rect 15979 16572 15991 16575
rect 17034 16572 17040 16584
rect 15979 16544 17040 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 10008 16476 10548 16504
rect 10008 16464 10014 16476
rect 11698 16464 11704 16516
rect 11756 16504 11762 16516
rect 12526 16504 12532 16516
rect 11756 16476 12532 16504
rect 11756 16464 11762 16476
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 15764 16504 15792 16532
rect 12636 16476 15792 16504
rect 7285 16439 7343 16445
rect 7285 16405 7297 16439
rect 7331 16436 7343 16439
rect 7558 16436 7564 16448
rect 7331 16408 7564 16436
rect 7331 16405 7343 16408
rect 7285 16399 7343 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 8386 16436 8392 16448
rect 8347 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12636 16436 12664 16476
rect 12032 16408 12664 16436
rect 12032 16396 12038 16408
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 13817 16439 13875 16445
rect 13817 16436 13829 16439
rect 13780 16408 13829 16436
rect 13780 16396 13786 16408
rect 13817 16405 13829 16408
rect 13863 16436 13875 16439
rect 14090 16436 14096 16448
rect 13863 16408 14096 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 14090 16396 14096 16408
rect 14148 16436 14154 16448
rect 14185 16439 14243 16445
rect 14185 16436 14197 16439
rect 14148 16408 14197 16436
rect 14148 16396 14154 16408
rect 14185 16405 14197 16408
rect 14231 16405 14243 16439
rect 14185 16399 14243 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2682 16192 2688 16244
rect 2740 16232 2746 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2740 16204 2973 16232
rect 2740 16192 2746 16204
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 2961 16195 3019 16201
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 4798 16232 4804 16244
rect 4755 16204 4804 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5442 16232 5448 16244
rect 5215 16204 5448 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 8294 16232 8300 16244
rect 8255 16204 8300 16232
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 8570 16232 8576 16244
rect 8531 16204 8576 16232
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 9858 16232 9864 16244
rect 9815 16204 9864 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10870 16232 10876 16244
rect 10831 16204 10876 16232
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11756 16204 11805 16232
rect 11756 16192 11762 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 12342 16232 12348 16244
rect 12299 16204 12348 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 15197 16235 15255 16241
rect 15197 16201 15209 16235
rect 15243 16232 15255 16235
rect 15838 16232 15844 16244
rect 15243 16204 15844 16232
rect 15243 16201 15255 16204
rect 15197 16195 15255 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16022 16232 16028 16244
rect 15983 16204 16028 16232
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 10226 16164 10232 16176
rect 9723 16136 10232 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 10226 16124 10232 16136
rect 10284 16124 10290 16176
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 15565 16167 15623 16173
rect 12216 16136 13032 16164
rect 12216 16124 12222 16136
rect 13004 16108 13032 16136
rect 15565 16133 15577 16167
rect 15611 16164 15623 16167
rect 15930 16164 15936 16176
rect 15611 16136 15936 16164
rect 15611 16133 15623 16136
rect 15565 16127 15623 16133
rect 15930 16124 15936 16136
rect 15988 16124 15994 16176
rect 3326 16096 3332 16108
rect 3287 16068 3332 16096
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16096 4215 16099
rect 5534 16096 5540 16108
rect 4203 16068 5540 16096
rect 4203 16065 4215 16068
rect 4157 16059 4215 16065
rect 5534 16056 5540 16068
rect 5592 16056 5598 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6086 16096 6092 16108
rect 5859 16068 6092 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 6914 16096 6920 16108
rect 6144 16068 6920 16096
rect 6144 16056 6150 16068
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7558 16096 7564 16108
rect 7515 16068 7564 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 9950 16056 9956 16108
rect 10008 16096 10014 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10008 16068 10333 16096
rect 10008 16056 10014 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 10321 16059 10379 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 12618 16096 12624 16108
rect 12579 16068 12624 16096
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13722 16096 13728 16108
rect 13044 16068 13728 16096
rect 13044 16056 13050 16068
rect 13722 16056 13728 16068
rect 13780 16096 13786 16108
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 13780 16068 13829 16096
rect 13780 16056 13786 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 16574 16096 16580 16108
rect 16535 16068 16580 16096
rect 13817 16059 13875 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 3878 16028 3884 16040
rect 3839 16000 3884 16028
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 5994 16028 6000 16040
rect 5675 16000 6000 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 5994 15988 6000 16000
rect 6052 16028 6058 16040
rect 6181 16031 6239 16037
rect 6181 16028 6193 16031
rect 6052 16000 6193 16028
rect 6052 15988 6058 16000
rect 6181 15997 6193 16000
rect 6227 16028 6239 16031
rect 6549 16031 6607 16037
rect 6549 16028 6561 16031
rect 6227 16000 6561 16028
rect 6227 15997 6239 16000
rect 6181 15991 6239 15997
rect 6549 15997 6561 16000
rect 6595 16028 6607 16031
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6595 16000 7297 16028
rect 6595 15997 6607 16000
rect 6549 15991 6607 15997
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 7285 15991 7343 15997
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 10229 16031 10287 16037
rect 10229 15997 10241 16031
rect 10275 16028 10287 16031
rect 10870 16028 10876 16040
rect 10275 16000 10876 16028
rect 10275 15997 10287 16000
rect 10229 15991 10287 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12492 16000 13185 16028
rect 12492 15988 12498 16000
rect 13173 15997 13185 16000
rect 13219 15997 13231 16031
rect 13173 15991 13231 15997
rect 1848 15963 1906 15969
rect 1848 15929 1860 15963
rect 1894 15960 1906 15963
rect 2038 15960 2044 15972
rect 1894 15932 2044 15960
rect 1894 15929 1906 15932
rect 1848 15923 1906 15929
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 7834 15960 7840 15972
rect 5552 15932 7840 15960
rect 5552 15904 5580 15932
rect 7834 15920 7840 15932
rect 7892 15920 7898 15972
rect 10134 15960 10140 15972
rect 10047 15932 10140 15960
rect 10134 15920 10140 15932
rect 10192 15960 10198 15972
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 10192 15932 11161 15960
rect 10192 15920 10198 15932
rect 11149 15929 11161 15932
rect 11195 15929 11207 15963
rect 14062 15963 14120 15969
rect 14062 15960 14074 15963
rect 11149 15923 11207 15929
rect 13648 15932 14074 15960
rect 3694 15892 3700 15904
rect 3655 15864 3700 15892
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15892 5135 15895
rect 5166 15892 5172 15904
rect 5123 15864 5172 15892
rect 5123 15861 5135 15864
rect 5077 15855 5135 15861
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 7064 15864 7205 15892
rect 7064 15852 7070 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13648 15901 13676 15932
rect 14062 15929 14074 15932
rect 14108 15960 14120 15963
rect 14182 15960 14188 15972
rect 14108 15932 14188 15960
rect 14108 15929 14120 15932
rect 14062 15923 14120 15929
rect 14182 15920 14188 15932
rect 14240 15920 14246 15972
rect 15746 15920 15752 15972
rect 15804 15960 15810 15972
rect 15933 15963 15991 15969
rect 15933 15960 15945 15963
rect 15804 15932 15945 15960
rect 15804 15920 15810 15932
rect 15933 15929 15945 15932
rect 15979 15960 15991 15963
rect 16942 15960 16948 15972
rect 15979 15932 16948 15960
rect 15979 15929 15991 15932
rect 15933 15923 15991 15929
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 13633 15895 13691 15901
rect 13633 15892 13645 15895
rect 13412 15864 13645 15892
rect 13412 15852 13418 15864
rect 13633 15861 13645 15864
rect 13679 15861 13691 15895
rect 16390 15892 16396 15904
rect 16351 15864 16396 15892
rect 13633 15855 13691 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 17494 15892 17500 15904
rect 16540 15864 16585 15892
rect 17455 15864 17500 15892
rect 16540 15852 16546 15864
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 2038 15688 2044 15700
rect 1719 15660 2044 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 2372 15660 2421 15688
rect 2372 15648 2378 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 2409 15651 2467 15657
rect 2777 15691 2835 15697
rect 2777 15657 2789 15691
rect 2823 15688 2835 15691
rect 3050 15688 3056 15700
rect 2823 15660 3056 15688
rect 2823 15657 2835 15660
rect 2777 15651 2835 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4893 15691 4951 15697
rect 4893 15688 4905 15691
rect 4212 15660 4905 15688
rect 4212 15648 4218 15660
rect 4893 15657 4905 15660
rect 4939 15688 4951 15691
rect 5534 15688 5540 15700
rect 4939 15660 5540 15688
rect 4939 15657 4951 15660
rect 4893 15651 4951 15657
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 6086 15688 6092 15700
rect 6047 15660 6092 15688
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 6638 15688 6644 15700
rect 6599 15660 6644 15688
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 10042 15688 10048 15700
rect 9539 15660 10048 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 12345 15691 12403 15697
rect 12345 15657 12357 15691
rect 12391 15688 12403 15691
rect 12802 15688 12808 15700
rect 12391 15660 12808 15688
rect 12391 15657 12403 15660
rect 12345 15651 12403 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15749 15691 15807 15697
rect 15749 15688 15761 15691
rect 15436 15660 15761 15688
rect 15436 15648 15442 15660
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 5258 15620 5264 15632
rect 4663 15592 5264 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 6454 15580 6460 15632
rect 6512 15620 6518 15632
rect 8478 15620 8484 15632
rect 6512 15592 8331 15620
rect 8439 15592 8484 15620
rect 6512 15580 6518 15592
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2740 15524 2881 15552
rect 2740 15512 2746 15524
rect 2869 15521 2881 15524
rect 2915 15552 2927 15555
rect 3421 15555 3479 15561
rect 3421 15552 3433 15555
rect 2915 15524 3433 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 3421 15521 3433 15524
rect 3467 15521 3479 15555
rect 3421 15515 3479 15521
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 5442 15552 5448 15564
rect 4764 15524 5448 15552
rect 4764 15512 4770 15524
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 6270 15552 6276 15564
rect 5583 15524 6276 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6788 15524 7021 15552
rect 6788 15512 6794 15524
rect 7009 15521 7021 15524
rect 7055 15552 7067 15555
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7055 15524 8033 15552
rect 7055 15521 7067 15524
rect 7009 15515 7067 15521
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 8021 15515 8079 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8303 15552 8331 15592
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 9030 15620 9036 15632
rect 8943 15592 9036 15620
rect 9030 15580 9036 15592
rect 9088 15620 9094 15632
rect 9582 15620 9588 15632
rect 9088 15592 9588 15620
rect 9088 15580 9094 15592
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 9950 15620 9956 15632
rect 9911 15592 9956 15620
rect 9950 15580 9956 15592
rect 10008 15580 10014 15632
rect 9490 15552 9496 15564
rect 8303 15524 9496 15552
rect 9490 15512 9496 15524
rect 9548 15552 9554 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 9548 15524 10425 15552
rect 9548 15512 9554 15524
rect 10413 15521 10425 15524
rect 10459 15552 10471 15555
rect 12066 15552 12072 15564
rect 10459 15524 12072 15552
rect 10459 15521 10471 15524
rect 10413 15515 10471 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13061 15555 13119 15561
rect 13061 15552 13073 15555
rect 12952 15524 13073 15552
rect 12952 15512 12958 15524
rect 13061 15521 13073 15524
rect 13107 15552 13119 15555
rect 14461 15555 14519 15561
rect 14461 15552 14473 15555
rect 13107 15524 14473 15552
rect 13107 15521 13119 15524
rect 13061 15515 13119 15521
rect 14461 15521 14473 15524
rect 14507 15552 14519 15555
rect 14550 15552 14556 15564
rect 14507 15524 14556 15552
rect 14507 15521 14519 15524
rect 14461 15515 14519 15521
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 2961 15487 3019 15493
rect 2961 15484 2973 15487
rect 2096 15456 2973 15484
rect 2096 15444 2102 15456
rect 2961 15453 2973 15456
rect 3007 15484 3019 15487
rect 3234 15484 3240 15496
rect 3007 15456 3240 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5258 15484 5264 15496
rect 5132 15456 5264 15484
rect 5132 15444 5138 15456
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5721 15487 5779 15493
rect 5721 15453 5733 15487
rect 5767 15484 5779 15487
rect 6454 15484 6460 15496
rect 5767 15456 6460 15484
rect 5767 15453 5779 15456
rect 5721 15447 5779 15453
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15484 6607 15487
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 6595 15456 7113 15484
rect 6595 15453 6607 15456
rect 6549 15447 6607 15453
rect 7101 15453 7113 15456
rect 7147 15484 7159 15487
rect 7190 15484 7196 15496
rect 7147 15456 7196 15484
rect 7147 15453 7159 15456
rect 7101 15447 7159 15453
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 7285 15487 7343 15493
rect 7285 15453 7297 15487
rect 7331 15484 7343 15487
rect 7650 15484 7656 15496
rect 7331 15456 7656 15484
rect 7331 15453 7343 15456
rect 7285 15447 7343 15453
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 9916 15456 10517 15484
rect 9916 15444 9922 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 11054 15484 11060 15496
rect 10735 15456 11060 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 11054 15444 11060 15456
rect 11112 15444 11118 15496
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15484 11851 15487
rect 12526 15484 12532 15496
rect 11839 15456 12532 15484
rect 11839 15453 11851 15456
rect 11793 15447 11851 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12805 15487 12863 15493
rect 12805 15453 12817 15487
rect 12851 15453 12863 15487
rect 12805 15447 12863 15453
rect 3878 15416 3884 15428
rect 3791 15388 3884 15416
rect 3878 15376 3884 15388
rect 3936 15416 3942 15428
rect 9582 15416 9588 15428
rect 3936 15388 9588 15416
rect 3936 15376 3942 15388
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 5074 15348 5080 15360
rect 5035 15320 5080 15348
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 8018 15348 8024 15360
rect 7791 15320 8024 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 8018 15308 8024 15320
rect 8076 15348 8082 15360
rect 8570 15348 8576 15360
rect 8076 15320 8576 15348
rect 8076 15308 8082 15320
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12713 15351 12771 15357
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 12820 15348 12848 15447
rect 13906 15376 13912 15428
rect 13964 15416 13970 15428
rect 15289 15419 15347 15425
rect 15289 15416 15301 15419
rect 13964 15388 15301 15416
rect 13964 15376 13970 15388
rect 15289 15385 15301 15388
rect 15335 15385 15347 15419
rect 15488 15416 15516 15660
rect 15749 15657 15761 15660
rect 15795 15657 15807 15691
rect 15749 15651 15807 15657
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 16540 15660 16865 15688
rect 16540 15648 16546 15660
rect 16853 15657 16865 15660
rect 16899 15688 16911 15691
rect 17770 15688 17776 15700
rect 16899 15660 17776 15688
rect 16899 15657 16911 15660
rect 16853 15651 16911 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 16666 15620 16672 15632
rect 16627 15592 16672 15620
rect 16666 15580 16672 15592
rect 16724 15620 16730 15632
rect 17313 15623 17371 15629
rect 17313 15620 17325 15623
rect 16724 15592 17325 15620
rect 16724 15580 16730 15592
rect 17313 15589 17325 15592
rect 17359 15589 17371 15623
rect 17313 15583 17371 15589
rect 21082 15580 21088 15632
rect 21140 15620 21146 15632
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 21140 15592 21189 15620
rect 21140 15580 21146 15592
rect 21177 15589 21189 15592
rect 21223 15589 21235 15623
rect 21177 15583 21235 15589
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 15620 15524 15669 15552
rect 15620 15512 15626 15524
rect 15657 15521 15669 15524
rect 15703 15552 15715 15555
rect 15930 15552 15936 15564
rect 15703 15524 15936 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 17494 15552 17500 15564
rect 17267 15524 17500 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 17494 15512 17500 15524
rect 17552 15552 17558 15564
rect 17862 15552 17868 15564
rect 17552 15524 17868 15552
rect 17552 15512 17558 15524
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 20898 15552 20904 15564
rect 20859 15524 20904 15552
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 15838 15484 15844 15496
rect 15799 15456 15844 15484
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 17402 15484 17408 15496
rect 17363 15456 17408 15484
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 15562 15416 15568 15428
rect 15488 15388 15568 15416
rect 15289 15379 15347 15385
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 12986 15348 12992 15360
rect 12759 15320 12992 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 15105 15351 15163 15357
rect 15105 15317 15117 15351
rect 15151 15348 15163 15351
rect 15378 15348 15384 15360
rect 15151 15320 15384 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 16393 15351 16451 15357
rect 16393 15317 16405 15351
rect 16439 15348 16451 15351
rect 16482 15348 16488 15360
rect 16439 15320 16488 15348
rect 16439 15317 16451 15320
rect 16393 15311 16451 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 18138 15348 18144 15360
rect 18051 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15348 18202 15360
rect 18506 15348 18512 15360
rect 18196 15320 18512 15348
rect 18196 15308 18202 15320
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3234 15144 3240 15156
rect 3195 15116 3240 15144
rect 3234 15104 3240 15116
rect 3292 15144 3298 15156
rect 3513 15147 3571 15153
rect 3513 15144 3525 15147
rect 3292 15116 3525 15144
rect 3292 15104 3298 15116
rect 3513 15113 3525 15116
rect 3559 15113 3571 15147
rect 3513 15107 3571 15113
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 5905 15147 5963 15153
rect 5500 15116 5672 15144
rect 5500 15104 5506 15116
rect 5534 15076 5540 15088
rect 5495 15048 5540 15076
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 5644 15076 5672 15116
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 6270 15144 6276 15156
rect 5951 15116 6276 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10045 15147 10103 15153
rect 10045 15113 10057 15147
rect 10091 15144 10103 15147
rect 10134 15144 10140 15156
rect 10091 15116 10140 15144
rect 10091 15113 10103 15116
rect 10045 15107 10103 15113
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 11020 15116 11069 15144
rect 11020 15104 11026 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11057 15107 11115 15113
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13814 15144 13820 15156
rect 12492 15116 12537 15144
rect 13775 15116 13820 15144
rect 12492 15104 12498 15116
rect 13814 15104 13820 15116
rect 13872 15144 13878 15156
rect 14458 15144 14464 15156
rect 13872 15116 14464 15144
rect 13872 15104 13878 15116
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 17678 15104 17684 15156
rect 17736 15144 17742 15156
rect 17773 15147 17831 15153
rect 17773 15144 17785 15147
rect 17736 15116 17785 15144
rect 17736 15104 17742 15116
rect 17773 15113 17785 15116
rect 17819 15113 17831 15147
rect 17773 15107 17831 15113
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 18012 15116 18061 15144
rect 18012 15104 18018 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 20898 15144 20904 15156
rect 20859 15116 20904 15144
rect 18049 15107 18107 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 6181 15079 6239 15085
rect 6181 15076 6193 15079
rect 5644 15048 6193 15076
rect 6181 15045 6193 15048
rect 6227 15045 6239 15079
rect 6181 15039 6239 15045
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1857 15011 1915 15017
rect 1857 15008 1869 15011
rect 1636 14980 1869 15008
rect 1636 14968 1642 14980
rect 1857 14977 1869 14980
rect 1903 14977 1915 15011
rect 10686 15008 10692 15020
rect 10599 14980 10692 15008
rect 1857 14971 1915 14977
rect 1872 14940 1900 14971
rect 10686 14968 10692 14980
rect 10744 15008 10750 15020
rect 10980 15008 11008 15104
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 12584 15048 13461 15076
rect 12584 15036 12590 15048
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 13449 15039 13507 15045
rect 10744 14980 11008 15008
rect 12253 15011 12311 15017
rect 10744 14968 10750 14980
rect 12253 14977 12265 15011
rect 12299 15008 12311 15011
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12299 14980 13001 15008
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 12989 14977 13001 14980
rect 13035 15008 13047 15011
rect 13354 15008 13360 15020
rect 13035 14980 13360 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 4154 14940 4160 14952
rect 1872 14912 4160 14940
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 6914 14940 6920 14952
rect 6871 14912 6920 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 13464 14940 13492 15039
rect 14550 15008 14556 15020
rect 14511 14980 14556 15008
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 13464 14912 14381 14940
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 14516 14912 14561 14940
rect 14516 14900 14522 14912
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 15436 14912 15761 14940
rect 15436 14900 15442 14912
rect 15749 14909 15761 14912
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18616 14940 18644 14971
rect 18012 14912 18644 14940
rect 18012 14900 18018 14912
rect 1765 14875 1823 14881
rect 1765 14841 1777 14875
rect 1811 14872 1823 14875
rect 2102 14875 2160 14881
rect 2102 14872 2114 14875
rect 1811 14844 2114 14872
rect 1811 14841 1823 14844
rect 1765 14835 1823 14841
rect 2102 14841 2114 14844
rect 2148 14872 2160 14875
rect 2222 14872 2228 14884
rect 2148 14844 2228 14872
rect 2148 14841 2160 14844
rect 2102 14835 2160 14841
rect 2222 14832 2228 14844
rect 2280 14832 2286 14884
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 4065 14875 4123 14881
rect 4065 14872 4077 14875
rect 3660 14844 4077 14872
rect 3660 14832 3666 14844
rect 4065 14841 4077 14844
rect 4111 14872 4123 14875
rect 4424 14875 4482 14881
rect 4424 14872 4436 14875
rect 4111 14844 4436 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4424 14841 4436 14844
rect 4470 14872 4482 14875
rect 4522 14872 4528 14884
rect 4470 14844 4528 14872
rect 4470 14841 4482 14844
rect 4424 14835 4482 14841
rect 4522 14832 4528 14844
rect 4580 14832 4586 14884
rect 7006 14832 7012 14884
rect 7064 14881 7070 14884
rect 7064 14875 7128 14881
rect 7064 14841 7082 14875
rect 7116 14841 7128 14875
rect 7064 14835 7128 14841
rect 9217 14875 9275 14881
rect 9217 14841 9229 14875
rect 9263 14872 9275 14875
rect 10413 14875 10471 14881
rect 9263 14844 10364 14872
rect 9263 14841 9275 14844
rect 9217 14835 9275 14841
rect 7064 14832 7070 14835
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6512 14776 6561 14804
rect 6512 14764 6518 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7708 14776 8217 14804
rect 7708 14764 7714 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8205 14767 8263 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10336 14804 10364 14844
rect 10413 14841 10425 14875
rect 10459 14872 10471 14875
rect 10962 14872 10968 14884
rect 10459 14844 10968 14872
rect 10459 14841 10471 14844
rect 10413 14835 10471 14841
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14872 11943 14875
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 11931 14844 12817 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12805 14841 12817 14844
rect 12851 14872 12863 14875
rect 16016 14875 16074 14881
rect 12851 14844 14044 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 10336 14776 10517 14804
rect 10505 14773 10517 14776
rect 10551 14804 10563 14807
rect 11146 14804 11152 14816
rect 10551 14776 11152 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11514 14804 11520 14816
rect 11475 14776 11520 14804
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 14016 14813 14044 14844
rect 16016 14841 16028 14875
rect 16062 14872 16074 14875
rect 16298 14872 16304 14884
rect 16062 14844 16304 14872
rect 16062 14841 16074 14844
rect 16016 14835 16074 14841
rect 16298 14832 16304 14844
rect 16356 14872 16362 14884
rect 17402 14872 17408 14884
rect 16356 14844 17408 14872
rect 16356 14832 16362 14844
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 17678 14832 17684 14884
rect 17736 14872 17742 14884
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 17736 14844 18429 14872
rect 17736 14832 17742 14844
rect 18417 14841 18429 14844
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12584 14776 12909 14804
rect 12584 14764 12590 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 14001 14807 14059 14813
rect 14001 14773 14013 14807
rect 14047 14773 14059 14807
rect 14001 14767 14059 14773
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14804 15439 14807
rect 15930 14804 15936 14816
rect 15427 14776 15936 14804
rect 15427 14773 15439 14776
rect 15381 14767 15439 14773
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 17126 14804 17132 14816
rect 17087 14776 17132 14804
rect 17126 14764 17132 14776
rect 17184 14764 17190 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2682 14600 2688 14612
rect 2455 14572 2688 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 2832 14572 4997 14600
rect 2832 14560 2838 14572
rect 4985 14569 4997 14572
rect 5031 14569 5043 14603
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 4985 14563 5043 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10686 14600 10692 14612
rect 10643 14572 10692 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 15562 14600 15568 14612
rect 15523 14572 15568 14600
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 1820 14504 2912 14532
rect 1820 14492 1826 14504
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2774 14464 2780 14476
rect 2188 14436 2780 14464
rect 2188 14424 2194 14436
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 2884 14473 2912 14504
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 7650 14541 7656 14544
rect 6917 14535 6975 14541
rect 4212 14504 5580 14532
rect 4212 14492 4218 14504
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14464 2927 14467
rect 3789 14467 3847 14473
rect 3789 14464 3801 14467
rect 2915 14436 3801 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 3789 14433 3801 14436
rect 3835 14433 3847 14467
rect 4062 14464 4068 14476
rect 4023 14436 4068 14464
rect 3789 14427 3847 14433
rect 4062 14424 4068 14436
rect 4120 14464 4126 14476
rect 5184 14473 5212 14504
rect 5442 14473 5448 14476
rect 4617 14467 4675 14473
rect 4617 14464 4629 14467
rect 4120 14436 4629 14464
rect 4120 14424 4126 14436
rect 4617 14433 4629 14436
rect 4663 14433 4675 14467
rect 4617 14427 4675 14433
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5436 14464 5448 14473
rect 5403 14436 5448 14464
rect 5169 14427 5227 14433
rect 5436 14427 5448 14436
rect 5442 14424 5448 14427
rect 5500 14424 5506 14476
rect 5552 14464 5580 14504
rect 6917 14501 6929 14535
rect 6963 14532 6975 14535
rect 7644 14532 7656 14541
rect 6963 14504 7656 14532
rect 6963 14501 6975 14504
rect 6917 14495 6975 14501
rect 7644 14495 7656 14504
rect 7650 14492 7656 14495
rect 7708 14492 7714 14544
rect 10778 14492 10784 14544
rect 10836 14532 10842 14544
rect 11026 14535 11084 14541
rect 11026 14532 11038 14535
rect 10836 14504 11038 14532
rect 10836 14492 10842 14504
rect 11026 14501 11038 14504
rect 11072 14501 11084 14535
rect 11026 14495 11084 14501
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 12986 14532 12992 14544
rect 11572 14504 12992 14532
rect 11572 14492 11578 14504
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 16574 14492 16580 14544
rect 16632 14532 16638 14544
rect 16752 14535 16810 14541
rect 16752 14532 16764 14535
rect 16632 14504 16764 14532
rect 16632 14492 16638 14504
rect 16752 14501 16764 14504
rect 16798 14532 16810 14535
rect 17126 14532 17132 14544
rect 16798 14504 17132 14532
rect 16798 14501 16810 14504
rect 16752 14495 16810 14501
rect 17126 14492 17132 14504
rect 17184 14492 17190 14544
rect 7377 14467 7435 14473
rect 5552 14436 6960 14464
rect 6932 14408 6960 14436
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 8938 14464 8944 14476
rect 7423 14436 8944 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2280 14368 3065 14396
rect 2280 14356 2286 14368
rect 3053 14365 3065 14368
rect 3099 14396 3111 14399
rect 3694 14396 3700 14408
rect 3099 14368 3700 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7392 14396 7420 14427
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9490 14464 9496 14476
rect 9403 14436 9496 14464
rect 9490 14424 9496 14436
rect 9548 14464 9554 14476
rect 11532 14464 11560 14492
rect 9548 14436 11560 14464
rect 9548 14424 9554 14436
rect 6972 14368 7420 14396
rect 9677 14399 9735 14405
rect 6972 14356 6978 14368
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 10042 14396 10048 14408
rect 9723 14368 10048 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 10796 14405 10824 14436
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 13245 14467 13303 14473
rect 13245 14464 13257 14467
rect 12768 14436 13257 14464
rect 12768 14424 12774 14436
rect 13245 14433 13257 14436
rect 13291 14433 13303 14467
rect 13245 14427 13303 14433
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14365 10839 14399
rect 12986 14396 12992 14408
rect 12947 14368 12992 14396
rect 10781 14359 10839 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 15378 14396 15384 14408
rect 15151 14368 15384 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 15378 14356 15384 14368
rect 15436 14396 15442 14408
rect 16482 14396 16488 14408
rect 15436 14368 16488 14396
rect 15436 14356 15442 14368
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 4028 14300 4261 14328
rect 4028 14288 4034 14300
rect 4249 14297 4261 14300
rect 4295 14297 4307 14331
rect 4249 14291 4307 14297
rect 10229 14331 10287 14337
rect 10229 14297 10241 14331
rect 10275 14328 10287 14331
rect 12161 14331 12219 14337
rect 10275 14300 10640 14328
rect 10275 14297 10287 14300
rect 10229 14291 10287 14297
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1581 14263 1639 14269
rect 1581 14260 1593 14263
rect 1452 14232 1593 14260
rect 1452 14220 1458 14232
rect 1581 14229 1593 14232
rect 1627 14229 1639 14263
rect 3418 14260 3424 14272
rect 3379 14232 3424 14260
rect 1581 14223 1639 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 6420 14232 6561 14260
rect 6420 14220 6426 14232
rect 6549 14229 6561 14232
rect 6595 14260 6607 14263
rect 7006 14260 7012 14272
rect 6595 14232 7012 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 7006 14220 7012 14232
rect 7064 14260 7070 14272
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 7064 14232 7205 14260
rect 7064 14220 7070 14232
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 8757 14263 8815 14269
rect 8757 14260 8769 14263
rect 8628 14232 8769 14260
rect 8628 14220 8634 14232
rect 8757 14229 8769 14232
rect 8803 14229 8815 14263
rect 10612 14260 10640 14300
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12710 14328 12716 14340
rect 12207 14300 12716 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 15838 14328 15844 14340
rect 15799 14300 15844 14328
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 10962 14260 10968 14272
rect 10612 14232 10968 14260
rect 8757 14223 8815 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 12250 14220 12256 14272
rect 12308 14260 12314 14272
rect 12805 14263 12863 14269
rect 12805 14260 12817 14263
rect 12308 14232 12817 14260
rect 12308 14220 12314 14232
rect 12805 14229 12817 14232
rect 12851 14260 12863 14263
rect 12894 14260 12900 14272
rect 12851 14232 12900 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 12894 14220 12900 14232
rect 12952 14260 12958 14272
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 12952 14232 14381 14260
rect 12952 14220 12958 14232
rect 14369 14229 14381 14232
rect 14415 14229 14427 14263
rect 16298 14260 16304 14272
rect 16259 14232 16304 14260
rect 14369 14223 14427 14229
rect 16298 14220 16304 14232
rect 16356 14260 16362 14272
rect 16850 14260 16856 14272
rect 16356 14232 16856 14260
rect 16356 14220 16362 14232
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17862 14260 17868 14272
rect 17823 14232 17868 14260
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18141 14263 18199 14269
rect 18141 14260 18153 14263
rect 18012 14232 18153 14260
rect 18012 14220 18018 14232
rect 18141 14229 18153 14232
rect 18187 14229 18199 14263
rect 18141 14223 18199 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2409 14059 2467 14065
rect 2409 14056 2421 14059
rect 2372 14028 2421 14056
rect 2372 14016 2378 14028
rect 2409 14025 2421 14028
rect 2455 14025 2467 14059
rect 5442 14056 5448 14068
rect 5403 14028 5448 14056
rect 2409 14019 2467 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5592 14028 5733 14056
rect 5592 14016 5598 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 5721 14019 5779 14025
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6549 14059 6607 14065
rect 6549 14025 6561 14059
rect 6595 14056 6607 14059
rect 6914 14056 6920 14068
rect 6595 14028 6920 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7650 14056 7656 14068
rect 7515 14028 7656 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 7929 14059 7987 14065
rect 7929 14025 7941 14059
rect 7975 14056 7987 14059
rect 8478 14056 8484 14068
rect 7975 14028 8484 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 10778 14056 10784 14068
rect 9508 14028 10784 14056
rect 3878 13948 3884 14000
rect 3936 13988 3942 14000
rect 3973 13991 4031 13997
rect 3973 13988 3985 13991
rect 3936 13960 3985 13988
rect 3936 13948 3942 13960
rect 3973 13957 3985 13960
rect 4019 13957 4031 13991
rect 9508 13988 9536 14028
rect 10778 14016 10784 14028
rect 10836 14056 10842 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 10836 14028 10885 14056
rect 10836 14016 10842 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 12526 14056 12532 14068
rect 11563 14028 12532 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14056 15439 14059
rect 15470 14056 15476 14068
rect 15427 14028 15476 14056
rect 15427 14025 15439 14028
rect 15381 14019 15439 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 16850 14056 16856 14068
rect 16811 14028 16856 14056
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 25777 14059 25835 14065
rect 25777 14056 25789 14059
rect 19392 14028 25789 14056
rect 19392 14016 19398 14028
rect 25777 14025 25789 14028
rect 25823 14025 25835 14059
rect 25777 14019 25835 14025
rect 3973 13951 4031 13957
rect 8496 13960 9536 13988
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2590 13920 2596 13932
rect 1995 13892 2596 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2590 13880 2596 13892
rect 2648 13920 2654 13932
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2648 13892 2881 13920
rect 2648 13880 2654 13892
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 3050 13920 3056 13932
rect 2963 13892 3056 13920
rect 2869 13883 2927 13889
rect 3050 13880 3056 13892
rect 3108 13920 3114 13932
rect 4522 13920 4528 13932
rect 3108 13892 4528 13920
rect 3108 13880 3114 13892
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4982 13920 4988 13932
rect 4663 13892 4988 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 8496 13929 8524 13960
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 12618 13988 12624 14000
rect 11204 13960 12624 13988
rect 11204 13948 11210 13960
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 7883 13892 8493 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 12161 13923 12219 13929
rect 9447 13892 9628 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2332 13824 2789 13852
rect 1397 13787 1455 13793
rect 1397 13753 1409 13787
rect 1443 13784 1455 13787
rect 1486 13784 1492 13796
rect 1443 13756 1492 13784
rect 1443 13753 1455 13756
rect 1397 13747 1455 13753
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 2332 13728 2360 13824
rect 2777 13821 2789 13824
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3881 13855 3939 13861
rect 3559 13824 3832 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3804 13784 3832 13824
rect 3881 13821 3893 13855
rect 3927 13852 3939 13855
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 3927 13824 4445 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4433 13821 4445 13824
rect 4479 13852 4491 13855
rect 4890 13852 4896 13864
rect 4479 13824 4896 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 6178 13852 6184 13864
rect 5583 13824 6184 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 9490 13852 9496 13864
rect 9451 13824 9496 13852
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9600 13852 9628 13892
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12250 13920 12256 13932
rect 12207 13892 12256 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 15488 13920 15516 14016
rect 24305 13923 24363 13929
rect 13044 13892 13584 13920
rect 15488 13892 15608 13920
rect 13044 13880 13050 13892
rect 13556 13864 13584 13892
rect 9760 13855 9818 13861
rect 9760 13852 9772 13855
rect 9600 13824 9772 13852
rect 9760 13821 9772 13824
rect 9806 13852 9818 13855
rect 10134 13852 10140 13864
rect 9806 13824 10140 13852
rect 9806 13821 9818 13824
rect 9760 13815 9818 13821
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13170 13852 13176 13864
rect 13127 13824 13176 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 15378 13852 15384 13864
rect 13596 13824 15384 13852
rect 13596 13812 13602 13824
rect 15378 13812 15384 13824
rect 15436 13852 15442 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15436 13824 15485 13852
rect 15436 13812 15442 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15580 13852 15608 13892
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 24351 13892 24532 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 15729 13855 15787 13861
rect 15729 13852 15741 13855
rect 15580 13824 15741 13852
rect 15473 13815 15531 13821
rect 15729 13821 15741 13824
rect 15775 13852 15787 13855
rect 16482 13852 16488 13864
rect 15775 13824 16488 13852
rect 15775 13821 15787 13824
rect 15729 13815 15787 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 24394 13852 24400 13864
rect 24355 13824 24400 13852
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24504 13852 24532 13892
rect 24670 13861 24676 13864
rect 24664 13852 24676 13861
rect 24504 13824 24676 13852
rect 24664 13815 24676 13824
rect 24670 13812 24676 13815
rect 24728 13812 24734 13864
rect 3804 13756 4384 13784
rect 4356 13728 4384 13756
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 7374 13784 7380 13796
rect 6696 13756 7380 13784
rect 6696 13744 6702 13756
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 8297 13787 8355 13793
rect 8297 13753 8309 13787
rect 8343 13784 8355 13787
rect 11425 13787 11483 13793
rect 8343 13756 9076 13784
rect 8343 13753 8355 13756
rect 8297 13747 8355 13753
rect 9048 13728 9076 13756
rect 11425 13753 11437 13787
rect 11471 13784 11483 13787
rect 11885 13787 11943 13793
rect 11885 13784 11897 13787
rect 11471 13756 11897 13784
rect 11471 13753 11483 13756
rect 11425 13747 11483 13753
rect 11885 13753 11897 13756
rect 11931 13784 11943 13787
rect 12158 13784 12164 13796
rect 11931 13756 12164 13784
rect 11931 13753 11943 13756
rect 11885 13747 11943 13753
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 16500 13784 16528 13812
rect 17954 13784 17960 13796
rect 16500 13756 17960 13784
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 4338 13716 4344 13728
rect 4299 13688 4344 13716
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 4982 13716 4988 13728
rect 4943 13688 4988 13716
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 8386 13716 8392 13728
rect 8347 13688 8392 13716
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 9030 13716 9036 13728
rect 8991 13688 9036 13716
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 11974 13676 11980 13728
rect 12032 13716 12038 13728
rect 12032 13688 12077 13716
rect 12032 13676 12038 13688
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 12400 13688 14473 13716
rect 12400 13676 12406 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 1995 13484 2881 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2869 13481 2881 13484
rect 2915 13512 2927 13515
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2915 13484 4077 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 5813 13515 5871 13521
rect 5813 13481 5825 13515
rect 5859 13512 5871 13515
rect 6730 13512 6736 13524
rect 5859 13484 6736 13512
rect 5859 13481 5871 13484
rect 5813 13475 5871 13481
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7006 13512 7012 13524
rect 6963 13484 7012 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 7248 13484 7389 13512
rect 7248 13472 7254 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 7377 13475 7435 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 8938 13512 8944 13524
rect 8899 13484 8944 13512
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9088 13484 9689 13512
rect 9088 13472 9094 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 10042 13512 10048 13524
rect 10003 13484 10048 13512
rect 9677 13475 9735 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13512 11483 13515
rect 11974 13512 11980 13524
rect 11471 13484 11980 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11974 13472 11980 13484
rect 12032 13512 12038 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 12032 13484 12357 13512
rect 12032 13472 12038 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12345 13475 12403 13481
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 12802 13512 12808 13524
rect 12759 13484 12808 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 13538 13512 13544 13524
rect 13495 13484 13544 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 16390 13512 16396 13524
rect 15611 13484 16396 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 3050 13444 3056 13456
rect 2363 13416 3056 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 7837 13447 7895 13453
rect 7837 13444 7849 13447
rect 7208 13416 7849 13444
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 3881 13379 3939 13385
rect 3881 13345 3893 13379
rect 3927 13376 3939 13379
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 3927 13348 4445 13376
rect 3927 13345 3939 13348
rect 3881 13339 3939 13345
rect 4433 13345 4445 13348
rect 4479 13376 4491 13379
rect 4798 13376 4804 13388
rect 4479 13348 4804 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 2682 13308 2688 13320
rect 1443 13280 2688 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 2406 13240 2412 13252
rect 2367 13212 2412 13240
rect 2406 13200 2412 13212
rect 2464 13200 2470 13252
rect 2792 13240 2820 13339
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5534 13376 5540 13388
rect 5399 13348 5540 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 5534 13336 5540 13348
rect 5592 13376 5598 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 5592 13348 6193 13376
rect 5592 13336 5598 13348
rect 6181 13345 6193 13348
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7208 13385 7236 13416
rect 7837 13413 7849 13416
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 7193 13379 7251 13385
rect 7193 13376 7205 13379
rect 6972 13348 7205 13376
rect 6972 13336 6978 13348
rect 7193 13345 7205 13348
rect 7239 13345 7251 13379
rect 8772 13376 8800 13472
rect 12069 13447 12127 13453
rect 9140 13416 11744 13444
rect 9140 13385 9168 13416
rect 11716 13388 11744 13416
rect 12069 13413 12081 13447
rect 12115 13444 12127 13447
rect 12250 13444 12256 13456
rect 12115 13416 12256 13444
rect 12115 13413 12127 13416
rect 12069 13407 12127 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 16574 13404 16580 13456
rect 16632 13444 16638 13456
rect 16669 13447 16727 13453
rect 16669 13444 16681 13447
rect 16632 13416 16681 13444
rect 16632 13404 16638 13416
rect 16669 13413 16681 13416
rect 16715 13444 16727 13447
rect 17586 13444 17592 13456
rect 16715 13416 17592 13444
rect 16715 13413 16727 13416
rect 16669 13407 16727 13413
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 24394 13444 24400 13456
rect 24355 13416 24400 13444
rect 24394 13404 24400 13416
rect 24452 13404 24458 13456
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8772 13348 9137 13376
rect 7193 13339 7251 13345
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 11698 13376 11704 13388
rect 9732 13348 10824 13376
rect 11611 13348 11704 13376
rect 9732 13336 9738 13348
rect 10796 13320 10824 13348
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 12342 13376 12348 13388
rect 11756 13348 12348 13376
rect 11756 13336 11762 13348
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13376 12863 13379
rect 12986 13376 12992 13388
rect 12851 13348 12992 13376
rect 12851 13345 12863 13348
rect 12805 13339 12863 13345
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 15105 13379 15163 13385
rect 15105 13345 15117 13379
rect 15151 13376 15163 13379
rect 15746 13376 15752 13388
rect 15151 13348 15752 13376
rect 15151 13345 15163 13348
rect 15105 13339 15163 13345
rect 15746 13336 15752 13348
rect 15804 13376 15810 13388
rect 15933 13379 15991 13385
rect 15933 13376 15945 13379
rect 15804 13348 15945 13376
rect 15804 13336 15810 13348
rect 15933 13345 15945 13348
rect 15979 13345 15991 13379
rect 15933 13339 15991 13345
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4212 13280 4537 13308
rect 4212 13268 4218 13280
rect 4525 13277 4537 13280
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 4890 13308 4896 13320
rect 4755 13280 4896 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5721 13311 5779 13317
rect 5721 13277 5733 13311
rect 5767 13308 5779 13311
rect 5994 13308 6000 13320
rect 5767 13280 6000 13308
rect 5767 13277 5779 13280
rect 5721 13271 5779 13277
rect 5994 13268 6000 13280
rect 6052 13308 6058 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6052 13280 6285 13308
rect 6052 13268 6058 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 6420 13280 7941 13308
rect 6420 13268 6426 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9456 13280 10149 13308
rect 9456 13268 9462 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10318 13308 10324 13320
rect 10279 13280 10324 13308
rect 10137 13271 10195 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 12897 13271 12955 13277
rect 2792 13212 4108 13240
rect 4080 13184 4108 13212
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8481 13243 8539 13249
rect 8481 13240 8493 13243
rect 8444 13212 8493 13240
rect 8444 13200 8450 13212
rect 8481 13209 8493 13212
rect 8527 13240 8539 13243
rect 9582 13240 9588 13252
rect 8527 13212 9588 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 11514 13240 11520 13252
rect 11475 13212 11520 13240
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 12912 13240 12940 13271
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 16298 13308 16304 13320
rect 16255 13280 16304 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 12768 13212 12940 13240
rect 13464 13212 14473 13240
rect 12768 13200 12774 13212
rect 3510 13172 3516 13184
rect 3471 13144 3516 13172
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 4062 13132 4068 13184
rect 4120 13132 4126 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 9272 13144 9413 13172
rect 9272 13132 9278 13144
rect 9401 13141 9413 13144
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 13464 13172 13492 13212
rect 14461 13209 14473 13212
rect 14507 13240 14519 13243
rect 16758 13240 16764 13252
rect 14507 13212 16764 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 11112 13144 13492 13172
rect 11112 13132 11118 13144
rect 13538 13132 13544 13184
rect 13596 13172 13602 13184
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13596 13144 13737 13172
rect 13596 13132 13602 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 13964 13144 14105 13172
rect 13964 13132 13970 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1670 12968 1676 12980
rect 1627 12940 1676 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2958 12968 2964 12980
rect 2547 12940 2964 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 4948 12940 5825 12968
rect 4948 12928 4954 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 7374 12968 7380 12980
rect 7335 12940 7380 12968
rect 5813 12931 5871 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8662 12928 8668 12980
rect 8720 12928 8726 12980
rect 8846 12968 8852 12980
rect 8759 12940 8852 12968
rect 8846 12928 8852 12940
rect 8904 12968 8910 12980
rect 9306 12968 9312 12980
rect 8904 12940 9312 12968
rect 8904 12928 8910 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10100 12940 10609 12968
rect 10100 12928 10106 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 11609 12971 11667 12977
rect 11609 12937 11621 12971
rect 11655 12968 11667 12971
rect 11698 12968 11704 12980
rect 11655 12940 11704 12968
rect 11655 12937 11667 12940
rect 11609 12931 11667 12937
rect 11698 12928 11704 12940
rect 11756 12968 11762 12980
rect 11974 12968 11980 12980
rect 11756 12940 11980 12968
rect 11756 12928 11762 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12710 12968 12716 12980
rect 12299 12940 12716 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14884 12940 14933 12968
rect 14884 12928 14890 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 14921 12931 14979 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16080 12940 17141 12968
rect 16080 12928 16086 12940
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 17129 12931 17187 12937
rect 3973 12903 4031 12909
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 4522 12900 4528 12912
rect 4019 12872 4528 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 1544 12736 2605 12764
rect 1544 12724 1550 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 1412 12696 1440 12724
rect 2038 12696 2044 12708
rect 1412 12668 2044 12696
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 2133 12699 2191 12705
rect 2133 12665 2145 12699
rect 2179 12696 2191 12699
rect 2860 12699 2918 12705
rect 2860 12696 2872 12699
rect 2179 12668 2872 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 2860 12665 2872 12668
rect 2906 12696 2918 12699
rect 3142 12696 3148 12708
rect 2906 12668 3148 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 3988 12628 4016 12863
rect 4522 12860 4528 12872
rect 4580 12900 4586 12912
rect 4908 12900 4936 12928
rect 6638 12900 6644 12912
rect 4580 12872 4936 12900
rect 5451 12872 6644 12900
rect 4580 12860 4586 12872
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 5353 12835 5411 12841
rect 5353 12832 5365 12835
rect 5040 12804 5365 12832
rect 5040 12792 5046 12804
rect 5353 12801 5365 12804
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 4387 12736 5181 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 5169 12733 5181 12736
rect 5215 12764 5227 12767
rect 5258 12764 5264 12776
rect 5215 12736 5264 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 5368 12696 5396 12795
rect 4856 12668 5396 12696
rect 4856 12656 4862 12668
rect 2648 12600 4016 12628
rect 2648 12588 2654 12600
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4212 12600 4721 12628
rect 4212 12588 4218 12600
rect 4709 12597 4721 12600
rect 4755 12628 4767 12631
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4755 12600 5273 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5261 12597 5273 12600
rect 5307 12628 5319 12631
rect 5451 12628 5479 12872
rect 6638 12860 6644 12872
rect 6696 12900 6702 12912
rect 8680 12900 8708 12928
rect 10318 12900 10324 12912
rect 6696 12872 8708 12900
rect 10231 12872 10324 12900
rect 6696 12860 6702 12872
rect 10318 12860 10324 12872
rect 10376 12900 10382 12912
rect 10965 12903 11023 12909
rect 10965 12900 10977 12903
rect 10376 12872 10977 12900
rect 10376 12860 10382 12872
rect 10965 12869 10977 12872
rect 11011 12869 11023 12903
rect 16390 12900 16396 12912
rect 10965 12863 11023 12869
rect 16224 12872 16396 12900
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 8067 12804 8524 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 6914 12764 6920 12776
rect 6687 12736 6920 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 6914 12724 6920 12736
rect 6972 12764 6978 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 6972 12736 7757 12764
rect 6972 12724 6978 12736
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 7837 12699 7895 12705
rect 7837 12696 7849 12699
rect 7331 12668 7849 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7837 12665 7849 12668
rect 7883 12696 7895 12699
rect 7926 12696 7932 12708
rect 7883 12668 7932 12696
rect 7883 12665 7895 12668
rect 7837 12659 7895 12665
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8496 12705 8524 12804
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 8938 12832 8944 12844
rect 8720 12804 8944 12832
rect 8720 12792 8726 12804
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10336 12832 10364 12860
rect 10100 12804 10364 12832
rect 12713 12835 12771 12841
rect 10100 12792 10106 12804
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 12802 12832 12808 12844
rect 12759 12804 12808 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 13538 12832 13544 12844
rect 13499 12804 13544 12832
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 15562 12832 15568 12844
rect 15523 12804 15568 12832
rect 15562 12792 15568 12804
rect 15620 12832 15626 12844
rect 16224 12841 16252 12872
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 16761 12903 16819 12909
rect 16761 12900 16773 12903
rect 16540 12872 16773 12900
rect 16540 12860 16546 12872
rect 16761 12869 16773 12872
rect 16807 12869 16819 12903
rect 16761 12863 16819 12869
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15620 12804 16221 12832
rect 15620 12792 15626 12804
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16500 12832 16528 12860
rect 16347 12804 16528 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 9214 12773 9220 12776
rect 9208 12764 9220 12773
rect 9175 12736 9220 12764
rect 9208 12727 9220 12736
rect 9214 12724 9220 12727
rect 9272 12724 9278 12776
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 14734 12764 14740 12776
rect 14608 12736 14740 12764
rect 14608 12724 14614 12736
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 15335 12736 16129 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 16117 12733 16129 12736
rect 16163 12764 16175 12767
rect 17126 12764 17132 12776
rect 16163 12736 17132 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 8481 12699 8539 12705
rect 8481 12665 8493 12699
rect 8527 12696 8539 12699
rect 13449 12699 13507 12705
rect 8527 12668 8984 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 8956 12640 8984 12668
rect 13449 12665 13461 12699
rect 13495 12696 13507 12699
rect 13786 12699 13844 12705
rect 13786 12696 13798 12699
rect 13495 12668 13798 12696
rect 13495 12665 13507 12668
rect 13449 12659 13507 12665
rect 13786 12665 13798 12668
rect 13832 12696 13844 12699
rect 14090 12696 14096 12708
rect 13832 12668 14096 12696
rect 13832 12665 13844 12668
rect 13786 12659 13844 12665
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 5307 12600 5479 12628
rect 6273 12631 6331 12637
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 6273 12597 6285 12631
rect 6319 12628 6331 12631
rect 6362 12628 6368 12640
rect 6319 12600 6368 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 6362 12588 6368 12600
rect 6420 12628 6426 12640
rect 7006 12628 7012 12640
rect 6420 12600 7012 12628
rect 6420 12588 6426 12600
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 8938 12588 8944 12640
rect 8996 12588 9002 12640
rect 10778 12588 10784 12640
rect 10836 12628 10842 12640
rect 11054 12628 11060 12640
rect 10836 12600 11060 12628
rect 10836 12588 10842 12600
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 3016 12396 3157 12424
rect 3016 12384 3022 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3145 12387 3203 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4062 12424 4068 12436
rect 3975 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 5592 12396 5733 12424
rect 5592 12384 5598 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7064 12396 7205 12424
rect 7064 12384 7070 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 7193 12387 7251 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 12897 12427 12955 12433
rect 12897 12393 12909 12427
rect 12943 12393 12955 12427
rect 13538 12424 13544 12436
rect 13499 12396 13544 12424
rect 12897 12387 12955 12393
rect 1673 12359 1731 12365
rect 1673 12325 1685 12359
rect 1719 12356 1731 12359
rect 4080 12356 4108 12384
rect 1719 12328 4108 12356
rect 1719 12325 1731 12328
rect 1673 12319 1731 12325
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 6178 12356 6184 12368
rect 4580 12328 4752 12356
rect 6139 12328 6184 12356
rect 4580 12316 4586 12328
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1544 12260 1777 12288
rect 1544 12248 1550 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 2021 12291 2079 12297
rect 2021 12288 2033 12291
rect 1912 12260 2033 12288
rect 1912 12248 1918 12260
rect 2021 12257 2033 12260
rect 2067 12288 2079 12291
rect 2590 12288 2596 12300
rect 2067 12260 2596 12288
rect 2067 12257 2079 12260
rect 2021 12251 2079 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4028 12260 4445 12288
rect 4028 12248 4034 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4724 12232 4752 12328
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6917 12359 6975 12365
rect 6917 12325 6929 12359
rect 6963 12356 6975 12359
rect 7742 12356 7748 12368
rect 6963 12328 7748 12356
rect 6963 12325 6975 12328
rect 6917 12319 6975 12325
rect 7742 12316 7748 12328
rect 7800 12316 7806 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11762 12359 11820 12365
rect 11762 12356 11774 12359
rect 11572 12328 11774 12356
rect 11572 12316 11578 12328
rect 11762 12325 11774 12328
rect 11808 12325 11820 12359
rect 12912 12356 12940 12387
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 15013 12427 15071 12433
rect 15013 12424 15025 12427
rect 14700 12396 15025 12424
rect 14700 12384 14706 12396
rect 15013 12393 15025 12396
rect 15059 12424 15071 12427
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15059 12396 15761 12424
rect 15059 12393 15071 12396
rect 15013 12387 15071 12393
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 16298 12424 16304 12436
rect 16259 12396 16304 12424
rect 15749 12387 15807 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 17310 12424 17316 12436
rect 17223 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12424 17374 12436
rect 18598 12424 18604 12436
rect 17368 12396 18604 12424
rect 17368 12384 17374 12396
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 12986 12356 12992 12368
rect 12899 12328 12992 12356
rect 11762 12319 11820 12325
rect 12986 12316 12992 12328
rect 13044 12356 13050 12368
rect 13044 12328 14596 12356
rect 13044 12316 13050 12328
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6822 12288 6828 12300
rect 6135 12260 6828 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7644 12291 7702 12297
rect 7644 12257 7656 12291
rect 7690 12288 7702 12291
rect 8202 12288 8208 12300
rect 7690 12260 8208 12288
rect 7690 12257 7702 12260
rect 7644 12251 7702 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10686 12288 10692 12300
rect 10091 12260 10692 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 14568 12232 14596 12328
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 17221 12359 17279 12365
rect 17221 12356 17233 12359
rect 16724 12328 17233 12356
rect 16724 12316 16730 12328
rect 17221 12325 17233 12328
rect 17267 12325 17279 12359
rect 17221 12319 17279 12325
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14967 12260 15669 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15657 12257 15669 12260
rect 15703 12288 15715 12291
rect 15703 12260 16896 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4120 12192 4537 12220
rect 4120 12180 4126 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 4525 12183 4583 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 7374 12220 7380 12232
rect 6328 12192 6373 12220
rect 7335 12192 7380 12220
rect 6328 12180 6334 12192
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 5629 12155 5687 12161
rect 5629 12152 5641 12155
rect 5592 12124 5641 12152
rect 5592 12112 5598 12124
rect 5629 12121 5641 12124
rect 5675 12152 5687 12155
rect 6288 12152 6316 12180
rect 5675 12124 6316 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 10689 12155 10747 12161
rect 10689 12152 10701 12155
rect 10560 12124 10701 12152
rect 10560 12112 10566 12124
rect 10689 12121 10701 12124
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 2924 12056 3433 12084
rect 2924 12044 2930 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 3421 12047 3479 12053
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4856 12056 5089 12084
rect 4856 12044 4862 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12084 8815 12087
rect 9214 12084 9220 12096
rect 8803 12056 9220 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 9214 12044 9220 12056
rect 9272 12084 9278 12096
rect 9398 12084 9404 12096
rect 9272 12056 9404 12084
rect 9272 12044 9278 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10594 12084 10600 12096
rect 9732 12056 10600 12084
rect 9732 12044 9738 12056
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 11425 12087 11483 12093
rect 11425 12053 11437 12087
rect 11471 12084 11483 12087
rect 11532 12084 11560 12183
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 14608 12192 15853 12220
rect 14608 12180 14614 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 13538 12152 13544 12164
rect 13096 12124 13544 12152
rect 12250 12084 12256 12096
rect 11471 12056 12256 12084
rect 11471 12053 11483 12056
rect 11425 12047 11483 12053
rect 12250 12044 12256 12056
rect 12308 12084 12314 12096
rect 13096 12084 13124 12124
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 16868 12161 16896 12260
rect 17494 12220 17500 12232
rect 17455 12192 17500 12220
rect 17494 12180 17500 12192
rect 17552 12220 17558 12232
rect 17862 12220 17868 12232
rect 17552 12192 17868 12220
rect 17552 12180 17558 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 13262 12084 13268 12096
rect 12308 12056 13124 12084
rect 13223 12056 13268 12084
rect 12308 12044 12314 12056
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13906 12084 13912 12096
rect 13819 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12084 13970 12096
rect 14274 12084 14280 12096
rect 13964 12056 14280 12084
rect 13964 12044 13970 12056
rect 14274 12044 14280 12056
rect 14332 12084 14338 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14332 12056 14657 12084
rect 14332 12044 14338 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 14645 12047 14703 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14792 12056 14933 12084
rect 14792 12044 14798 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 15286 12084 15292 12096
rect 15247 12056 15292 12084
rect 14921 12047 14979 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 2832 11852 3433 11880
rect 2832 11840 2838 11852
rect 3421 11849 3433 11852
rect 3467 11880 3479 11883
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3467 11852 3709 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 4764 11852 5365 11880
rect 4764 11840 4770 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 5353 11843 5411 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 6822 11880 6828 11892
rect 6687 11852 6828 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7834 11880 7840 11892
rect 7616 11852 7840 11880
rect 7616 11840 7622 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 9309 11883 9367 11889
rect 9309 11849 9321 11883
rect 9355 11880 9367 11883
rect 10134 11880 10140 11892
rect 9355 11852 10140 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 10134 11840 10140 11852
rect 10192 11880 10198 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10192 11852 10701 11880
rect 10192 11840 10198 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 14090 11880 14096 11892
rect 14051 11852 14096 11880
rect 10689 11843 10747 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14550 11880 14556 11892
rect 14511 11852 14556 11880
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 16022 11880 16028 11892
rect 15427 11852 16028 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16482 11880 16488 11892
rect 16443 11852 16488 11880
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17310 11880 17316 11892
rect 17271 11852 17316 11880
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17589 11883 17647 11889
rect 17589 11880 17601 11883
rect 17552 11852 17601 11880
rect 17552 11840 17558 11852
rect 17589 11849 17601 11852
rect 17635 11849 17647 11883
rect 17589 11843 17647 11849
rect 3142 11812 3148 11824
rect 3103 11784 3148 11812
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 3970 11812 3976 11824
rect 3931 11784 3976 11812
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 8202 11812 8208 11824
rect 8163 11784 8208 11812
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 8849 11815 8907 11821
rect 8849 11781 8861 11815
rect 8895 11812 8907 11815
rect 10042 11812 10048 11824
rect 8895 11784 10048 11812
rect 8895 11781 8907 11784
rect 8849 11775 8907 11781
rect 10042 11772 10048 11784
rect 10100 11812 10106 11824
rect 10318 11812 10324 11824
rect 10100 11784 10324 11812
rect 10100 11772 10106 11784
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 13906 11772 13912 11824
rect 13964 11812 13970 11824
rect 14660 11812 14688 11840
rect 13964 11784 14688 11812
rect 13964 11772 13970 11784
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1544 11716 1777 11744
rect 1544 11704 1550 11716
rect 1765 11713 1777 11716
rect 1811 11713 1823 11747
rect 3160 11744 3188 11772
rect 3878 11744 3884 11756
rect 3160 11716 3884 11744
rect 1765 11707 1823 11713
rect 3878 11704 3884 11716
rect 3936 11744 3942 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 3936 11716 4537 11744
rect 3936 11704 3942 11716
rect 4525 11713 4537 11716
rect 4571 11744 4583 11747
rect 4798 11744 4804 11756
rect 4571 11716 4804 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4798 11704 4804 11716
rect 4856 11744 4862 11756
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4856 11716 4997 11744
rect 4856 11704 4862 11716
rect 4985 11713 4997 11716
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9456 11716 9873 11744
rect 9456 11704 9462 11716
rect 9861 11713 9873 11716
rect 9907 11713 9919 11747
rect 10502 11744 10508 11756
rect 9861 11707 9919 11713
rect 9968 11716 10508 11744
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 3743 11648 4353 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 4341 11639 4399 11645
rect 6822 11636 6828 11648
rect 6880 11676 6886 11688
rect 7374 11676 7380 11688
rect 6880 11648 7380 11676
rect 6880 11636 6886 11648
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9968 11676 9996 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16500 11744 16528 11840
rect 16071 11716 16528 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 8812 11648 9996 11676
rect 8812 11636 8818 11648
rect 10134 11636 10140 11688
rect 10192 11676 10198 11688
rect 10870 11676 10876 11688
rect 10192 11648 10876 11676
rect 10192 11636 10198 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 11848 11648 12173 11676
rect 11848 11636 11854 11648
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 12161 11639 12219 11645
rect 1673 11611 1731 11617
rect 1673 11577 1685 11611
rect 1719 11608 1731 11611
rect 2010 11611 2068 11617
rect 2010 11608 2022 11611
rect 1719 11580 2022 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 2010 11577 2022 11580
rect 2056 11608 2068 11611
rect 2314 11608 2320 11620
rect 2056 11580 2320 11608
rect 2056 11577 2068 11580
rect 2010 11571 2068 11577
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 7092 11611 7150 11617
rect 7092 11577 7104 11611
rect 7138 11608 7150 11611
rect 7466 11608 7472 11620
rect 7138 11580 7472 11608
rect 7138 11577 7150 11580
rect 7092 11571 7150 11577
rect 7466 11568 7472 11580
rect 7524 11568 7530 11620
rect 9398 11568 9404 11620
rect 9456 11608 9462 11620
rect 9766 11608 9772 11620
rect 9456 11580 9772 11608
rect 9456 11568 9462 11580
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 10100 11580 11345 11608
rect 10100 11568 10106 11580
rect 11333 11577 11345 11580
rect 11379 11577 11391 11611
rect 12176 11608 12204 11639
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12986 11685 12992 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12400 11648 12725 11676
rect 12400 11636 12406 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12980 11676 12992 11685
rect 12713 11639 12771 11645
rect 12912 11648 12992 11676
rect 12912 11608 12940 11648
rect 12980 11639 12992 11648
rect 12986 11636 12992 11639
rect 13044 11636 13050 11688
rect 15194 11608 15200 11620
rect 12176 11580 12940 11608
rect 15155 11580 15200 11608
rect 11333 11571 11391 11577
rect 15194 11568 15200 11580
rect 15252 11608 15258 11620
rect 15470 11608 15476 11620
rect 15252 11580 15476 11608
rect 15252 11568 15258 11580
rect 15470 11568 15476 11580
rect 15528 11608 15534 11620
rect 15749 11611 15807 11617
rect 15749 11608 15761 11611
rect 15528 11580 15761 11608
rect 15528 11568 15534 11580
rect 15749 11577 15761 11580
rect 15795 11577 15807 11611
rect 15749 11571 15807 11577
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3789 11543 3847 11549
rect 3789 11540 3801 11543
rect 3108 11512 3801 11540
rect 3108 11500 3114 11512
rect 3789 11509 3801 11512
rect 3835 11540 3847 11543
rect 4246 11540 4252 11552
rect 3835 11512 4252 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4246 11500 4252 11512
rect 4304 11540 4310 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4304 11512 4445 11540
rect 4304 11500 4310 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 4433 11503 4491 11509
rect 5721 11543 5779 11549
rect 5721 11509 5733 11543
rect 5767 11540 5779 11543
rect 6086 11540 6092 11552
rect 5767 11512 6092 11540
rect 5767 11509 5779 11512
rect 5721 11503 5779 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 9217 11543 9275 11549
rect 9217 11509 9229 11543
rect 9263 11540 9275 11543
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9263 11512 9689 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 9677 11509 9689 11512
rect 9723 11540 9735 11543
rect 10134 11540 10140 11552
rect 9723 11512 10140 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10686 11540 10692 11552
rect 10459 11512 10692 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11572 11512 11805 11540
rect 11572 11500 11578 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 14921 11543 14979 11549
rect 14921 11509 14933 11543
rect 14967 11540 14979 11543
rect 15102 11540 15108 11552
rect 14967 11512 15108 11540
rect 14967 11509 14979 11512
rect 14921 11503 14979 11509
rect 15102 11500 15108 11512
rect 15160 11540 15166 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15160 11512 15853 11540
rect 15160 11500 15166 11512
rect 15841 11509 15853 11512
rect 15887 11509 15899 11543
rect 15841 11503 15899 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16724 11512 16865 11540
rect 16724 11500 16730 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 16853 11503 16911 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4062 11336 4068 11348
rect 3927 11308 4068 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5629 11339 5687 11345
rect 5629 11305 5641 11339
rect 5675 11336 5687 11339
rect 5994 11336 6000 11348
rect 5675 11308 6000 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 7469 11339 7527 11345
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 8202 11336 8208 11348
rect 7515 11308 8208 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 11146 11336 11152 11348
rect 9723 11308 11152 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 13446 11336 13452 11348
rect 12851 11308 13452 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14734 11336 14740 11348
rect 14695 11308 14740 11336
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 15151 11308 15761 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15749 11305 15761 11308
rect 15795 11336 15807 11339
rect 16853 11339 16911 11345
rect 16853 11336 16865 11339
rect 15795 11308 16865 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16853 11305 16865 11308
rect 16899 11305 16911 11339
rect 16853 11299 16911 11305
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 17310 11336 17316 11348
rect 17267 11308 17316 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 1578 11228 1584 11280
rect 1636 11268 1642 11280
rect 2498 11268 2504 11280
rect 1636 11240 2504 11268
rect 1636 11228 1642 11240
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 3513 11271 3571 11277
rect 3513 11237 3525 11271
rect 3559 11268 3571 11271
rect 3970 11268 3976 11280
rect 3559 11240 3976 11268
rect 3559 11237 3571 11240
rect 3513 11231 3571 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4430 11268 4436 11280
rect 4343 11240 4436 11268
rect 4430 11228 4436 11240
rect 4488 11268 4494 11280
rect 4706 11268 4712 11280
rect 4488 11240 4712 11268
rect 4488 11228 4494 11240
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 8478 11268 8484 11280
rect 8439 11240 8484 11268
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 11164 11268 11192 11296
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 11164 11240 11621 11268
rect 11609 11237 11621 11240
rect 11655 11237 11667 11271
rect 11609 11231 11667 11237
rect 13173 11271 13231 11277
rect 13173 11237 13185 11271
rect 13219 11268 13231 11271
rect 13262 11268 13268 11280
rect 13219 11240 13268 11268
rect 13219 11237 13231 11240
rect 13173 11231 13231 11237
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 4246 11200 4252 11212
rect 3844 11172 4252 11200
rect 3844 11160 3850 11172
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5592 11172 6009 11200
rect 5592 11160 5598 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11200 6147 11203
rect 6362 11200 6368 11212
rect 6135 11172 6368 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 8386 11200 8392 11212
rect 7800 11172 8392 11200
rect 7800 11160 7806 11172
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 9582 11200 9588 11212
rect 8496 11172 9588 11200
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 2593 11095 2651 11101
rect 4356 11104 4537 11132
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 2406 11064 2412 11076
rect 2087 11036 2412 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 2608 10996 2636 11095
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 3053 11067 3111 11073
rect 3053 11064 3065 11067
rect 2740 11036 3065 11064
rect 2740 11024 2746 11036
rect 3053 11033 3065 11036
rect 3099 11033 3111 11067
rect 3053 11027 3111 11033
rect 4356 11008 4384 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4798 11132 4804 11144
rect 4755 11104 4804 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5307 11036 5580 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 2556 10968 2636 10996
rect 2556 10956 2562 10968
rect 4338 10956 4344 11008
rect 4396 10956 4402 11008
rect 5552 10996 5580 11036
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 7834 11064 7840 11076
rect 7432 11036 7696 11064
rect 7795 11036 7840 11064
rect 7432 11024 7438 11036
rect 5994 10996 6000 11008
rect 5552 10968 6000 10996
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7466 10996 7472 11008
rect 6963 10968 7472 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7668 10996 7696 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8496 11064 8524 11172
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 10376 11172 12633 11200
rect 10376 11160 10382 11172
rect 12621 11169 12633 11172
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8067 11036 8524 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8588 10996 8616 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9916 11104 10149 11132
rect 9916 11092 9922 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11132 10287 11135
rect 11514 11132 11520 11144
rect 10275 11104 11520 11132
rect 10275 11101 10287 11104
rect 10229 11095 10287 11101
rect 10244 11064 10272 11095
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11698 11132 11704 11144
rect 11659 11104 11704 11132
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 11848 11104 11893 11132
rect 11848 11092 11854 11104
rect 9600 11036 10272 11064
rect 10873 11067 10931 11073
rect 9398 10996 9404 11008
rect 7668 10968 9404 10996
rect 9398 10956 9404 10968
rect 9456 10996 9462 11008
rect 9600 10996 9628 11036
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 10962 11064 10968 11076
rect 10919 11036 10968 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 10962 11024 10968 11036
rect 11020 11064 11026 11076
rect 11241 11067 11299 11073
rect 11020 11036 11100 11064
rect 11020 11024 11026 11036
rect 9456 10968 9628 10996
rect 11072 10996 11100 11036
rect 11241 11033 11253 11067
rect 11287 11064 11299 11067
rect 13188 11064 13216 11231
rect 13262 11228 13268 11240
rect 13320 11228 13326 11280
rect 14274 11228 14280 11280
rect 14332 11268 14338 11280
rect 16574 11268 16580 11280
rect 14332 11240 16580 11268
rect 14332 11228 14338 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 16758 11268 16764 11280
rect 16719 11240 16764 11268
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 15378 11200 15384 11212
rect 14056 11172 15384 11200
rect 14056 11160 14062 11172
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15620 11172 15669 11200
rect 15620 11160 15626 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11200 17371 11203
rect 17586 11200 17592 11212
rect 17359 11172 17592 11200
rect 17359 11169 17371 11172
rect 17313 11163 17371 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13354 11132 13360 11144
rect 13311 11104 13360 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13538 11132 13544 11144
rect 13495 11104 13544 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 13538 11092 13544 11104
rect 13596 11132 13602 11144
rect 14090 11132 14096 11144
rect 13596 11104 14096 11132
rect 13596 11092 13602 11104
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 17494 11132 17500 11144
rect 17455 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 11287 11036 13216 11064
rect 15289 11067 15347 11073
rect 11287 11033 11299 11036
rect 11241 11027 11299 11033
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 16206 11064 16212 11076
rect 15335 11036 16212 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 11146 10996 11152 11008
rect 11072 10968 11152 10996
rect 9456 10956 9462 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 12526 10996 12532 11008
rect 12487 10968 12532 10996
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12621 10999 12679 11005
rect 12621 10965 12633 10999
rect 12667 10996 12679 10999
rect 13998 10996 14004 11008
rect 12667 10968 14004 10996
rect 12667 10965 12679 10968
rect 12621 10959 12679 10965
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 14093 10999 14151 11005
rect 14093 10965 14105 10999
rect 14139 10996 14151 10999
rect 14274 10996 14280 11008
rect 14139 10968 14280 10996
rect 14139 10965 14151 10968
rect 14093 10959 14151 10965
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 16114 10956 16120 11008
rect 16172 10996 16178 11008
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 16172 10968 16313 10996
rect 16172 10956 16178 10968
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1394 10792 1400 10804
rect 1307 10764 1400 10792
rect 1394 10752 1400 10764
rect 1452 10792 1458 10804
rect 2774 10792 2780 10804
rect 1452 10764 2780 10792
rect 1452 10752 1458 10764
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 2958 10792 2964 10804
rect 2915 10764 2964 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6328 10764 6561 10792
rect 6328 10752 6334 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 6549 10755 6607 10761
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7432 10764 7481 10792
rect 7432 10752 7438 10764
rect 7469 10761 7481 10764
rect 7515 10761 7527 10795
rect 10042 10792 10048 10804
rect 10003 10764 10048 10792
rect 7469 10755 7527 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12124 10764 12173 10792
rect 12124 10752 12130 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 13538 10792 13544 10804
rect 13499 10764 13544 10792
rect 12161 10755 12219 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17310 10792 17316 10804
rect 16991 10764 17316 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 1946 10656 1952 10668
rect 1907 10628 1952 10656
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 2976 10656 3004 10752
rect 5442 10684 5448 10736
rect 5500 10724 5506 10736
rect 7742 10724 7748 10736
rect 5500 10696 7748 10724
rect 5500 10684 5506 10696
rect 7742 10684 7748 10696
rect 7800 10724 7806 10736
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 7800 10696 7849 10724
rect 7800 10684 7806 10696
rect 7837 10693 7849 10696
rect 7883 10693 7895 10727
rect 7837 10687 7895 10693
rect 9401 10727 9459 10733
rect 9401 10693 9413 10727
rect 9447 10724 9459 10727
rect 9950 10724 9956 10736
rect 9447 10696 9956 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 16960 10724 16988 10755
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 12860 10696 16988 10724
rect 12860 10684 12866 10696
rect 5813 10659 5871 10665
rect 2976 10628 3096 10656
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2832 10560 2973 10588
rect 2832 10548 2838 10560
rect 2961 10557 2973 10560
rect 3007 10557 3019 10591
rect 3068 10588 3096 10628
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6086 10656 6092 10668
rect 5859 10628 6092 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9824 10628 10609 10656
rect 9824 10616 9830 10628
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 11422 10656 11428 10668
rect 10643 10628 11192 10656
rect 11335 10628 11428 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 3217 10591 3275 10597
rect 3217 10588 3229 10591
rect 3068 10560 3229 10588
rect 2961 10551 3019 10557
rect 3217 10557 3229 10560
rect 3263 10557 3275 10591
rect 3217 10551 3275 10557
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4396 10560 4629 10588
rect 4396 10548 4402 10560
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 4617 10551 4675 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 7116 10588 7144 10616
rect 8018 10588 8024 10600
rect 5675 10560 7144 10588
rect 7979 10560 8024 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8288 10591 8346 10597
rect 8288 10557 8300 10591
rect 8334 10588 8346 10591
rect 8570 10588 8576 10600
rect 8334 10560 8576 10588
rect 8334 10557 8346 10560
rect 8288 10551 8346 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 11164 10597 11192 10628
rect 11422 10616 11428 10628
rect 11480 10656 11486 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11480 10628 11897 10656
rect 11480 10616 11486 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 12986 10656 12992 10668
rect 11931 10628 12992 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10656 13967 10659
rect 14550 10656 14556 10668
rect 13955 10628 14556 10656
rect 13955 10625 13967 10628
rect 13909 10619 13967 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 16114 10656 16120 10668
rect 16075 10628 16120 10656
rect 16114 10616 16120 10628
rect 16172 10656 16178 10668
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 16172 10628 17233 10656
rect 16172 10616 16178 10628
rect 17221 10625 17233 10628
rect 17267 10656 17279 10659
rect 17494 10656 17500 10668
rect 17267 10628 17500 10656
rect 17267 10625 17279 10628
rect 17221 10619 17279 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12584 10560 12817 10588
rect 12584 10548 12590 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 15194 10588 15200 10600
rect 14424 10560 15200 10588
rect 14424 10548 14430 10560
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15436 10560 16037 10588
rect 15436 10548 15442 10560
rect 16025 10557 16037 10560
rect 16071 10588 16083 10591
rect 16071 10560 16160 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 16132 10532 16160 10560
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2682 10520 2688 10532
rect 1903 10492 2688 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2682 10480 2688 10492
rect 2740 10480 2746 10532
rect 12066 10480 12072 10532
rect 12124 10520 12130 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12124 10492 12909 10520
rect 12124 10480 12130 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 14461 10523 14519 10529
rect 14461 10520 14473 10523
rect 13872 10492 14473 10520
rect 13872 10480 13878 10492
rect 14461 10489 14473 10492
rect 14507 10489 14519 10523
rect 15010 10520 15016 10532
rect 14971 10492 15016 10520
rect 14461 10483 14519 10489
rect 15010 10480 15016 10492
rect 15068 10520 15074 10532
rect 15933 10523 15991 10529
rect 15933 10520 15945 10523
rect 15068 10492 15945 10520
rect 15068 10480 15074 10492
rect 15933 10489 15945 10492
rect 15979 10489 15991 10523
rect 15933 10483 15991 10489
rect 16114 10480 16120 10532
rect 16172 10480 16178 10532
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 2222 10452 2228 10464
rect 1811 10424 2228 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4614 10452 4620 10464
rect 4387 10424 4620 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4706 10412 4712 10464
rect 4764 10452 4770 10464
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4764 10424 4997 10452
rect 4764 10412 4770 10424
rect 4985 10421 4997 10424
rect 5031 10421 5043 10455
rect 6270 10452 6276 10464
rect 6231 10424 6276 10452
rect 4985 10415 5043 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 9769 10455 9827 10461
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 9858 10452 9864 10464
rect 9815 10424 9864 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10778 10452 10784 10464
rect 10739 10424 10784 10452
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 14001 10455 14059 10461
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14090 10452 14096 10464
rect 14047 10424 14096 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14332 10424 14381 10452
rect 14332 10412 14338 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 14369 10415 14427 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 17586 10452 17592 10464
rect 17547 10424 17592 10452
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2682 10248 2688 10260
rect 2455 10220 2688 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3510 10248 3516 10260
rect 2823 10220 3516 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3510 10208 3516 10220
rect 3568 10248 3574 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3568 10220 4077 10248
rect 3568 10208 3574 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 7466 10248 7472 10260
rect 7427 10220 7472 10248
rect 4065 10211 4123 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 11422 10248 11428 10260
rect 11383 10220 11428 10248
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11790 10248 11796 10260
rect 11751 10220 11796 10248
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 15562 10248 15568 10260
rect 14783 10220 15568 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 16758 10248 16764 10260
rect 16719 10220 16764 10248
rect 16758 10208 16764 10220
rect 16816 10248 16822 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16816 10220 17049 10248
rect 16816 10208 16822 10220
rect 17037 10217 17049 10220
rect 17083 10248 17095 10251
rect 17862 10248 17868 10260
rect 17083 10220 17868 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 2280 10152 3433 10180
rect 2280 10140 2286 10152
rect 3421 10149 3433 10152
rect 3467 10149 3479 10183
rect 3878 10180 3884 10192
rect 3839 10152 3884 10180
rect 3421 10143 3479 10149
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 4433 10183 4491 10189
rect 4433 10149 4445 10183
rect 4479 10180 4491 10183
rect 4522 10180 4528 10192
rect 4479 10152 4528 10180
rect 4479 10149 4491 10152
rect 4433 10143 4491 10149
rect 4522 10140 4528 10152
rect 4580 10180 4586 10192
rect 4982 10180 4988 10192
rect 4580 10152 4988 10180
rect 4580 10140 4586 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 6822 10180 6828 10192
rect 6104 10152 6828 10180
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2869 10115 2927 10121
rect 2869 10112 2881 10115
rect 2363 10084 2881 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2869 10081 2881 10084
rect 2915 10112 2927 10115
rect 4062 10112 4068 10124
rect 2915 10084 4068 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 5626 10112 5632 10124
rect 5587 10084 5632 10112
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6104 10121 6132 10152
rect 6822 10140 6828 10152
rect 6880 10180 6886 10192
rect 8018 10180 8024 10192
rect 6880 10152 8024 10180
rect 6880 10140 6886 10152
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 14090 10180 14096 10192
rect 13780 10152 14096 10180
rect 13780 10140 13786 10152
rect 14090 10140 14096 10152
rect 14148 10140 14154 10192
rect 14642 10140 14648 10192
rect 14700 10180 14706 10192
rect 15013 10183 15071 10189
rect 15013 10180 15025 10183
rect 14700 10152 15025 10180
rect 14700 10140 14706 10152
rect 15013 10149 15025 10152
rect 15059 10149 15071 10183
rect 16022 10180 16028 10192
rect 15013 10143 15071 10149
rect 15488 10152 16028 10180
rect 6362 10121 6368 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 6052 10084 6101 10112
rect 6052 10072 6058 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6356 10112 6368 10121
rect 6323 10084 6368 10112
rect 6089 10075 6147 10081
rect 6356 10075 6368 10084
rect 6362 10072 6368 10075
rect 6420 10072 6426 10124
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7800 10084 8125 10112
rect 7800 10072 7806 10084
rect 8113 10081 8125 10084
rect 8159 10112 8171 10115
rect 8478 10112 8484 10124
rect 8159 10084 8484 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9766 10112 9772 10124
rect 8619 10084 9772 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 9950 10121 9956 10124
rect 9944 10112 9956 10121
rect 9911 10084 9956 10112
rect 9944 10075 9956 10084
rect 9950 10072 9956 10075
rect 10008 10072 10014 10124
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12158 10112 12164 10124
rect 12032 10084 12164 10112
rect 12032 10072 12038 10084
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12342 10112 12348 10124
rect 12268 10084 12348 10112
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2130 10044 2136 10056
rect 1443 10016 2136 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3142 10044 3148 10056
rect 3099 10016 3148 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4488 10016 4537 10044
rect 4488 10004 4494 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4672 10016 4717 10044
rect 4672 10004 4678 10016
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 12268 10053 12296 10084
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12520 10115 12578 10121
rect 12520 10081 12532 10115
rect 12566 10112 12578 10115
rect 12986 10112 12992 10124
rect 12566 10084 12992 10112
rect 12566 10081 12578 10084
rect 12520 10075 12578 10081
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 9732 10016 9777 10044
rect 11992 10016 12265 10044
rect 9732 10004 9738 10016
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5258 9908 5264 9920
rect 5215 9880 5264 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11992 9917 12020 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15488 10044 15516 10152
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15620 10084 15669 10112
rect 15620 10072 15626 10084
rect 15657 10081 15669 10084
rect 15703 10112 15715 10115
rect 16482 10112 16488 10124
rect 15703 10084 16488 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15436 10016 15761 10044
rect 15436 10004 15442 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 15896 10016 15941 10044
rect 15896 10004 15902 10016
rect 15289 9979 15347 9985
rect 15289 9945 15301 9979
rect 15335 9976 15347 9979
rect 17586 9976 17592 9988
rect 15335 9948 17592 9976
rect 15335 9945 15347 9948
rect 15289 9939 15347 9945
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11204 9880 11989 9908
rect 11204 9868 11210 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 13633 9911 13691 9917
rect 13633 9908 13645 9911
rect 13504 9880 13645 9908
rect 13504 9868 13510 9880
rect 13633 9877 13645 9880
rect 13679 9877 13691 9911
rect 13633 9871 13691 9877
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13872 9880 14013 9908
rect 13872 9868 13878 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 14001 9871 14059 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 7190 9704 7196 9716
rect 6788 9676 7196 9704
rect 6788 9664 6794 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 13446 9704 13452 9716
rect 13407 9676 13452 9704
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14608 9676 14933 9704
rect 14608 9664 14614 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 18506 9704 18512 9716
rect 17000 9676 18184 9704
rect 17000 9664 17006 9676
rect 2682 9636 2688 9648
rect 2643 9608 2688 9636
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4212 9608 4997 9636
rect 4212 9596 4218 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6604 9608 6837 9636
rect 6604 9596 6610 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 7484 9608 10180 9636
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 7484 9577 7512 9608
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 4672 9540 5549 9568
rect 4672 9528 4678 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 6687 9540 7481 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 7469 9531 7527 9537
rect 7852 9540 8861 9568
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2774 9460 2780 9512
rect 2832 9509 2838 9512
rect 3050 9509 3056 9512
rect 2832 9500 2842 9509
rect 3044 9500 3056 9509
rect 2832 9472 2877 9500
rect 3011 9472 3056 9500
rect 2832 9463 2842 9472
rect 3044 9463 3056 9472
rect 2832 9460 2838 9463
rect 3050 9460 3056 9463
rect 3108 9460 3114 9512
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 6914 9500 6920 9512
rect 3476 9472 6920 9500
rect 3476 9460 3482 9472
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7852 9509 7880 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9568 8999 9571
rect 10152 9568 10180 9608
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11756 9608 11805 9636
rect 11756 9596 11762 9608
rect 11793 9605 11805 9608
rect 11839 9605 11851 9639
rect 12250 9636 12256 9648
rect 12211 9608 12256 9636
rect 11793 9599 11851 9605
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12437 9571 12495 9577
rect 8987 9540 9720 9568
rect 10152 9540 10272 9568
rect 8987 9537 8999 9540
rect 8941 9531 8999 9537
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 7248 9472 7849 9500
rect 7248 9460 7254 9472
rect 7837 9469 7849 9472
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8297 9503 8355 9509
rect 8297 9469 8309 9503
rect 8343 9500 8355 9503
rect 8757 9503 8815 9509
rect 8343 9472 8708 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 6181 9435 6239 9441
rect 3660 9404 6132 9432
rect 3660 9392 3666 9404
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 1728 9336 2329 9364
rect 1728 9324 1734 9336
rect 2317 9333 2329 9336
rect 2363 9364 2375 9367
rect 3142 9364 3148 9376
rect 2363 9336 3148 9364
rect 2363 9333 2375 9336
rect 2317 9327 2375 9333
rect 3142 9324 3148 9336
rect 3200 9364 3206 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3200 9336 4169 9364
rect 3200 9324 3206 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4430 9364 4436 9376
rect 4391 9336 4436 9364
rect 4157 9327 4215 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4580 9336 4813 9364
rect 4580 9324 4586 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 4801 9327 4859 9333
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 5316 9336 5365 9364
rect 5316 9324 5322 9336
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5353 9327 5411 9333
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 6104 9364 6132 9404
rect 6181 9401 6193 9435
rect 6227 9432 6239 9435
rect 6362 9432 6368 9444
rect 6227 9404 6368 9432
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 6362 9392 6368 9404
rect 6420 9432 6426 9444
rect 7098 9432 7104 9444
rect 6420 9404 7104 9432
rect 6420 9392 6426 9404
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 8680 9432 8708 9472
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9030 9500 9036 9512
rect 8803 9472 9036 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9140 9432 9168 9540
rect 9692 9441 9720 9540
rect 10134 9500 10140 9512
rect 10095 9472 10140 9500
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10244 9500 10272 9540
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 12526 9568 12532 9580
rect 12483 9540 12532 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 13464 9568 13492 9664
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 15565 9639 15623 9645
rect 15565 9636 15577 9639
rect 15528 9608 15577 9636
rect 15528 9596 15534 9608
rect 15565 9605 15577 9608
rect 15611 9605 15623 9639
rect 15565 9599 15623 9605
rect 13464 9540 13676 9568
rect 10404 9503 10462 9509
rect 10404 9500 10416 9503
rect 10244 9472 10416 9500
rect 10404 9469 10416 9472
rect 10450 9500 10462 9503
rect 10962 9500 10968 9512
rect 10450 9472 10968 9500
rect 10450 9469 10462 9472
rect 10404 9463 10462 9469
rect 8680 9404 9168 9432
rect 9677 9435 9735 9441
rect 9677 9401 9689 9435
rect 9723 9432 9735 9435
rect 10045 9435 10103 9441
rect 9723 9404 9976 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 9948 9376 9976 9404
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 10419 9432 10447 9463
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13648 9500 13676 9540
rect 13797 9503 13855 9509
rect 13797 9500 13809 9503
rect 13648 9472 13809 9500
rect 13797 9469 13809 9472
rect 13843 9469 13855 9503
rect 15580 9500 15608 9599
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16632 9608 16773 9636
rect 16632 9596 16638 9608
rect 16761 9605 16773 9608
rect 16807 9605 16819 9639
rect 16761 9599 16819 9605
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18156 9636 18184 9676
rect 18104 9608 18184 9636
rect 18248 9676 18512 9704
rect 18104 9596 18110 9608
rect 18248 9580 18276 9676
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 16298 9568 16304 9580
rect 16259 9540 16304 9568
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 15580 9472 16129 9500
rect 13797 9463 13855 9469
rect 16117 9469 16129 9472
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 10091 9404 10447 9432
rect 15304 9404 16221 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 15304 9376 15332 9404
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 16209 9395 16267 9401
rect 7006 9364 7012 9376
rect 5500 9336 5545 9364
rect 6104 9336 7012 9364
rect 5500 9324 5506 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 8018 9364 8024 9376
rect 7331 9336 8024 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 8018 9324 8024 9336
rect 8076 9364 8082 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 8076 9336 8401 9364
rect 8076 9324 8082 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 9930 9324 9936 9376
rect 9988 9324 9994 9376
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11112 9336 11529 9364
rect 11112 9324 11118 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 12986 9364 12992 9376
rect 12947 9336 12992 9364
rect 11517 9327 11575 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 15286 9364 15292 9376
rect 15247 9336 15292 9364
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17221 9367 17279 9373
rect 17221 9364 17233 9367
rect 16724 9336 17233 9364
rect 16724 9324 16730 9336
rect 17221 9333 17233 9336
rect 17267 9364 17279 9367
rect 17494 9364 17500 9376
rect 17267 9336 17500 9364
rect 17267 9333 17279 9336
rect 17221 9327 17279 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9364 17647 9367
rect 17862 9364 17868 9376
rect 17635 9336 17868 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2004 9132 2789 9160
rect 2004 9120 2010 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 2777 9123 2835 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4614 9160 4620 9172
rect 4448 9132 4620 9160
rect 1670 9101 1676 9104
rect 1664 9092 1676 9101
rect 1631 9064 1676 9092
rect 1664 9055 1676 9064
rect 1670 9052 1676 9055
rect 1728 9052 1734 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3108 9064 3801 9092
rect 3108 9052 3114 9064
rect 3789 9061 3801 9064
rect 3835 9092 3847 9095
rect 4448 9092 4476 9132
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 7650 9160 7656 9172
rect 6840 9132 7656 9160
rect 3835 9064 4476 9092
rect 4525 9095 4583 9101
rect 3835 9061 3847 9064
rect 3789 9055 3847 9061
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4890 9092 4896 9104
rect 4571 9064 4896 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 4890 9052 4896 9064
rect 4948 9092 4954 9104
rect 6840 9092 6868 9132
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8018 9160 8024 9172
rect 7975 9132 8024 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 4948 9064 6868 9092
rect 4948 9052 4954 9064
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 9401 9095 9459 9101
rect 9401 9092 9413 9095
rect 7248 9064 9413 9092
rect 7248 9052 7254 9064
rect 9401 9061 9413 9064
rect 9447 9092 9459 9095
rect 9692 9092 9720 9123
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 9824 9132 10057 9160
rect 9824 9120 9830 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 12345 9163 12403 9169
rect 12345 9129 12357 9163
rect 12391 9160 12403 9163
rect 12434 9160 12440 9172
rect 12391 9132 12440 9160
rect 12391 9129 12403 9132
rect 12345 9123 12403 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12894 9160 12900 9172
rect 12855 9132 12900 9160
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 16761 9163 16819 9169
rect 16761 9160 16773 9163
rect 16356 9132 16773 9160
rect 16356 9120 16362 9132
rect 16761 9129 16773 9132
rect 16807 9160 16819 9163
rect 16942 9160 16948 9172
rect 16807 9132 16948 9160
rect 16807 9129 16819 9132
rect 16761 9123 16819 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 9447 9064 9720 9092
rect 10137 9095 10195 9101
rect 9447 9061 9459 9064
rect 9401 9055 9459 9061
rect 10137 9061 10149 9095
rect 10183 9061 10195 9095
rect 10137 9055 10195 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1486 9024 1492 9036
rect 1443 8996 1492 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1486 8984 1492 8996
rect 1544 9024 1550 9036
rect 2774 9024 2780 9036
rect 1544 8996 2780 9024
rect 1544 8984 1550 8996
rect 2774 8984 2780 8996
rect 2832 8984 2838 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4798 9024 4804 9036
rect 4479 8996 4804 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 5902 9024 5908 9036
rect 5859 8996 5908 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6080 9027 6138 9033
rect 6080 8993 6092 9027
rect 6126 9024 6138 9027
rect 6454 9024 6460 9036
rect 6126 8996 6460 9024
rect 6126 8993 6138 8996
rect 6080 8987 6138 8993
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 8018 9024 8024 9036
rect 7064 8996 8024 9024
rect 7064 8984 7070 8996
rect 8018 8984 8024 8996
rect 8076 9024 8082 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8076 8996 8401 9024
rect 8076 8984 8082 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 10152 9024 10180 9055
rect 10410 9052 10416 9104
rect 10468 9092 10474 9104
rect 11146 9092 11152 9104
rect 10468 9064 11152 9092
rect 10468 9052 10474 9064
rect 11146 9052 11152 9064
rect 11204 9092 11210 9104
rect 13449 9095 13507 9101
rect 13449 9092 13461 9095
rect 11204 9064 13461 9092
rect 11204 9052 11210 9064
rect 13449 9061 13461 9064
rect 13495 9092 13507 9095
rect 13538 9092 13544 9104
rect 13495 9064 13544 9092
rect 13495 9061 13507 9064
rect 13449 9055 13507 9061
rect 13538 9052 13544 9064
rect 13596 9092 13602 9104
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 13596 9064 13829 9092
rect 13596 9052 13602 9064
rect 13817 9061 13829 9064
rect 13863 9092 13875 9095
rect 14182 9092 14188 9104
rect 13863 9064 14188 9092
rect 13863 9061 13875 9064
rect 13817 9055 13875 9061
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 10778 9024 10784 9036
rect 8389 8987 8447 8993
rect 10060 8996 10180 9024
rect 10739 8996 10784 9024
rect 4614 8956 4620 8968
rect 4575 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8956 4678 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 4672 8928 5457 8956
rect 4672 8916 4678 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7926 8956 7932 8968
rect 6972 8928 7932 8956
rect 6972 8916 6978 8928
rect 7926 8916 7932 8928
rect 7984 8956 7990 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 7984 8928 8493 8956
rect 7984 8916 7990 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8628 8928 9045 8956
rect 8628 8916 8634 8928
rect 9033 8925 9045 8928
rect 9079 8956 9091 8959
rect 9122 8956 9128 8968
rect 9079 8928 9128 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 8021 8891 8079 8897
rect 8021 8857 8033 8891
rect 8067 8888 8079 8891
rect 10060 8888 10088 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12492 8996 12817 9024
rect 12492 8984 12498 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 15286 9024 15292 9036
rect 13044 8996 15292 9024
rect 13044 8984 13050 8996
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 16022 9024 16028 9036
rect 15703 8996 16028 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 13081 8959 13139 8965
rect 10284 8928 10329 8956
rect 10284 8916 10290 8928
rect 13081 8925 13093 8959
rect 13127 8956 13139 8959
rect 13446 8956 13452 8968
rect 13127 8928 13452 8956
rect 13127 8925 13139 8928
rect 13081 8919 13139 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 15378 8956 15384 8968
rect 15151 8928 15384 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 15378 8916 15384 8928
rect 15436 8956 15442 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15436 8928 15761 8956
rect 15436 8916 15442 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15749 8919 15807 8925
rect 10318 8888 10324 8900
rect 8067 8860 10324 8888
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 11609 8891 11667 8897
rect 11609 8857 11621 8891
rect 11655 8888 11667 8891
rect 11974 8888 11980 8900
rect 11655 8860 11980 8888
rect 11655 8857 11667 8860
rect 11609 8851 11667 8857
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12437 8891 12495 8897
rect 12437 8857 12449 8891
rect 12483 8888 12495 8891
rect 14274 8888 14280 8900
rect 12483 8860 14280 8888
rect 12483 8857 12495 8860
rect 12437 8851 12495 8857
rect 14274 8848 14280 8860
rect 14332 8848 14338 8900
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5442 8820 5448 8832
rect 5215 8792 5448 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 7190 8820 7196 8832
rect 7151 8792 7196 8820
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7466 8820 7472 8832
rect 7427 8792 7472 8820
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10226 8820 10232 8832
rect 10008 8792 10232 8820
rect 10008 8780 10014 8792
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 11238 8820 11244 8832
rect 11199 8792 11244 8820
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11848 8792 11897 8820
rect 11848 8780 11854 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 14642 8820 14648 8832
rect 14603 8792 14648 8820
rect 11885 8783 11943 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15764 8820 15792 8919
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 15838 8820 15844 8832
rect 15764 8792 15844 8820
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17221 8823 17279 8829
rect 17221 8789 17233 8823
rect 17267 8820 17279 8823
rect 17494 8820 17500 8832
rect 17267 8792 17500 8820
rect 17267 8789 17279 8792
rect 17221 8783 17279 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17589 8823 17647 8829
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 17862 8820 17868 8832
rect 17635 8792 17868 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 1854 8616 1860 8628
rect 1811 8588 1860 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 4890 8616 4896 8628
rect 3651 8588 4896 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6236 8588 6561 8616
rect 6236 8576 6242 8588
rect 6549 8585 6561 8588
rect 6595 8616 6607 8619
rect 8018 8616 8024 8628
rect 6595 8588 7328 8616
rect 7979 8588 8024 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 4062 8548 4068 8560
rect 4023 8520 4068 8548
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1544 8452 1869 8480
rect 1544 8440 1550 8452
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 4614 8480 4620 8492
rect 4575 8452 4620 8480
rect 1857 8443 1915 8449
rect 4614 8440 4620 8452
rect 4672 8480 4678 8492
rect 7300 8489 7328 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 9030 8616 9036 8628
rect 8619 8588 9036 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 11790 8616 11796 8628
rect 10827 8588 11796 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12894 8576 12900 8628
rect 12952 8616 12958 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 12952 8588 13553 8616
rect 12952 8576 12958 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8616 14151 8619
rect 14550 8616 14556 8628
rect 14139 8588 14556 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16390 8616 16396 8628
rect 16347 8588 16396 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 10597 8551 10655 8557
rect 10597 8548 10609 8551
rect 9364 8520 10609 8548
rect 9364 8508 9370 8520
rect 10597 8517 10609 8520
rect 10643 8517 10655 8551
rect 10597 8511 10655 8517
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 4672 8452 5457 8480
rect 4672 8440 4678 8452
rect 5445 8449 5457 8452
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7379 8452 7472 8480
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8480 7530 8492
rect 8018 8480 8024 8492
rect 7524 8452 8024 8480
rect 7524 8440 7530 8452
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2113 8415 2171 8421
rect 2113 8412 2125 8415
rect 2004 8384 2125 8412
rect 2004 8372 2010 8384
rect 2113 8381 2125 8384
rect 2159 8381 2171 8415
rect 2113 8375 2171 8381
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4430 8412 4436 8424
rect 4019 8384 4292 8412
rect 4391 8384 4436 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 4062 8344 4068 8356
rect 2832 8316 4068 8344
rect 2832 8304 2838 8316
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4264 8344 4292 8384
rect 4430 8372 4436 8384
rect 4488 8412 4494 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4488 8384 5089 8412
rect 4488 8372 4494 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 8386 8412 8392 8424
rect 8347 8384 8392 8412
rect 5077 8375 5135 8381
rect 8386 8372 8392 8384
rect 8444 8412 8450 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8444 8384 8953 8412
rect 8444 8372 8450 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8381 10379 8415
rect 10612 8412 10640 8511
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 11296 8452 11345 8480
rect 11296 8440 11302 8452
rect 11333 8449 11345 8452
rect 11379 8480 11391 8483
rect 11698 8480 11704 8492
rect 11379 8452 11704 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11808 8480 11836 8576
rect 12529 8551 12587 8557
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 13262 8548 13268 8560
rect 12575 8520 13268 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 13262 8508 13268 8520
rect 13320 8508 13326 8560
rect 15378 8508 15384 8560
rect 15436 8548 15442 8560
rect 15565 8551 15623 8557
rect 15565 8548 15577 8551
rect 15436 8520 15577 8548
rect 15436 8508 15442 8520
rect 15565 8517 15577 8520
rect 15611 8517 15623 8551
rect 15565 8511 15623 8517
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16022 8548 16028 8560
rect 15979 8520 16028 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 11808 8452 13001 8480
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 14182 8480 14188 8492
rect 14143 8452 14188 8480
rect 13173 8443 13231 8449
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10612 8384 11161 8412
rect 10321 8375 10379 8381
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8412 11943 8415
rect 11931 8384 13032 8412
rect 11931 8381 11943 8384
rect 11885 8375 11943 8381
rect 4798 8344 4804 8356
rect 4264 8316 4804 8344
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5629 8347 5687 8353
rect 5500 8316 5580 8344
rect 5500 8304 5506 8316
rect 3234 8276 3240 8288
rect 3195 8248 3240 8276
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 4304 8248 4537 8276
rect 4304 8236 4310 8248
rect 4525 8245 4537 8248
rect 4571 8245 4583 8279
rect 5552 8276 5580 8316
rect 5629 8313 5641 8347
rect 5675 8344 5687 8347
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5675 8316 6285 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 6273 8313 6285 8316
rect 6319 8344 6331 8347
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6319 8316 7205 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 9674 8344 9680 8356
rect 9587 8316 9680 8344
rect 7193 8307 7251 8313
rect 6546 8276 6552 8288
rect 5552 8248 6552 8276
rect 4525 8239 4583 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6822 8276 6828 8288
rect 6783 8248 6828 8276
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 9033 8279 9091 8285
rect 9033 8245 9045 8279
rect 9079 8276 9091 8279
rect 9122 8276 9128 8288
rect 9079 8248 9128 8276
rect 9079 8245 9091 8248
rect 9033 8239 9091 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9600 8276 9628 8316
rect 9674 8304 9680 8316
rect 9732 8344 9738 8356
rect 9732 8316 10180 8344
rect 9732 8304 9738 8316
rect 10152 8285 10180 8316
rect 9548 8248 9628 8276
rect 10137 8279 10195 8285
rect 9548 8236 9554 8248
rect 10137 8245 10149 8279
rect 10183 8245 10195 8279
rect 10336 8276 10364 8375
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11241 8347 11299 8353
rect 11241 8344 11253 8347
rect 11020 8316 11253 8344
rect 11020 8304 11026 8316
rect 11241 8313 11253 8316
rect 11287 8313 11299 8347
rect 11241 8307 11299 8313
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 12158 8344 12164 8356
rect 11388 8316 12164 8344
rect 11388 8304 11394 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 13004 8344 13032 8384
rect 13188 8344 13216 8443
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16448 8384 16865 8412
rect 16448 8372 16454 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 17494 8412 17500 8424
rect 17455 8384 17500 8412
rect 16853 8375 16911 8381
rect 17494 8372 17500 8384
rect 17552 8372 17558 8424
rect 13538 8344 13544 8356
rect 13004 8316 13544 8344
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 14452 8347 14510 8353
rect 14452 8313 14464 8347
rect 14498 8344 14510 8347
rect 14550 8344 14556 8356
rect 14498 8316 14556 8344
rect 14498 8313 14510 8316
rect 14452 8307 14510 8313
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 16482 8344 16488 8356
rect 15344 8316 16488 8344
rect 15344 8304 15350 8316
rect 16482 8304 16488 8316
rect 16540 8344 16546 8356
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 16540 8316 16773 8344
rect 16540 8304 16546 8316
rect 16761 8313 16773 8316
rect 16807 8313 16819 8347
rect 17862 8344 17868 8356
rect 17823 8316 17868 8344
rect 16761 8307 16819 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 12066 8276 12072 8288
rect 10336 8248 12072 8276
rect 10137 8239 10195 8245
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 16390 8276 16396 8288
rect 16351 8248 16396 8276
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 2682 8072 2688 8084
rect 2639 8044 2688 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 3200 8044 3249 8072
rect 3200 8032 3206 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 3237 8035 3295 8041
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4614 8072 4620 8084
rect 3927 8044 4620 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8041 4951 8075
rect 5534 8072 5540 8084
rect 5447 8044 5540 8072
rect 4893 8035 4951 8041
rect 2866 7964 2872 8016
rect 2924 8004 2930 8016
rect 4908 8004 4936 8035
rect 5534 8032 5540 8044
rect 5592 8072 5598 8084
rect 6822 8072 6828 8084
rect 5592 8044 6828 8072
rect 5592 8032 5598 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7374 8072 7380 8084
rect 7239 8044 7380 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 4982 8004 4988 8016
rect 2924 7976 4988 8004
rect 2924 7964 2930 7976
rect 4982 7964 4988 7976
rect 5040 8004 5046 8016
rect 5040 7976 6316 8004
rect 5040 7964 5046 7976
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 6178 7936 6184 7948
rect 5123 7908 6184 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6288 7936 6316 7976
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 7208 8004 7236 8035
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7984 8044 8033 8072
rect 7984 8032 7990 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 8570 8072 8576 8084
rect 8527 8044 8576 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9950 8072 9956 8084
rect 9911 8044 9956 8072
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10229 8075 10287 8081
rect 10229 8072 10241 8075
rect 10192 8044 10241 8072
rect 10192 8032 10198 8044
rect 10229 8041 10241 8044
rect 10275 8041 10287 8075
rect 10229 8035 10287 8041
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 12894 8072 12900 8084
rect 12216 8044 12900 8072
rect 12216 8032 12222 8044
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13630 8072 13636 8084
rect 13403 8044 13636 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 13817 8075 13875 8081
rect 13817 8072 13829 8075
rect 13780 8044 13829 8072
rect 13780 8032 13786 8044
rect 13817 8041 13829 8044
rect 13863 8041 13875 8075
rect 13817 8035 13875 8041
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14366 8072 14372 8084
rect 13964 8044 14372 8072
rect 13964 8032 13970 8044
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 15286 8072 15292 8084
rect 15247 8044 15292 8072
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 15988 8044 16221 8072
rect 15988 8032 15994 8044
rect 16209 8041 16221 8044
rect 16255 8072 16267 8075
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16255 8044 17693 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 8754 8004 8760 8016
rect 6604 7976 7236 8004
rect 7291 7976 8760 8004
rect 6604 7964 6610 7976
rect 7291 7936 7319 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 16568 8007 16626 8013
rect 16568 7973 16580 8007
rect 16614 8004 16626 8007
rect 16666 8004 16672 8016
rect 16614 7976 16672 8004
rect 16614 7973 16626 7976
rect 16568 7967 16626 7973
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 18966 8004 18972 8016
rect 16776 7976 18972 8004
rect 8570 7936 8576 7948
rect 6288 7908 7319 7936
rect 8531 7908 8576 7936
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 10686 7936 10692 7948
rect 9539 7908 10692 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 10962 7945 10968 7948
rect 10945 7939 10968 7945
rect 10945 7936 10957 7939
rect 10836 7908 10957 7936
rect 10836 7896 10842 7908
rect 10945 7905 10957 7908
rect 11020 7936 11026 7948
rect 11020 7908 11093 7936
rect 10945 7899 10968 7905
rect 10962 7896 10968 7899
rect 11020 7896 11026 7908
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 13354 7936 13360 7948
rect 12492 7908 13360 7936
rect 12492 7896 12498 7908
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 13725 7939 13783 7945
rect 13725 7936 13737 7939
rect 13688 7908 13737 7936
rect 13688 7896 13694 7908
rect 13725 7905 13737 7908
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 16776 7936 16804 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 18874 7936 18880 7948
rect 13872 7908 16804 7936
rect 18835 7908 18880 7936
rect 13872 7896 13878 7908
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3142 7868 3148 7880
rect 2915 7840 3148 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 5224 7840 5641 7868
rect 5224 7828 5230 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7800 4859 7803
rect 5736 7800 5764 7831
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7248 7840 7297 7868
rect 7248 7828 7254 7840
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 13446 7868 13452 7880
rect 12575 7840 13452 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 13446 7828 13452 7840
rect 13504 7868 13510 7880
rect 13909 7871 13967 7877
rect 13909 7868 13921 7871
rect 13504 7840 13921 7868
rect 13504 7828 13510 7840
rect 13909 7837 13921 7840
rect 13955 7837 13967 7871
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 13909 7831 13967 7837
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 6086 7800 6092 7812
rect 4847 7772 6092 7800
rect 4847 7769 4859 7772
rect 4801 7763 4859 7769
rect 6086 7760 6092 7772
rect 6144 7760 6150 7812
rect 6641 7803 6699 7809
rect 6641 7769 6653 7803
rect 6687 7800 6699 7803
rect 7374 7800 7380 7812
rect 6687 7772 7380 7800
rect 6687 7769 6699 7772
rect 6641 7763 6699 7769
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 11974 7760 11980 7812
rect 12032 7800 12038 7812
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 12032 7772 14565 7800
rect 12032 7760 12038 7772
rect 14553 7769 14565 7772
rect 14599 7800 14611 7803
rect 14642 7800 14648 7812
rect 14599 7772 14648 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 16316 7800 16344 7831
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 19061 7871 19119 7877
rect 19061 7868 19073 7871
rect 17828 7840 19073 7868
rect 17828 7828 17834 7840
rect 19061 7837 19073 7840
rect 19107 7837 19119 7871
rect 19061 7831 19119 7837
rect 14844 7772 16344 7800
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5169 7735 5227 7741
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5442 7732 5448 7744
rect 5215 7704 5448 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6454 7732 6460 7744
rect 6319 7704 6460 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6730 7732 6736 7744
rect 6691 7704 6736 7732
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 9122 7732 9128 7744
rect 9083 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 12066 7732 12072 7744
rect 12027 7704 12072 7732
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 13446 7732 13452 7744
rect 13219 7704 13452 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14090 7732 14096 7744
rect 13964 7704 14096 7732
rect 13964 7692 13970 7704
rect 14090 7692 14096 7704
rect 14148 7692 14154 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14844 7741 14872 7772
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14240 7704 14841 7732
rect 14240 7692 14246 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 18012 7704 18061 7732
rect 18012 7692 18018 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18506 7732 18512 7744
rect 18467 7704 18512 7732
rect 18049 7695 18107 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6546 7528 6552 7540
rect 6319 7500 6552 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 2501 7463 2559 7469
rect 2501 7460 2513 7463
rect 1820 7432 2513 7460
rect 1820 7420 1826 7432
rect 2501 7429 2513 7432
rect 2547 7429 2559 7463
rect 2501 7423 2559 7429
rect 4709 7463 4767 7469
rect 4709 7429 4721 7463
rect 4755 7460 4767 7463
rect 5350 7460 5356 7472
rect 4755 7432 5356 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2516 7392 2544 7423
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 6288 7460 6316 7491
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7156 7500 7849 7528
rect 7156 7488 7162 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 10778 7528 10784 7540
rect 10739 7500 10784 7528
rect 7837 7491 7895 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 12250 7528 12256 7540
rect 11664 7500 12256 7528
rect 11664 7488 11670 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13354 7528 13360 7540
rect 13035 7500 13360 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16448 7500 16957 7528
rect 16448 7488 16454 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 16945 7491 17003 7497
rect 17402 7488 17408 7500
rect 17460 7528 17466 7540
rect 18598 7528 18604 7540
rect 17460 7500 18604 7528
rect 17460 7488 17466 7500
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 19024 7500 19073 7528
rect 19024 7488 19030 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19061 7491 19119 7497
rect 5684 7432 6316 7460
rect 5684 7420 5690 7432
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 10744 7432 11805 7460
rect 10744 7420 10750 7432
rect 11793 7429 11805 7432
rect 11839 7429 11851 7463
rect 15470 7460 15476 7472
rect 15383 7432 15476 7460
rect 11793 7423 11851 7429
rect 15470 7420 15476 7432
rect 15528 7460 15534 7472
rect 15528 7432 16160 7460
rect 15528 7420 15534 7432
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2516 7364 3525 7392
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 3786 7392 3792 7404
rect 3651 7364 3792 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1728 7296 1869 7324
rect 1728 7284 1734 7296
rect 1857 7293 1869 7296
rect 1903 7324 1915 7327
rect 2774 7324 2780 7336
rect 1903 7296 2780 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3007 7296 3433 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3421 7293 3433 7296
rect 3467 7324 3479 7327
rect 3694 7324 3700 7336
rect 3467 7296 3700 7324
rect 3467 7293 3479 7296
rect 3421 7287 3479 7293
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 5368 7324 5396 7420
rect 16132 7404 16160 7432
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5994 7392 6000 7404
rect 5859 7364 6000 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 8570 7352 8576 7404
rect 8628 7392 8634 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8628 7364 8677 7392
rect 8628 7352 8634 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 8665 7355 8723 7361
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5368 7296 5549 7324
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 7193 7327 7251 7333
rect 7193 7293 7205 7327
rect 7239 7324 7251 7327
rect 7282 7324 7288 7336
rect 7239 7296 7288 7324
rect 7239 7293 7251 7296
rect 7193 7287 7251 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8680 7324 8708 7355
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12176 7364 13093 7392
rect 9490 7324 9496 7336
rect 8680 7296 9496 7324
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10413 7327 10471 7333
rect 10413 7324 10425 7327
rect 9732 7296 10425 7324
rect 9732 7284 9738 7296
rect 10413 7293 10425 7296
rect 10459 7324 10471 7327
rect 11974 7324 11980 7336
rect 10459 7296 11980 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 1995 7228 3096 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 3068 7200 3096 7228
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 4985 7259 5043 7265
rect 4985 7256 4997 7259
rect 3936 7228 4997 7256
rect 3936 7216 3942 7228
rect 4985 7225 4997 7228
rect 5031 7256 5043 7259
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 5031 7228 5641 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 5629 7225 5641 7228
rect 5675 7256 5687 7259
rect 6270 7256 6276 7268
rect 5675 7228 6276 7256
rect 5675 7225 5687 7228
rect 5629 7219 5687 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 8938 7265 8944 7268
rect 8573 7259 8631 7265
rect 6564 7228 7328 7256
rect 6564 7200 6592 7228
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4890 7188 4896 7200
rect 4387 7160 4896 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 6914 7188 6920 7200
rect 6871 7160 6920 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7300 7197 7328 7228
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8932 7256 8944 7265
rect 8619 7228 8944 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 8932 7219 8944 7228
rect 8938 7216 8944 7219
rect 8996 7216 9002 7268
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 11330 7256 11336 7268
rect 10008 7228 11336 7256
rect 10008 7216 10014 7228
rect 11330 7216 11336 7228
rect 11388 7216 11394 7268
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 12176 7265 12204 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15746 7392 15752 7404
rect 15151 7364 15752 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15746 7352 15752 7364
rect 15804 7392 15810 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15804 7364 16037 7392
rect 15804 7352 15810 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 16172 7364 16265 7392
rect 16172 7352 16178 7364
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18012 7364 18613 7392
rect 18012 7352 18018 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7324 15991 7327
rect 16390 7324 16396 7336
rect 15979 7296 16396 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 17770 7324 17776 7336
rect 17731 7296 17776 7324
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18230 7324 18236 7336
rect 18104 7296 18236 7324
rect 18104 7284 18110 7296
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7324 18570 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18564 7296 19441 7324
rect 18564 7284 18570 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 12124 7228 12173 7256
rect 12124 7216 12130 7228
rect 12161 7225 12173 7228
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 13348 7259 13406 7265
rect 13348 7225 13360 7259
rect 13394 7256 13406 7259
rect 13446 7256 13452 7268
rect 13394 7228 13452 7256
rect 13394 7225 13406 7228
rect 13348 7219 13406 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7157 7343 7191
rect 7285 7151 7343 7157
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10134 7188 10140 7200
rect 10091 7160 10140 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 11149 7191 11207 7197
rect 11149 7157 11161 7191
rect 11195 7188 11207 7191
rect 11238 7188 11244 7200
rect 11195 7160 11244 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15565 7191 15623 7197
rect 15565 7188 15577 7191
rect 15252 7160 15577 7188
rect 15252 7148 15258 7160
rect 15565 7157 15577 7160
rect 15611 7157 15623 7191
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 15565 7151 15623 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 18046 7188 18052 7200
rect 18007 7160 18052 7188
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18598 7188 18604 7200
rect 18555 7160 18604 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3605 6987 3663 6993
rect 3605 6984 3617 6987
rect 3108 6956 3617 6984
rect 3108 6944 3114 6956
rect 3605 6953 3617 6956
rect 3651 6953 3663 6987
rect 3605 6947 3663 6953
rect 4709 6987 4767 6993
rect 4709 6953 4721 6987
rect 4755 6984 4767 6987
rect 5166 6984 5172 6996
rect 4755 6956 5172 6984
rect 4755 6953 4767 6956
rect 4709 6947 4767 6953
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 6181 6987 6239 6993
rect 6181 6984 6193 6987
rect 6144 6956 6193 6984
rect 6144 6944 6150 6956
rect 6181 6953 6193 6956
rect 6227 6953 6239 6987
rect 6181 6947 6239 6953
rect 6549 6987 6607 6993
rect 6549 6953 6561 6987
rect 6595 6984 6607 6987
rect 7190 6984 7196 6996
rect 6595 6956 7196 6984
rect 6595 6953 6607 6956
rect 6549 6947 6607 6953
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 8754 6984 8760 6996
rect 8715 6956 8760 6984
rect 8754 6944 8760 6956
rect 8812 6944 8818 6996
rect 13449 6987 13507 6993
rect 13449 6953 13461 6987
rect 13495 6984 13507 6987
rect 13538 6984 13544 6996
rect 13495 6956 13544 6984
rect 13495 6953 13507 6956
rect 13449 6947 13507 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 13722 6984 13728 6996
rect 13683 6956 13728 6984
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 18785 6987 18843 6993
rect 18785 6953 18797 6987
rect 18831 6984 18843 6987
rect 18874 6984 18880 6996
rect 18831 6956 18880 6984
rect 18831 6953 18843 6956
rect 18785 6947 18843 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 1848 6919 1906 6925
rect 1848 6885 1860 6919
rect 1894 6916 1906 6919
rect 2038 6916 2044 6928
rect 1894 6888 2044 6916
rect 1894 6885 1906 6888
rect 1848 6879 1906 6885
rect 2038 6876 2044 6888
rect 2096 6876 2102 6928
rect 3329 6919 3387 6925
rect 3329 6885 3341 6919
rect 3375 6916 3387 6919
rect 3786 6916 3792 6928
rect 3375 6888 3792 6916
rect 3375 6885 3387 6888
rect 3329 6879 3387 6885
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 4982 6916 4988 6928
rect 4816 6888 4988 6916
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 1452 6820 1593 6848
rect 1452 6808 1458 6820
rect 1581 6817 1593 6820
rect 1627 6848 1639 6851
rect 2866 6848 2872 6860
rect 1627 6820 2872 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4816 6857 4844 6888
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 7276 6919 7334 6925
rect 7276 6885 7288 6919
rect 7322 6916 7334 6919
rect 7374 6916 7380 6928
rect 7322 6888 7380 6916
rect 7322 6885 7334 6888
rect 7276 6879 7334 6885
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 12526 6876 12532 6928
rect 12584 6876 12590 6928
rect 16114 6876 16120 6928
rect 16172 6925 16178 6928
rect 16172 6919 16236 6925
rect 16172 6885 16190 6919
rect 16224 6885 16236 6919
rect 16172 6879 16236 6885
rect 16172 6876 16178 6879
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5068 6851 5126 6857
rect 5068 6848 5080 6851
rect 4948 6820 5080 6848
rect 4948 6808 4954 6820
rect 5068 6817 5080 6820
rect 5114 6848 5126 6851
rect 5994 6848 6000 6860
rect 5114 6820 6000 6848
rect 5114 6817 5126 6820
rect 5068 6811 5126 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 8570 6848 8576 6860
rect 7055 6820 8576 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9933 6851 9991 6857
rect 9933 6848 9945 6851
rect 9824 6820 9945 6848
rect 9824 6808 9830 6820
rect 9933 6817 9945 6820
rect 9979 6817 9991 6851
rect 9933 6811 9991 6817
rect 12336 6851 12394 6857
rect 12336 6817 12348 6851
rect 12382 6848 12394 6851
rect 12544 6848 12572 6876
rect 17589 6851 17647 6857
rect 17589 6848 17601 6851
rect 12382 6820 12572 6848
rect 15948 6820 17601 6848
rect 12382 6817 12394 6820
rect 12336 6811 12394 6817
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9416 6752 9689 6780
rect 5902 6672 5908 6724
rect 5960 6712 5966 6724
rect 6270 6712 6276 6724
rect 5960 6684 6276 6712
rect 5960 6672 5966 6684
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2372 6616 2973 6644
rect 2372 6604 2378 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 5534 6644 5540 6656
rect 4387 6616 5540 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7282 6644 7288 6656
rect 6963 6616 7288 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 8076 6616 8401 6644
rect 8076 6604 8082 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 8389 6607 8447 6613
rect 9030 6604 9036 6616
rect 9088 6644 9094 6656
rect 9416 6653 9444 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 12066 6780 12072 6792
rect 9677 6743 9735 6749
rect 11164 6752 12072 6780
rect 11054 6712 11060 6724
rect 11015 6684 11060 6712
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9088 6616 9413 6644
rect 9088 6604 9094 6616
rect 9401 6613 9413 6616
rect 9447 6644 9459 6647
rect 11164 6644 11192 6752
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14734 6780 14740 6792
rect 14516 6752 14740 6780
rect 14516 6740 14522 6752
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15948 6789 15976 6820
rect 17589 6817 17601 6820
rect 17635 6848 17647 6851
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17635 6820 17969 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 19426 6848 19432 6860
rect 18187 6820 19432 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15344 6752 15945 6780
rect 15344 6740 15350 6752
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 17972 6780 18000 6811
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 19061 6783 19119 6789
rect 19061 6780 19073 6783
rect 17972 6752 19073 6780
rect 15933 6743 15991 6749
rect 19061 6749 19073 6752
rect 19107 6780 19119 6783
rect 19150 6780 19156 6792
rect 19107 6752 19156 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 15194 6712 15200 6724
rect 14752 6684 15200 6712
rect 14752 6656 14780 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 19518 6712 19524 6724
rect 19431 6684 19524 6712
rect 19518 6672 19524 6684
rect 19576 6712 19582 6724
rect 20438 6712 20444 6724
rect 19576 6684 20444 6712
rect 19576 6672 19582 6684
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 9447 6616 11192 6644
rect 11425 6647 11483 6653
rect 9447 6613 9459 6616
rect 9401 6607 9459 6613
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11514 6644 11520 6656
rect 11471 6616 11520 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11664 6616 11713 6644
rect 11664 6604 11670 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 13630 6644 13636 6656
rect 12032 6616 13636 6644
rect 12032 6604 12038 6616
rect 13630 6604 13636 6616
rect 13688 6644 13694 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13688 6616 14105 6644
rect 13688 6604 13694 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 14093 6607 14151 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15105 6647 15163 6653
rect 15105 6613 15117 6647
rect 15151 6644 15163 6647
rect 15562 6644 15568 6656
rect 15151 6616 15568 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15841 6647 15899 6653
rect 15841 6613 15853 6647
rect 15887 6644 15899 6647
rect 16298 6644 16304 6656
rect 15887 6616 16304 6644
rect 15887 6613 15899 6616
rect 15841 6607 15899 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 17313 6647 17371 6653
rect 17313 6644 17325 6647
rect 16724 6616 17325 6644
rect 16724 6604 16730 6616
rect 17313 6613 17325 6616
rect 17359 6613 17371 6647
rect 17313 6607 17371 6613
rect 18325 6647 18383 6653
rect 18325 6613 18337 6647
rect 18371 6644 18383 6647
rect 18506 6644 18512 6656
rect 18371 6616 18512 6644
rect 18371 6613 18383 6616
rect 18325 6607 18383 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 19889 6647 19947 6653
rect 19889 6613 19901 6647
rect 19935 6644 19947 6647
rect 20254 6644 20260 6656
rect 19935 6616 20260 6644
rect 19935 6613 19947 6616
rect 19889 6607 19947 6613
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 3970 6440 3976 6452
rect 3651 6412 3976 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4890 6440 4896 6452
rect 4387 6412 4896 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6144 6412 6561 6440
rect 6144 6400 6150 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 5169 6375 5227 6381
rect 5169 6341 5181 6375
rect 5215 6372 5227 6375
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 5215 6344 6193 6372
rect 5215 6341 5227 6344
rect 5169 6335 5227 6341
rect 6181 6341 6193 6344
rect 6227 6341 6239 6375
rect 6181 6335 6239 6341
rect 1394 6264 1400 6316
rect 1452 6304 1458 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 1452 6276 1501 6304
rect 1452 6264 1458 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 2832 6276 3709 6304
rect 2832 6264 2838 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 5994 6264 6000 6276
rect 6052 6304 6058 6316
rect 6052 6276 6132 6304
rect 6052 6264 6058 6276
rect 1762 6177 1768 6180
rect 1756 6168 1768 6177
rect 1723 6140 1768 6168
rect 1756 6131 1768 6140
rect 1762 6128 1768 6131
rect 1820 6128 1826 6180
rect 5537 6171 5595 6177
rect 5537 6168 5549 6171
rect 4632 6140 5549 6168
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2866 6100 2872 6112
rect 2096 6072 2872 6100
rect 2096 6060 2102 6072
rect 2866 6060 2872 6072
rect 2924 6100 2930 6112
rect 3145 6103 3203 6109
rect 3145 6100 3157 6103
rect 2924 6072 3157 6100
rect 2924 6060 2930 6072
rect 3145 6069 3157 6072
rect 3191 6069 3203 6103
rect 3145 6063 3203 6069
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4632 6109 4660 6140
rect 5537 6137 5549 6140
rect 5583 6137 5595 6171
rect 6104 6168 6132 6276
rect 6196 6236 6224 6335
rect 6564 6304 6592 6403
rect 7374 6400 7380 6452
rect 7432 6440 7438 6452
rect 7650 6440 7656 6452
rect 7432 6412 7656 6440
rect 7432 6400 7438 6412
rect 7650 6400 7656 6412
rect 7708 6440 7714 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7708 6412 7849 6440
rect 7708 6400 7714 6412
rect 7837 6409 7849 6412
rect 7883 6440 7895 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 7883 6412 10057 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 11698 6400 11704 6452
rect 11756 6440 11762 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 11756 6412 12081 6440
rect 11756 6400 11762 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 12069 6403 12127 6409
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6440 15163 6443
rect 15470 6440 15476 6452
rect 15151 6412 15476 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 15470 6400 15476 6412
rect 15528 6440 15534 6452
rect 16758 6440 16764 6452
rect 15528 6412 16764 6440
rect 15528 6400 15534 6412
rect 16758 6400 16764 6412
rect 16816 6440 16822 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16816 6412 16957 6440
rect 16816 6400 16822 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 16945 6403 17003 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10321 6375 10379 6381
rect 10321 6372 10333 6375
rect 9824 6344 10333 6372
rect 9824 6332 9830 6344
rect 10321 6341 10333 6344
rect 10367 6341 10379 6375
rect 10321 6335 10379 6341
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 6564 6276 7389 6304
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 17788 6304 17816 6400
rect 18598 6304 18604 6316
rect 15519 6276 15700 6304
rect 17788 6276 18604 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6196 6208 7205 6236
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 11241 6239 11299 6245
rect 11241 6236 11253 6239
rect 7193 6199 7251 6205
rect 11164 6208 11253 6236
rect 8018 6168 8024 6180
rect 6104 6140 8024 6168
rect 5537 6131 5595 6137
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8573 6171 8631 6177
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 8932 6171 8990 6177
rect 8932 6168 8944 6171
rect 8619 6140 8944 6168
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 8932 6137 8944 6140
rect 8978 6168 8990 6171
rect 10134 6168 10140 6180
rect 8978 6140 10140 6168
rect 8978 6137 8990 6140
rect 8932 6131 8990 6137
rect 10134 6128 10140 6140
rect 10192 6128 10198 6180
rect 11164 6112 11192 6208
rect 11241 6205 11253 6208
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 12066 6196 12072 6248
rect 12124 6236 12130 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12124 6208 12725 6236
rect 12124 6196 12130 6208
rect 12713 6205 12725 6208
rect 12759 6236 12771 6239
rect 12759 6208 13216 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 12980 6171 13038 6177
rect 12980 6137 12992 6171
rect 13026 6137 13038 6171
rect 13188 6168 13216 6208
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 13320 6208 14381 6236
rect 13320 6196 13326 6208
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6205 15623 6239
rect 15672 6236 15700 6276
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 15832 6239 15890 6245
rect 15832 6236 15844 6239
rect 15672 6208 15844 6236
rect 15565 6199 15623 6205
rect 15832 6205 15844 6208
rect 15878 6236 15890 6239
rect 16206 6236 16212 6248
rect 15878 6208 16212 6236
rect 15878 6205 15890 6208
rect 15832 6199 15890 6205
rect 14182 6168 14188 6180
rect 13188 6140 14188 6168
rect 12980 6131 13038 6137
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4212 6072 4629 6100
rect 4212 6060 4218 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4617 6063 4675 6069
rect 4982 6060 4988 6072
rect 5040 6100 5046 6112
rect 5626 6100 5632 6112
rect 5040 6072 5632 6100
rect 5040 6060 5046 6072
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 7374 6100 7380 6112
rect 7331 6072 7380 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 10962 6100 10968 6112
rect 10827 6072 10968 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11422 6100 11428 6112
rect 11383 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 12995 6100 13023 6131
rect 14182 6128 14188 6140
rect 14240 6168 14246 6180
rect 15286 6168 15292 6180
rect 14240 6140 15292 6168
rect 14240 6128 14246 6140
rect 15286 6128 15292 6140
rect 15344 6168 15350 6180
rect 15580 6168 15608 6199
rect 16040 6180 16068 6208
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17920 6208 18429 6236
rect 17920 6196 17926 6208
rect 18417 6205 18429 6208
rect 18463 6236 18475 6239
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18463 6208 19073 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 15344 6140 15608 6168
rect 15344 6128 15350 6140
rect 16022 6128 16028 6180
rect 16080 6128 16086 6180
rect 17497 6171 17555 6177
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 17954 6168 17960 6180
rect 17543 6140 17960 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 17954 6128 17960 6140
rect 18012 6168 18018 6180
rect 18509 6171 18567 6177
rect 18509 6168 18521 6171
rect 18012 6140 18521 6168
rect 18012 6128 18018 6140
rect 18509 6137 18521 6140
rect 18555 6137 18567 6171
rect 18509 6131 18567 6137
rect 19150 6128 19156 6180
rect 19208 6168 19214 6180
rect 19889 6171 19947 6177
rect 19889 6168 19901 6171
rect 19208 6140 19901 6168
rect 19208 6128 19214 6140
rect 19889 6137 19901 6140
rect 19935 6168 19947 6171
rect 20622 6168 20628 6180
rect 19935 6140 20628 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 13538 6100 13544 6112
rect 12860 6072 13544 6100
rect 12860 6060 12866 6072
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15930 6100 15936 6112
rect 15528 6072 15936 6100
rect 15528 6060 15534 6072
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 20254 6100 20260 6112
rect 20167 6072 20260 6100
rect 20254 6060 20260 6072
rect 20312 6100 20318 6112
rect 20714 6100 20720 6112
rect 20312 6072 20720 6100
rect 20312 6060 20318 6072
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2038 5896 2044 5908
rect 1999 5868 2044 5896
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 3697 5899 3755 5905
rect 3697 5865 3709 5899
rect 3743 5896 3755 5899
rect 4062 5896 4068 5908
rect 3743 5868 4068 5896
rect 3743 5865 3755 5868
rect 3697 5859 3755 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4890 5896 4896 5908
rect 4851 5868 4896 5896
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7374 5896 7380 5908
rect 6963 5868 7380 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 9030 5896 9036 5908
rect 8619 5868 9036 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10045 5899 10103 5905
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 10686 5896 10692 5908
rect 10091 5868 10692 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3844 5800 4261 5828
rect 3844 5788 3850 5800
rect 4249 5797 4261 5800
rect 4295 5828 4307 5831
rect 4430 5828 4436 5840
rect 4295 5800 4436 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5436 5831 5494 5837
rect 5436 5828 5448 5831
rect 5316 5800 5448 5828
rect 5316 5788 5322 5800
rect 5436 5797 5448 5800
rect 5482 5828 5494 5831
rect 6086 5828 6092 5840
rect 5482 5800 6092 5828
rect 5482 5797 5494 5800
rect 5436 5791 5494 5797
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5828 8999 5831
rect 10060 5828 10088 5859
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11974 5896 11980 5908
rect 11287 5868 11980 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14792 5868 14872 5896
rect 14792 5856 14798 5868
rect 8987 5800 10088 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 11112 5800 11713 5828
rect 11112 5788 11118 5800
rect 11701 5797 11713 5800
rect 11747 5828 11759 5831
rect 11790 5828 11796 5840
rect 11747 5800 11796 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 14844 5828 14872 5868
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15930 5896 15936 5908
rect 15620 5868 15936 5896
rect 15620 5856 15626 5868
rect 15930 5856 15936 5868
rect 15988 5896 15994 5908
rect 16209 5899 16267 5905
rect 16209 5896 16221 5899
rect 15988 5868 16221 5896
rect 15988 5856 15994 5868
rect 16209 5865 16221 5868
rect 16255 5865 16267 5899
rect 16209 5859 16267 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16758 5896 16764 5908
rect 16540 5868 16764 5896
rect 16540 5856 16546 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 19334 5896 19340 5908
rect 17359 5868 19340 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 16117 5831 16175 5837
rect 16117 5828 16129 5831
rect 14844 5800 16129 5828
rect 16117 5797 16129 5800
rect 16163 5797 16175 5831
rect 16117 5791 16175 5797
rect 18230 5788 18236 5840
rect 18288 5828 18294 5840
rect 18325 5831 18383 5837
rect 18325 5828 18337 5831
rect 18288 5800 18337 5828
rect 18288 5788 18294 5800
rect 18325 5797 18337 5800
rect 18371 5797 18383 5831
rect 18690 5828 18696 5840
rect 18651 5800 18696 5828
rect 18325 5791 18383 5797
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 2590 5760 2596 5772
rect 2551 5732 2596 5760
rect 2590 5720 2596 5732
rect 2648 5760 2654 5772
rect 3237 5763 3295 5769
rect 3237 5760 3249 5763
rect 2648 5732 3249 5760
rect 2648 5720 2654 5732
rect 3237 5729 3249 5732
rect 3283 5729 3295 5763
rect 3237 5723 3295 5729
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 5132 5732 5181 5760
rect 5132 5720 5138 5732
rect 5169 5729 5181 5732
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 6972 5732 7757 5760
rect 6972 5720 6978 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11609 5763 11667 5769
rect 11609 5760 11621 5763
rect 11388 5732 11621 5760
rect 11388 5720 11394 5732
rect 11609 5729 11621 5732
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 13412 5732 14289 5760
rect 13412 5720 13418 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14642 5760 14648 5772
rect 14603 5732 14648 5760
rect 14277 5723 14335 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 17678 5760 17684 5772
rect 17639 5732 17684 5760
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 19242 5760 19248 5772
rect 19203 5732 19248 5760
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 7064 5664 7297 5692
rect 7064 5652 7070 5664
rect 7285 5661 7297 5664
rect 7331 5692 7343 5695
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7331 5664 7849 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 7837 5655 7895 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9824 5664 10149 5692
rect 9824 5652 9830 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 11885 5695 11943 5701
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 11885 5661 11897 5695
rect 11931 5692 11943 5695
rect 12342 5692 12348 5704
rect 11931 5664 12348 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13446 5692 13452 5704
rect 12860 5664 13452 5692
rect 12860 5652 12866 5664
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 14090 5692 14096 5704
rect 13504 5664 14096 5692
rect 13504 5652 13510 5664
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 15896 5664 16313 5692
rect 15896 5652 15902 5664
rect 16301 5661 16313 5664
rect 16347 5692 16359 5695
rect 16666 5692 16672 5704
rect 16347 5664 16672 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17368 5664 17785 5692
rect 17368 5652 17374 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5624 1731 5627
rect 1762 5624 1768 5636
rect 1719 5596 1768 5624
rect 1719 5593 1731 5596
rect 1673 5587 1731 5593
rect 1762 5584 1768 5596
rect 1820 5624 1826 5636
rect 3050 5624 3056 5636
rect 1820 5596 3056 5624
rect 1820 5584 1826 5596
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 9674 5624 9680 5636
rect 9635 5596 9680 5624
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 12894 5624 12900 5636
rect 12855 5596 12900 5624
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 13630 5584 13636 5636
rect 13688 5624 13694 5636
rect 14921 5627 14979 5633
rect 14921 5624 14933 5627
rect 13688 5596 14933 5624
rect 13688 5584 13694 5596
rect 14921 5593 14933 5596
rect 14967 5593 14979 5627
rect 14921 5587 14979 5593
rect 15657 5627 15715 5633
rect 15657 5593 15669 5627
rect 15703 5624 15715 5627
rect 16022 5624 16028 5636
rect 15703 5596 16028 5624
rect 15703 5593 15715 5596
rect 15657 5587 15715 5593
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 17129 5627 17187 5633
rect 17129 5624 17141 5627
rect 16632 5596 17141 5624
rect 16632 5584 16638 5596
rect 17129 5593 17141 5596
rect 17175 5593 17187 5627
rect 17129 5587 17187 5593
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 17880 5624 17908 5655
rect 18598 5652 18604 5704
rect 18656 5692 18662 5704
rect 19150 5692 19156 5704
rect 18656 5664 19156 5692
rect 18656 5652 18662 5664
rect 19150 5652 19156 5664
rect 19208 5692 19214 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19208 5664 19441 5692
rect 19208 5652 19214 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 20714 5692 20720 5704
rect 20675 5664 20720 5692
rect 19429 5655 19487 5661
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5692 22799 5695
rect 23474 5692 23480 5704
rect 22787 5664 23480 5692
rect 22787 5661 22799 5664
rect 22741 5655 22799 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 18874 5624 18880 5636
rect 17644 5596 17908 5624
rect 18835 5596 18880 5624
rect 17644 5584 17650 5596
rect 18874 5584 18880 5596
rect 18932 5584 18938 5636
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 6546 5556 6552 5568
rect 6507 5528 6552 5556
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 10781 5559 10839 5565
rect 10781 5556 10793 5559
rect 10744 5528 10793 5556
rect 10744 5516 10750 5528
rect 10781 5525 10793 5528
rect 10827 5525 10839 5559
rect 10781 5519 10839 5525
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12492 5528 12537 5556
rect 12492 5516 12498 5528
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 13909 5559 13967 5565
rect 13909 5556 13921 5559
rect 13872 5528 13921 5556
rect 13872 5516 13878 5528
rect 13909 5525 13921 5528
rect 13955 5525 13967 5559
rect 13909 5519 13967 5525
rect 14182 5516 14188 5568
rect 14240 5556 14246 5568
rect 14461 5559 14519 5565
rect 14461 5556 14473 5559
rect 14240 5528 14473 5556
rect 14240 5516 14246 5528
rect 14461 5525 14473 5528
rect 14507 5525 14519 5559
rect 14461 5519 14519 5525
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 16298 5556 16304 5568
rect 15795 5528 16304 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 19978 5556 19984 5568
rect 19939 5528 19984 5556
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20349 5559 20407 5565
rect 20349 5525 20361 5559
rect 20395 5556 20407 5559
rect 20438 5556 20444 5568
rect 20395 5528 20444 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2590 5352 2596 5364
rect 2455 5324 2596 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 5258 5352 5264 5364
rect 5219 5324 5264 5352
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5408 5324 5641 5352
rect 5408 5312 5414 5324
rect 5629 5321 5641 5324
rect 5675 5352 5687 5355
rect 6730 5352 6736 5364
rect 5675 5324 6736 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 8938 5312 8944 5364
rect 8996 5352 9002 5364
rect 9033 5355 9091 5361
rect 9033 5352 9045 5355
rect 8996 5324 9045 5352
rect 8996 5312 9002 5324
rect 9033 5321 9045 5324
rect 9079 5321 9091 5355
rect 9033 5315 9091 5321
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9582 5352 9588 5364
rect 9263 5324 9588 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 3973 5287 4031 5293
rect 3973 5284 3985 5287
rect 2832 5256 3985 5284
rect 2832 5244 2838 5256
rect 3973 5253 3985 5256
rect 4019 5253 4031 5287
rect 6178 5284 6184 5296
rect 6139 5256 6184 5284
rect 3973 5247 4031 5253
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 9048 5284 9076 5315
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10226 5352 10232 5364
rect 10187 5324 10232 5352
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 11790 5312 11796 5324
rect 11848 5352 11854 5364
rect 12066 5352 12072 5364
rect 11848 5324 12072 5352
rect 11848 5312 11854 5324
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12802 5352 12808 5364
rect 12763 5324 12808 5352
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 12897 5355 12955 5361
rect 12897 5321 12909 5355
rect 12943 5352 12955 5355
rect 13354 5352 13360 5364
rect 12943 5324 13360 5352
rect 12943 5321 12955 5324
rect 12897 5315 12955 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 15930 5312 15936 5364
rect 15988 5352 15994 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15988 5324 16037 5352
rect 15988 5312 15994 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 18012 5324 18061 5352
rect 18012 5312 18018 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 19153 5355 19211 5361
rect 19153 5321 19165 5355
rect 19199 5352 19211 5355
rect 19242 5352 19248 5364
rect 19199 5324 19248 5352
rect 19199 5321 19211 5324
rect 19153 5315 19211 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19392 5324 19809 5352
rect 19392 5312 19398 5324
rect 19797 5321 19809 5324
rect 19843 5321 19855 5355
rect 19797 5315 19855 5321
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 9048 5256 9812 5284
rect 3050 5216 3056 5228
rect 2963 5188 3056 5216
rect 3050 5176 3056 5188
rect 3108 5216 3114 5228
rect 4430 5216 4436 5228
rect 3108 5188 4436 5216
rect 3108 5176 3114 5188
rect 4430 5176 4436 5188
rect 4488 5216 4494 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4488 5188 4537 5216
rect 4488 5176 4494 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9784 5225 9812 5256
rect 13372 5256 14473 5284
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9364 5188 9689 5216
rect 9364 5176 9370 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 10744 5188 11345 5216
rect 10744 5176 10750 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 11333 5179 11391 5185
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 3513 5151 3571 5157
rect 2363 5120 2912 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2884 5089 2912 5120
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 6917 5151 6975 5157
rect 3559 5120 4476 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5080 2927 5083
rect 3970 5080 3976 5092
rect 2915 5052 3976 5080
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 4341 5083 4399 5089
rect 4341 5080 4353 5083
rect 4264 5052 4353 5080
rect 1578 4972 1584 5024
rect 1636 5012 1642 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1636 4984 1869 5012
rect 1636 4972 1642 4984
rect 1857 4981 1869 4984
rect 1903 5012 1915 5015
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 1903 4984 2789 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 3786 5012 3792 5024
rect 3747 4984 3792 5012
rect 2777 4975 2835 4981
rect 3786 4972 3792 4984
rect 3844 5012 3850 5024
rect 4264 5012 4292 5052
rect 4341 5049 4353 5052
rect 4387 5049 4399 5083
rect 4341 5043 4399 5049
rect 4448 5024 4476 5120
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 8570 5148 8576 5160
rect 6963 5120 8576 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 9490 5148 9496 5160
rect 8803 5120 9496 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 9548 5120 9597 5148
rect 9548 5108 9554 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 10652 5120 11253 5148
rect 10652 5108 10658 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 6546 5080 6552 5092
rect 6144 5052 6552 5080
rect 6144 5040 6150 5052
rect 6546 5040 6552 5052
rect 6604 5080 6610 5092
rect 7162 5083 7220 5089
rect 7162 5080 7174 5083
rect 6604 5052 7174 5080
rect 6604 5040 6610 5052
rect 7162 5049 7174 5052
rect 7208 5049 7220 5083
rect 7162 5043 7220 5049
rect 4430 5012 4436 5024
rect 3844 4984 4292 5012
rect 4391 4984 4436 5012
rect 3844 4972 3850 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 9398 5012 9404 5024
rect 8343 4984 9404 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 10962 5012 10968 5024
rect 10827 4984 10968 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11348 5012 11376 5179
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 13372 5225 13400 5256
rect 14461 5253 14473 5256
rect 14507 5253 14519 5287
rect 14461 5247 14519 5253
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 12492 5188 13369 5216
rect 12492 5176 12498 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13357 5179 13415 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 13998 5176 14004 5228
rect 14056 5176 14062 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14976 5188 15117 5216
rect 14976 5176 14982 5188
rect 15105 5185 15117 5188
rect 15151 5216 15163 5219
rect 15378 5216 15384 5228
rect 15151 5188 15384 5216
rect 15151 5185 15163 5188
rect 15105 5179 15163 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16577 5219 16635 5225
rect 16577 5216 16589 5219
rect 16540 5188 16589 5216
rect 16540 5176 16546 5188
rect 16577 5185 16589 5188
rect 16623 5185 16635 5219
rect 16577 5179 16635 5185
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17644 5188 18613 5216
rect 17644 5176 17650 5188
rect 18601 5185 18613 5188
rect 18647 5216 18659 5219
rect 19334 5216 19340 5228
rect 18647 5188 19340 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 19334 5176 19340 5188
rect 19392 5216 19398 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19392 5188 19441 5216
rect 19392 5176 19398 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 13265 5151 13323 5157
rect 13265 5148 13277 5151
rect 11480 5120 13277 5148
rect 11480 5108 11486 5120
rect 13265 5117 13277 5120
rect 13311 5148 13323 5151
rect 13722 5148 13728 5160
rect 13311 5120 13728 5148
rect 13311 5117 13323 5120
rect 13265 5111 13323 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 12526 5012 12532 5024
rect 11348 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12710 4972 12716 5024
rect 12768 5012 12774 5024
rect 13354 5012 13360 5024
rect 12768 4984 13360 5012
rect 12768 4972 12774 4984
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 14016 5021 14044 5176
rect 14090 5108 14096 5160
rect 14148 5148 14154 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14148 5120 14381 5148
rect 14148 5108 14154 5120
rect 14369 5117 14381 5120
rect 14415 5148 14427 5151
rect 14826 5148 14832 5160
rect 14415 5120 14832 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 18230 5108 18236 5160
rect 18288 5148 18294 5160
rect 18417 5151 18475 5157
rect 18417 5148 18429 5151
rect 18288 5120 18429 5148
rect 18288 5108 18294 5120
rect 18417 5117 18429 5120
rect 18463 5117 18475 5151
rect 18417 5111 18475 5117
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 18690 5148 18696 5160
rect 18555 5120 18696 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 20254 5148 20260 5160
rect 20215 5120 20260 5148
rect 20254 5108 20260 5120
rect 20312 5148 20318 5160
rect 20993 5151 21051 5157
rect 20993 5148 21005 5151
rect 20312 5120 21005 5148
rect 20312 5108 20318 5120
rect 20993 5117 21005 5120
rect 21039 5117 21051 5151
rect 22462 5148 22468 5160
rect 22423 5120 22468 5148
rect 20993 5111 21051 5117
rect 22462 5108 22468 5120
rect 22520 5108 22526 5160
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23532 5120 23673 5148
rect 23532 5108 23538 5120
rect 23661 5117 23673 5120
rect 23707 5148 23719 5151
rect 24213 5151 24271 5157
rect 24213 5148 24225 5151
rect 23707 5120 24225 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24213 5117 24225 5120
rect 24259 5117 24271 5151
rect 24213 5111 24271 5117
rect 15562 5040 15568 5092
rect 15620 5080 15626 5092
rect 16485 5083 16543 5089
rect 16485 5080 16497 5083
rect 15620 5052 16497 5080
rect 15620 5040 15626 5052
rect 16485 5049 16497 5052
rect 16531 5080 16543 5083
rect 16574 5080 16580 5092
rect 16531 5052 16580 5080
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 20530 5080 20536 5092
rect 20491 5052 20536 5080
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 14001 5015 14059 5021
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14047 4984 14933 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 14921 4981 14933 4984
rect 14967 5012 14979 5015
rect 15378 5012 15384 5024
rect 14967 4984 15384 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 17678 5012 17684 5024
rect 17639 4984 17684 5012
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 25314 5012 25320 5024
rect 23891 4984 25320 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 25314 4972 25320 4984
rect 25372 4972 25378 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1854 4808 1860 4820
rect 1815 4780 1860 4808
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 2280 4780 2329 4808
rect 2280 4768 2286 4780
rect 2317 4777 2329 4780
rect 2363 4808 2375 4811
rect 2682 4808 2688 4820
rect 2363 4780 2688 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2832 4780 3249 4808
rect 2832 4768 2838 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5592 4780 5825 4808
rect 5592 4768 5598 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 5905 4811 5963 4817
rect 5905 4777 5917 4811
rect 5951 4808 5963 4811
rect 5994 4808 6000 4820
rect 5951 4780 6000 4808
rect 5951 4777 5963 4780
rect 5905 4771 5963 4777
rect 2961 4743 3019 4749
rect 2961 4709 2973 4743
rect 3007 4740 3019 4743
rect 3050 4740 3056 4752
rect 3007 4712 3056 4740
rect 3007 4709 3019 4712
rect 2961 4703 3019 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 4338 4740 4344 4752
rect 4299 4712 4344 4740
rect 4338 4700 4344 4712
rect 4396 4700 4402 4752
rect 5828 4740 5856 4771
rect 5994 4768 6000 4780
rect 6052 4808 6058 4820
rect 6822 4808 6828 4820
rect 6052 4780 6828 4808
rect 6052 4768 6058 4780
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 7558 4808 7564 4820
rect 7423 4780 7564 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8018 4808 8024 4820
rect 7979 4780 8024 4808
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9582 4808 9588 4820
rect 9539 4780 9588 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 9916 4780 10885 4808
rect 9916 4768 9922 4780
rect 10873 4777 10885 4780
rect 10919 4808 10931 4811
rect 11146 4808 11152 4820
rect 10919 4780 11152 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11422 4808 11428 4820
rect 11383 4780 11428 4808
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 12158 4808 12164 4820
rect 11839 4780 12164 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13538 4808 13544 4820
rect 13035 4780 13544 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13722 4808 13728 4820
rect 13679 4780 13728 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14792 4780 15025 4808
rect 14792 4768 14798 4780
rect 15013 4777 15025 4780
rect 15059 4808 15071 4811
rect 15286 4808 15292 4820
rect 15059 4780 15292 4808
rect 15059 4777 15071 4780
rect 15013 4771 15071 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 16390 4808 16396 4820
rect 16172 4780 16396 4808
rect 16172 4768 16178 4780
rect 16390 4768 16396 4780
rect 16448 4808 16454 4820
rect 16945 4811 17003 4817
rect 16945 4808 16957 4811
rect 16448 4780 16957 4808
rect 16448 4768 16454 4780
rect 16945 4777 16957 4780
rect 16991 4777 17003 4811
rect 16945 4771 17003 4777
rect 17405 4811 17463 4817
rect 17405 4777 17417 4811
rect 17451 4808 17463 4811
rect 17586 4808 17592 4820
rect 17451 4780 17592 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 17862 4808 17868 4820
rect 17819 4780 17868 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 19150 4808 19156 4820
rect 19111 4780 19156 4808
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 20070 4808 20076 4820
rect 20031 4780 20076 4808
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22554 4808 22560 4820
rect 22152 4780 22560 4808
rect 22152 4768 22158 4780
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 6178 4740 6184 4752
rect 5828 4712 6184 4740
rect 6178 4700 6184 4712
rect 6236 4700 6242 4752
rect 6914 4740 6920 4752
rect 6875 4712 6920 4740
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 9950 4700 9956 4752
rect 10008 4740 10014 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 10008 4712 10057 4740
rect 10008 4700 10014 4712
rect 10045 4709 10057 4712
rect 10091 4740 10103 4743
rect 10134 4740 10140 4752
rect 10091 4712 10140 4740
rect 10091 4709 10103 4712
rect 10045 4703 10103 4709
rect 10134 4700 10140 4712
rect 10192 4700 10198 4752
rect 11330 4740 11336 4752
rect 11291 4712 11336 4740
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 17604 4740 17632 4768
rect 11756 4712 14780 4740
rect 17604 4712 18368 4740
rect 11756 4700 11762 4712
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 2222 4672 2228 4684
rect 1544 4644 2228 4672
rect 1544 4632 1550 4644
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 4062 4632 4068 4684
rect 4120 4681 4126 4684
rect 4120 4675 4133 4681
rect 4121 4672 4133 4675
rect 7469 4675 7527 4681
rect 4121 4644 4165 4672
rect 4121 4641 4133 4644
rect 4120 4635 4133 4641
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 7834 4672 7840 4684
rect 7515 4644 7840 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 4120 4632 4126 4635
rect 7834 4632 7840 4644
rect 7892 4672 7898 4684
rect 8294 4672 8300 4684
rect 7892 4644 8300 4672
rect 7892 4632 7898 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 2372 4576 2421 4604
rect 2372 4564 2378 4576
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 4080 4604 4108 4632
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4080 4576 4813 4604
rect 2409 4567 2467 4573
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 6086 4604 6092 4616
rect 6047 4576 6092 4604
rect 4801 4567 4859 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 7650 4604 7656 4616
rect 7611 4576 7656 4604
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9490 4604 9496 4616
rect 8619 4576 9496 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 10008 4576 10149 4604
rect 10008 4564 10014 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10686 4604 10692 4616
rect 10367 4576 10692 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 5261 4539 5319 4545
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5534 4536 5540 4548
rect 5307 4508 5540 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 9398 4496 9404 4548
rect 9456 4536 9462 4548
rect 10336 4536 10364 4567
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11992 4613 12020 4712
rect 14752 4681 14780 4712
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 14737 4675 14795 4681
rect 13587 4644 14320 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 14292 4616 14320 4644
rect 14737 4641 14749 4675
rect 14783 4672 14795 4675
rect 14918 4672 14924 4684
rect 14783 4644 14924 4672
rect 14783 4641 14795 4644
rect 14737 4635 14795 4641
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15832 4675 15890 4681
rect 15832 4641 15844 4675
rect 15878 4672 15890 4675
rect 16114 4672 16120 4684
rect 15878 4644 16120 4672
rect 15878 4641 15890 4644
rect 15832 4635 15890 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 17954 4632 17960 4684
rect 18012 4672 18018 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 18012 4644 18153 4672
rect 18012 4632 18018 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 9456 4508 10364 4536
rect 9456 4496 9462 4508
rect 11790 4496 11796 4548
rect 11848 4536 11854 4548
rect 11900 4536 11928 4567
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13872 4576 14105 4604
rect 13872 4564 13878 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14093 4567 14151 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4573 15623 4607
rect 18230 4604 18236 4616
rect 18191 4576 18236 4604
rect 15565 4567 15623 4573
rect 11848 4508 11928 4536
rect 11848 4496 11854 4508
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 15580 4536 15608 4567
rect 18230 4564 18236 4576
rect 18288 4564 18294 4616
rect 18340 4613 18368 4712
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 19613 4743 19671 4749
rect 19613 4740 19625 4743
rect 19484 4712 19625 4740
rect 19484 4700 19490 4712
rect 19613 4709 19625 4712
rect 19659 4709 19671 4743
rect 19613 4703 19671 4709
rect 19337 4675 19395 4681
rect 19337 4641 19349 4675
rect 19383 4672 19395 4675
rect 19518 4672 19524 4684
rect 19383 4644 19524 4672
rect 19383 4641 19395 4644
rect 19337 4635 19395 4641
rect 19518 4632 19524 4644
rect 19576 4632 19582 4684
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 20990 4672 20996 4684
rect 20588 4644 20996 4672
rect 20588 4632 20594 4644
rect 20990 4632 20996 4644
rect 21048 4672 21054 4684
rect 21177 4675 21235 4681
rect 21177 4672 21189 4675
rect 21048 4644 21189 4672
rect 21048 4632 21054 4644
rect 21177 4641 21189 4644
rect 21223 4641 21235 4675
rect 21177 4635 21235 4641
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 22152 4644 22293 4672
rect 22152 4632 22158 4644
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 20070 4564 20076 4616
rect 20128 4604 20134 4616
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 20128 4576 20453 4604
rect 20128 4564 20134 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 14240 4508 15608 4536
rect 14240 4496 14246 4508
rect 20714 4496 20720 4548
rect 20772 4536 20778 4548
rect 20772 4508 21864 4536
rect 20772 4496 20778 4508
rect 21836 4480 21864 4508
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4468 1731 4471
rect 2130 4468 2136 4480
rect 1719 4440 2136 4468
rect 1719 4437 1731 4440
rect 1673 4431 1731 4437
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 3694 4468 3700 4480
rect 3655 4440 3700 4468
rect 3694 4428 3700 4440
rect 3752 4428 3758 4480
rect 5442 4468 5448 4480
rect 5403 4440 5448 4468
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 6454 4468 6460 4480
rect 6415 4440 6460 4468
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 8478 4468 8484 4480
rect 8439 4440 8484 4468
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9674 4468 9680 4480
rect 9635 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 12529 4471 12587 4477
rect 12529 4437 12541 4471
rect 12575 4468 12587 4471
rect 12894 4468 12900 4480
rect 12575 4440 12900 4468
rect 12575 4437 12587 4440
rect 12529 4431 12587 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 14734 4468 14740 4480
rect 14424 4440 14740 4468
rect 14424 4428 14430 4440
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 18782 4468 18788 4480
rect 18743 4440 18788 4468
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 21361 4471 21419 4477
rect 21361 4437 21373 4471
rect 21407 4468 21419 4471
rect 21634 4468 21640 4480
rect 21407 4440 21640 4468
rect 21407 4437 21419 4440
rect 21361 4431 21419 4437
rect 21634 4428 21640 4440
rect 21692 4428 21698 4480
rect 21818 4468 21824 4480
rect 21779 4440 21824 4468
rect 21818 4428 21824 4440
rect 21876 4428 21882 4480
rect 22462 4468 22468 4480
rect 22423 4440 22468 4468
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 2280 4236 3004 4264
rect 2280 4224 2286 4236
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1762 4128 1768 4140
rect 1452 4100 1768 4128
rect 1452 4088 1458 4100
rect 1762 4088 1768 4100
rect 1820 4128 1826 4140
rect 1949 4131 2007 4137
rect 1949 4128 1961 4131
rect 1820 4100 1961 4128
rect 1820 4088 1826 4100
rect 1949 4097 1961 4100
rect 1995 4097 2007 4131
rect 2976 4128 3004 4236
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 3844 4236 6561 4264
rect 3844 4224 3850 4236
rect 6549 4233 6561 4236
rect 6595 4264 6607 4267
rect 7282 4264 7288 4276
rect 6595 4236 7288 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 7926 4264 7932 4276
rect 7576 4236 7932 4264
rect 7576 4208 7604 4236
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 13998 4264 14004 4276
rect 13959 4236 14004 4264
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19429 4267 19487 4273
rect 19429 4264 19441 4267
rect 19392 4236 19441 4264
rect 19392 4224 19398 4236
rect 19429 4233 19441 4236
rect 19475 4233 19487 4267
rect 19429 4227 19487 4233
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 20625 4267 20683 4273
rect 20625 4264 20637 4267
rect 19576 4236 20637 4264
rect 19576 4224 19582 4236
rect 20625 4233 20637 4236
rect 20671 4233 20683 4267
rect 20990 4264 20996 4276
rect 20951 4236 20996 4264
rect 20625 4227 20683 4233
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 3326 4196 3332 4208
rect 3239 4168 3332 4196
rect 3326 4156 3332 4168
rect 3384 4196 3390 4208
rect 6086 4196 6092 4208
rect 3384 4168 4660 4196
rect 3384 4156 3390 4168
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 2976 4100 3985 4128
rect 1949 4091 2007 4097
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4632 4060 4660 4168
rect 5460 4168 6092 4196
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5460 4128 5488 4168
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 7558 4196 7564 4208
rect 6840 4168 7564 4196
rect 5123 4100 5488 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5592 4100 5733 4128
rect 5592 4088 5598 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 6273 4131 6331 4137
rect 6273 4097 6285 4131
rect 6319 4128 6331 4131
rect 6840 4128 6868 4168
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 7708 4168 8248 4196
rect 7708 4156 7714 4168
rect 6319 4100 6868 4128
rect 7837 4131 7895 4137
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 8018 4128 8024 4140
rect 7883 4100 8024 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8220 4128 8248 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9030 4196 9036 4208
rect 8352 4168 9036 4196
rect 8352 4156 8358 4168
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 9122 4156 9128 4208
rect 9180 4196 9186 4208
rect 11698 4196 11704 4208
rect 9180 4168 9628 4196
rect 9180 4156 9186 4168
rect 9324 4137 9352 4168
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8220 4100 8585 4128
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9600 4128 9628 4168
rect 11072 4168 11704 4196
rect 9766 4128 9772 4140
rect 9600 4100 9772 4128
rect 9309 4091 9367 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4128 10747 4131
rect 11072 4128 11100 4168
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 18230 4196 18236 4208
rect 17880 4168 18236 4196
rect 11330 4128 11336 4140
rect 10735 4100 11100 4128
rect 11291 4100 11336 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 17770 4128 17776 4140
rect 17731 4100 17776 4128
rect 12989 4091 13047 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 4632 4032 5304 4060
rect 2216 3995 2274 4001
rect 2216 3961 2228 3995
rect 2262 3992 2274 3995
rect 3234 3992 3240 4004
rect 2262 3964 3240 3992
rect 2262 3961 2274 3964
rect 2216 3955 2274 3961
rect 3234 3952 3240 3964
rect 3292 3992 3298 4004
rect 3292 3964 3740 3992
rect 3292 3952 3298 3964
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 2314 3924 2320 3936
rect 1903 3896 2320 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 3712 3933 3740 3964
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 3786 3924 3792 3936
rect 3743 3896 3792 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4154 3924 4160 3936
rect 4115 3896 4160 3924
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4890 3924 4896 3936
rect 4755 3896 4896 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5276 3924 5304 4032
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5408 4032 5641 4060
rect 5408 4020 5414 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 5629 4023 5687 4029
rect 7024 4032 7665 4060
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 5718 3992 5724 4004
rect 5583 3964 5724 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 5718 3952 5724 3964
rect 5776 3992 5782 4004
rect 6454 3992 6460 4004
rect 5776 3964 6460 3992
rect 5776 3952 5782 3964
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 7024 3936 7052 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8444 4032 9137 4060
rect 8444 4020 8450 4032
rect 9125 4029 9137 4032
rect 9171 4060 9183 4063
rect 9582 4060 9588 4072
rect 9171 4032 9588 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4060 11207 4063
rect 11238 4060 11244 4072
rect 11195 4032 11244 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13630 4060 13636 4072
rect 12851 4032 13636 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14240 4032 14289 4060
rect 14240 4020 14246 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 15344 4032 16497 4060
rect 15344 4020 15350 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 16632 4032 17509 4060
rect 16632 4020 16638 4032
rect 17497 4029 17509 4032
rect 17543 4060 17555 4063
rect 17880 4060 17908 4168
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 20162 4156 20168 4208
rect 20220 4196 20226 4208
rect 20220 4168 20300 4196
rect 20220 4156 20226 4168
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 17543 4032 17908 4060
rect 17972 4100 18613 4128
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 8294 3992 8300 4004
rect 7208 3964 8300 3992
rect 6086 3924 6092 3936
rect 5276 3896 6092 3924
rect 6086 3884 6092 3896
rect 6144 3924 6150 3936
rect 6270 3924 6276 3936
rect 6144 3896 6276 3924
rect 6144 3884 6150 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7208 3933 7236 3964
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 8536 3964 9229 3992
rect 8536 3952 8542 3964
rect 9217 3961 9229 3964
rect 9263 3961 9275 3995
rect 9217 3955 9275 3961
rect 11532 3964 12480 3992
rect 11532 3936 11560 3964
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7340 3896 7573 3924
rect 7340 3884 7346 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 7561 3887 7619 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9732 3896 9781 3924
rect 9732 3884 9738 3896
rect 9769 3893 9781 3896
rect 9815 3924 9827 3927
rect 9950 3924 9956 3936
rect 9815 3896 9956 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10781 3927 10839 3933
rect 10781 3893 10793 3927
rect 10827 3924 10839 3927
rect 10870 3924 10876 3936
rect 10827 3896 10876 3924
rect 10827 3893 10839 3896
rect 10781 3887 10839 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11241 3927 11299 3933
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11514 3924 11520 3936
rect 11287 3896 11520 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12452 3933 12480 3964
rect 12710 3952 12716 4004
rect 12768 3992 12774 4004
rect 13725 3995 13783 4001
rect 13725 3992 13737 3995
rect 12768 3964 13737 3992
rect 12768 3952 12774 3964
rect 13725 3961 13737 3964
rect 13771 3992 13783 3995
rect 13814 3992 13820 4004
rect 13771 3964 13820 3992
rect 13771 3961 13783 3964
rect 13725 3955 13783 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 14522 3995 14580 4001
rect 14522 3992 14534 3995
rect 14424 3964 14534 3992
rect 14424 3952 14430 3964
rect 14522 3961 14534 3964
rect 14568 3961 14580 3995
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 14522 3955 14580 3961
rect 15580 3964 16313 3992
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12437 3887 12495 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 15580 3924 15608 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16758 3992 16764 4004
rect 16719 3964 16764 3992
rect 16301 3955 16359 3961
rect 13596 3896 15608 3924
rect 15657 3927 15715 3933
rect 13596 3884 13602 3896
rect 15657 3893 15669 3927
rect 15703 3924 15715 3927
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15703 3896 16037 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 16025 3893 16037 3896
rect 16071 3924 16083 3927
rect 16114 3924 16120 3936
rect 16071 3896 16120 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16316 3924 16344 3955
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 17972 3924 18000 4100
rect 18601 4097 18613 4100
rect 18647 4128 18659 4131
rect 19242 4128 19248 4140
rect 18647 4100 19248 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20272 4137 20300 4168
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 18046 4020 18052 4072
rect 18104 4060 18110 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18104 4032 18429 4060
rect 18104 4020 18110 4032
rect 18417 4029 18429 4032
rect 18463 4060 18475 4063
rect 18782 4060 18788 4072
rect 18463 4032 18788 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19978 4060 19984 4072
rect 19392 4032 19984 4060
rect 19392 4020 19398 4032
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 21174 4060 21180 4072
rect 21135 4032 21180 4060
rect 21174 4020 21180 4032
rect 21232 4060 21238 4072
rect 21729 4063 21787 4069
rect 21729 4060 21741 4063
rect 21232 4032 21741 4060
rect 21232 4020 21238 4032
rect 21729 4029 21741 4032
rect 21775 4029 21787 4063
rect 22278 4060 22284 4072
rect 22239 4032 22284 4060
rect 21729 4023 21787 4029
rect 22278 4020 22284 4032
rect 22336 4060 22342 4072
rect 22833 4063 22891 4069
rect 22833 4060 22845 4063
rect 22336 4032 22845 4060
rect 22336 4020 22342 4032
rect 22833 4029 22845 4032
rect 22879 4029 22891 4063
rect 22833 4023 22891 4029
rect 18138 3952 18144 4004
rect 18196 3992 18202 4004
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 18196 3964 18521 3992
rect 18196 3952 18202 3964
rect 18509 3961 18521 3964
rect 18555 3992 18567 3995
rect 19061 3995 19119 4001
rect 19061 3992 19073 3995
rect 18555 3964 19073 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 19061 3961 19073 3964
rect 19107 3961 19119 3995
rect 20346 3992 20352 4004
rect 19061 3955 19119 3961
rect 19628 3964 20352 3992
rect 16316 3896 18000 3924
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18322 3924 18328 3936
rect 18095 3896 18328 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 19628 3933 19656 3964
rect 20346 3952 20352 3964
rect 20404 3952 20410 4004
rect 22370 3992 22376 4004
rect 21376 3964 22376 3992
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3893 19671 3927
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 19613 3887 19671 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 21376 3933 21404 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3893 21419 3927
rect 21361 3887 21419 3893
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22462 3924 22468 3936
rect 22152 3896 22197 3924
rect 22423 3896 22468 3924
rect 22152 3884 22158 3896
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 2832 3692 3157 3720
rect 2832 3680 2838 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3145 3683 3203 3689
rect 3160 3652 3188 3683
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 5994 3720 6000 3732
rect 5859 3692 6000 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6178 3720 6184 3732
rect 6139 3692 6184 3720
rect 6178 3680 6184 3692
rect 6236 3680 6242 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 7742 3720 7748 3732
rect 7699 3692 7748 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8386 3720 8392 3732
rect 8347 3692 8392 3720
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 8849 3723 8907 3729
rect 8849 3689 8861 3723
rect 8895 3720 8907 3723
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8895 3692 9137 3720
rect 8895 3689 8907 3692
rect 8849 3683 8907 3689
rect 9125 3689 9137 3692
rect 9171 3720 9183 3723
rect 9398 3720 9404 3732
rect 9171 3692 9404 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11330 3720 11336 3732
rect 10919 3692 11336 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11330 3680 11336 3692
rect 11388 3680 11394 3732
rect 12434 3720 12440 3732
rect 11532 3692 12440 3720
rect 4062 3652 4068 3664
rect 3160 3624 4068 3652
rect 4062 3612 4068 3624
rect 4120 3652 4126 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 4120 3624 4322 3652
rect 4120 3612 4126 3624
rect 4310 3621 4322 3624
rect 4356 3621 4368 3655
rect 4310 3615 4368 3621
rect 5534 3612 5540 3664
rect 5592 3652 5598 3664
rect 6518 3655 6576 3661
rect 6518 3652 6530 3655
rect 5592 3624 6530 3652
rect 5592 3612 5598 3624
rect 6518 3621 6530 3624
rect 6564 3621 6576 3655
rect 6518 3615 6576 3621
rect 7834 3612 7840 3664
rect 7892 3652 7898 3664
rect 11532 3652 11560 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12584 3692 13093 3720
rect 12584 3680 12590 3692
rect 13081 3689 13093 3692
rect 13127 3720 13139 3723
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 13127 3692 13185 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3720 13415 3723
rect 13630 3720 13636 3732
rect 13403 3692 13636 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 15562 3720 15568 3732
rect 15523 3692 15568 3720
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 16022 3720 16028 3732
rect 15983 3692 16028 3720
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 17126 3720 17132 3732
rect 17087 3692 17132 3720
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17494 3720 17500 3732
rect 17455 3692 17500 3720
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18012 3692 18153 3720
rect 18012 3680 18018 3692
rect 18141 3689 18153 3692
rect 18187 3720 18199 3723
rect 19061 3723 19119 3729
rect 19061 3720 19073 3723
rect 18187 3692 19073 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 19061 3689 19073 3692
rect 19107 3689 19119 3723
rect 21450 3720 21456 3732
rect 21411 3692 21456 3720
rect 19061 3683 19119 3689
rect 21450 3680 21456 3692
rect 21508 3680 21514 3732
rect 21818 3720 21824 3732
rect 21779 3692 21824 3720
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 22554 3720 22560 3732
rect 22515 3692 22560 3720
rect 22554 3680 22560 3692
rect 22612 3720 22618 3732
rect 22925 3723 22983 3729
rect 22925 3720 22937 3723
rect 22612 3692 22937 3720
rect 22612 3680 22618 3692
rect 22925 3689 22937 3692
rect 22971 3689 22983 3723
rect 23658 3720 23664 3732
rect 23619 3692 23664 3720
rect 22925 3683 22983 3689
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 7892 3624 11560 3652
rect 7892 3612 7898 3624
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 13722 3652 13728 3664
rect 12124 3624 13728 3652
rect 12124 3612 12130 3624
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 15930 3652 15936 3664
rect 15843 3624 15936 3652
rect 15930 3612 15936 3624
rect 15988 3652 15994 3664
rect 16574 3652 16580 3664
rect 15988 3624 16580 3652
rect 15988 3612 15994 3624
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 18966 3652 18972 3664
rect 18555 3624 18972 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 18966 3612 18972 3624
rect 19024 3652 19030 3664
rect 19153 3655 19211 3661
rect 19153 3652 19165 3655
rect 19024 3624 19165 3652
rect 19024 3612 19030 3624
rect 19153 3621 19165 3624
rect 19199 3621 19211 3655
rect 19153 3615 19211 3621
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2038 3593 2044 3596
rect 2032 3584 2044 3593
rect 1951 3556 2044 3584
rect 2032 3547 2044 3556
rect 2096 3584 2102 3596
rect 2096 3556 2820 3584
rect 2038 3544 2044 3547
rect 2096 3544 2102 3556
rect 2792 3516 2820 3556
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 2924 3556 3433 3584
rect 2924 3544 2930 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8444 3556 8493 3584
rect 8444 3544 8450 3556
rect 8481 3553 8493 3556
rect 8527 3584 8539 3587
rect 8662 3584 8668 3596
rect 8527 3556 8668 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 10134 3584 10140 3596
rect 10095 3556 10140 3584
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 11416 3587 11474 3593
rect 11416 3553 11428 3587
rect 11462 3584 11474 3587
rect 11974 3584 11980 3596
rect 11462 3556 11980 3584
rect 11462 3553 11474 3556
rect 11416 3547 11474 3553
rect 11974 3544 11980 3556
rect 12032 3584 12038 3596
rect 12802 3584 12808 3596
rect 12032 3556 12808 3584
rect 12032 3544 12038 3556
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13817 3587 13875 3593
rect 13817 3553 13829 3587
rect 13863 3584 13875 3587
rect 13998 3584 14004 3596
rect 13863 3556 14004 3584
rect 13863 3553 13875 3556
rect 13817 3547 13875 3553
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 14550 3544 14556 3596
rect 14608 3584 14614 3596
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 14608 3556 16957 3584
rect 14608 3544 14614 3556
rect 16945 3553 16957 3556
rect 16991 3584 17003 3587
rect 17402 3584 17408 3596
rect 16991 3556 17408 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 17586 3584 17592 3596
rect 17547 3556 17592 3584
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 22002 3584 22008 3596
rect 21963 3556 22008 3584
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 23106 3584 23112 3596
rect 23067 3556 23112 3584
rect 23106 3544 23112 3556
rect 23164 3544 23170 3596
rect 3326 3516 3332 3528
rect 2792 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3804 3488 4077 3516
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 3804 3380 3832 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 4065 3479 4123 3485
rect 5083 3488 6285 3516
rect 4430 3380 4436 3392
rect 1820 3352 4436 3380
rect 1820 3340 1826 3352
rect 4430 3340 4436 3352
rect 4488 3380 4494 3392
rect 5083 3380 5111 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 8018 3516 8024 3528
rect 7931 3488 8024 3516
rect 6273 3479 6331 3485
rect 8018 3476 8024 3488
rect 8076 3516 8082 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8076 3488 8861 3516
rect 8076 3476 8082 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 11146 3516 11152 3528
rect 11107 3488 11152 3516
rect 8849 3479 8907 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13630 3516 13636 3528
rect 13127 3488 13636 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 13909 3519 13967 3525
rect 13909 3516 13921 3519
rect 13688 3488 13921 3516
rect 13688 3476 13694 3488
rect 13909 3485 13921 3488
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 14332 3488 15117 3516
rect 14332 3476 14338 3488
rect 15105 3485 15117 3488
rect 15151 3516 15163 3519
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 15151 3488 16221 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 16209 3485 16221 3488
rect 16255 3516 16267 3519
rect 16390 3516 16396 3528
rect 16255 3488 16396 3516
rect 16255 3485 16267 3488
rect 16209 3479 16267 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 17678 3516 17684 3528
rect 17639 3488 17684 3516
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 19242 3516 19248 3528
rect 19203 3488 19248 3516
rect 19242 3476 19248 3488
rect 19300 3516 19306 3528
rect 19705 3519 19763 3525
rect 19705 3516 19717 3519
rect 19300 3488 19717 3516
rect 19300 3476 19306 3488
rect 19705 3485 19717 3488
rect 19751 3516 19763 3519
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19751 3488 20085 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 20073 3485 20085 3488
rect 20119 3516 20131 3519
rect 20162 3516 20168 3528
rect 20119 3488 20168 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 18693 3451 18751 3457
rect 12492 3420 16804 3448
rect 12492 3408 12498 3420
rect 4488 3352 5111 3380
rect 5445 3383 5503 3389
rect 4488 3340 4494 3352
rect 5445 3349 5457 3383
rect 5491 3380 5503 3383
rect 5994 3380 6000 3392
rect 5491 3352 6000 3380
rect 5491 3349 5503 3352
rect 5445 3343 5503 3349
rect 5994 3340 6000 3352
rect 6052 3340 6058 3392
rect 8665 3383 8723 3389
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 8938 3380 8944 3392
rect 8711 3352 8944 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 12529 3383 12587 3389
rect 12529 3380 12541 3383
rect 11388 3352 12541 3380
rect 11388 3340 11394 3352
rect 12529 3349 12541 3352
rect 12575 3349 12587 3383
rect 12894 3380 12900 3392
rect 12855 3352 12900 3380
rect 12529 3343 12587 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 14366 3380 14372 3392
rect 14327 3352 14372 3380
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 16574 3380 16580 3392
rect 16535 3352 16580 3380
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 16776 3380 16804 3420
rect 18693 3417 18705 3451
rect 18739 3448 18751 3451
rect 18874 3448 18880 3460
rect 18739 3420 18880 3448
rect 18739 3417 18751 3420
rect 18693 3411 18751 3417
rect 18874 3408 18880 3420
rect 18932 3408 18938 3460
rect 20806 3408 20812 3460
rect 20864 3448 20870 3460
rect 22189 3451 22247 3457
rect 22189 3448 22201 3451
rect 20864 3420 22201 3448
rect 20864 3408 20870 3420
rect 22189 3417 22201 3420
rect 22235 3417 22247 3451
rect 22189 3411 22247 3417
rect 19426 3380 19432 3392
rect 16776 3352 19432 3380
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 20438 3380 20444 3392
rect 20399 3352 20444 3380
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 21082 3380 21088 3392
rect 21043 3352 21088 3380
rect 21082 3340 21088 3352
rect 21140 3340 21146 3392
rect 23290 3380 23296 3392
rect 23251 3352 23296 3380
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1394 3176 1400 3188
rect 1355 3148 1400 3176
rect 1394 3136 1400 3148
rect 1452 3136 1458 3188
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4172 3148 5479 3176
rect 2501 3111 2559 3117
rect 2501 3077 2513 3111
rect 2547 3108 2559 3111
rect 4172 3108 4200 3148
rect 2547 3080 4200 3108
rect 5451 3108 5479 3148
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5592 3148 5917 3176
rect 5592 3136 5598 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 8478 3176 8484 3188
rect 6963 3148 8484 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9732 3148 10609 3176
rect 9732 3136 9738 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 11974 3176 11980 3188
rect 11931 3148 11980 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 6089 3111 6147 3117
rect 6089 3108 6101 3111
rect 5451 3080 6101 3108
rect 2547 3077 2559 3080
rect 2501 3071 2559 3077
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2130 3040 2136 3052
rect 2087 3012 2136 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 3436 3049 3464 3080
rect 6089 3077 6101 3080
rect 6135 3077 6147 3111
rect 8018 3108 8024 3120
rect 7979 3080 8024 3108
rect 6089 3071 6147 3077
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 8386 3108 8392 3120
rect 8347 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 9858 3068 9864 3120
rect 9916 3108 9922 3120
rect 10137 3111 10195 3117
rect 10137 3108 10149 3111
rect 9916 3080 10149 3108
rect 9916 3068 9922 3080
rect 10137 3077 10149 3080
rect 10183 3077 10195 3111
rect 10137 3071 10195 3077
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3568 3012 3617 3040
rect 3568 3000 3574 3012
rect 3605 3009 3617 3012
rect 3651 3040 3663 3043
rect 3786 3040 3792 3052
rect 3651 3012 3792 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4488 3012 4537 3040
rect 4488 3000 4494 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 6972 3012 7573 3040
rect 6972 3000 6978 3012
rect 7561 3009 7573 3012
rect 7607 3040 7619 3043
rect 8036 3040 8064 3068
rect 7607 3012 8616 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 1728 2944 1777 2972
rect 1728 2932 1734 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3326 2972 3332 2984
rect 2915 2944 3332 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 3970 2972 3976 2984
rect 3804 2944 3976 2972
rect 3804 2916 3832 2944
rect 3970 2932 3976 2944
rect 4028 2972 4034 2984
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 4028 2944 6285 2972
rect 4028 2932 4034 2944
rect 6273 2941 6285 2944
rect 6319 2972 6331 2975
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6319 2944 7297 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 8478 2972 8484 2984
rect 8439 2944 8484 2972
rect 7285 2935 7343 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8588 2972 8616 3012
rect 8737 2975 8795 2981
rect 8737 2972 8749 2975
rect 8588 2944 8749 2972
rect 8737 2941 8749 2944
rect 8783 2941 8795 2975
rect 8737 2935 8795 2941
rect 3786 2864 3792 2916
rect 3844 2864 3850 2916
rect 4792 2907 4850 2913
rect 4792 2873 4804 2907
rect 4838 2904 4850 2907
rect 4890 2904 4896 2916
rect 4838 2876 4896 2904
rect 4838 2873 4850 2876
rect 4792 2867 4850 2873
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 5994 2904 6000 2916
rect 4948 2876 6000 2904
rect 4948 2864 4954 2876
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 6546 2904 6552 2916
rect 6507 2876 6552 2904
rect 6546 2864 6552 2876
rect 6604 2904 6610 2916
rect 7377 2907 7435 2913
rect 7377 2904 7389 2907
rect 6604 2876 7389 2904
rect 6604 2864 6610 2876
rect 7377 2873 7389 2876
rect 7423 2904 7435 2907
rect 9490 2904 9496 2916
rect 7423 2876 9496 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 10612 2904 10640 3139
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 10744 3080 11468 3108
rect 10744 3068 10750 3080
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11440 3049 11468 3080
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 11112 3012 11253 3040
rect 11112 3000 11118 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11425 3043 11483 3049
rect 11425 3009 11437 3043
rect 11471 3040 11483 3043
rect 11900 3040 11928 3139
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 13780 3148 14381 3176
rect 13780 3136 13786 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14369 3139 14427 3145
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15470 3176 15476 3188
rect 15243 3148 15476 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15657 3179 15715 3185
rect 15657 3145 15669 3179
rect 15703 3176 15715 3179
rect 16022 3176 16028 3188
rect 15703 3148 16028 3176
rect 15703 3145 15715 3148
rect 15657 3139 15715 3145
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 17221 3179 17279 3185
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 17494 3176 17500 3188
rect 17267 3148 17500 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18414 3176 18420 3188
rect 18095 3148 18420 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 19426 3136 19432 3148
rect 19484 3176 19490 3188
rect 20070 3176 20076 3188
rect 19484 3148 20076 3176
rect 19484 3136 19490 3148
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 20898 3176 20904 3188
rect 20859 3148 20904 3176
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 22002 3176 22008 3188
rect 21963 3148 22008 3176
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 23382 3176 23388 3188
rect 23164 3148 23388 3176
rect 23164 3136 23170 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15565 3111 15623 3117
rect 15565 3108 15577 3111
rect 15160 3080 15577 3108
rect 15160 3068 15166 3080
rect 15565 3077 15577 3080
rect 15611 3108 15623 3111
rect 15930 3108 15936 3120
rect 15611 3080 15936 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20622 3108 20628 3120
rect 19659 3080 20628 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 11471 3012 11928 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12032 3012 12848 3040
rect 12032 3000 12038 3012
rect 11146 2932 11152 2984
rect 11204 2972 11210 2984
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 11204 2944 12725 2972
rect 11204 2932 11210 2944
rect 12713 2941 12725 2944
rect 12759 2941 12771 2975
rect 12820 2972 12848 3012
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 16172 3012 16313 3040
rect 16172 3000 16178 3012
rect 16301 3009 16313 3012
rect 16347 3040 16359 3043
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16347 3012 16681 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17460 3012 18613 3040
rect 17460 3000 17466 3012
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 12969 2975 13027 2981
rect 12969 2972 12981 2975
rect 12820 2944 12981 2972
rect 12713 2935 12771 2941
rect 12969 2941 12981 2944
rect 13015 2941 13027 2975
rect 12969 2935 13027 2941
rect 10612 2876 11192 2904
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 2958 2836 2964 2848
rect 2919 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 6089 2839 6147 2845
rect 6089 2805 6101 2839
rect 6135 2836 6147 2839
rect 8110 2836 8116 2848
rect 6135 2808 8116 2836
rect 6135 2805 6147 2808
rect 6089 2799 6147 2805
rect 8110 2796 8116 2808
rect 8168 2836 8174 2848
rect 8386 2836 8392 2848
rect 8168 2808 8392 2836
rect 8168 2796 8174 2808
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 9824 2808 9873 2836
rect 9824 2796 9830 2808
rect 9861 2805 9873 2808
rect 9907 2836 9919 2839
rect 10686 2836 10692 2848
rect 9907 2808 10692 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 10781 2839 10839 2845
rect 10781 2805 10793 2839
rect 10827 2836 10839 2839
rect 10962 2836 10968 2848
rect 10827 2808 10968 2836
rect 10827 2805 10839 2808
rect 10781 2799 10839 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11164 2845 11192 2876
rect 11330 2864 11336 2916
rect 11388 2904 11394 2916
rect 11974 2904 11980 2916
rect 11388 2876 11980 2904
rect 11388 2864 11394 2876
rect 11974 2864 11980 2876
rect 12032 2904 12038 2916
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 12032 2876 12173 2904
rect 12032 2864 12038 2876
rect 12161 2873 12173 2876
rect 12207 2873 12219 2907
rect 12728 2904 12756 2935
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15620 2944 16037 2972
rect 15620 2932 15626 2944
rect 16025 2941 16037 2944
rect 16071 2941 16083 2975
rect 16025 2935 16083 2941
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 19628 2972 19656 3071
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3040 21511 3043
rect 22020 3040 22048 3136
rect 22649 3111 22707 3117
rect 22649 3077 22661 3111
rect 22695 3108 22707 3111
rect 23658 3108 23664 3120
rect 22695 3080 23664 3108
rect 22695 3077 22707 3080
rect 22649 3071 22707 3077
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 21499 3012 22048 3040
rect 21499 3009 21511 3012
rect 21453 3003 21511 3009
rect 20070 2972 20076 2984
rect 18463 2944 19656 2972
rect 20031 2944 20076 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 21177 2975 21235 2981
rect 21177 2941 21189 2975
rect 21223 2972 21235 2975
rect 21358 2972 21364 2984
rect 21223 2944 21364 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 22465 2975 22523 2981
rect 22465 2972 22477 2975
rect 22244 2944 22477 2972
rect 22244 2932 22250 2944
rect 22465 2941 22477 2944
rect 22511 2972 22523 2975
rect 23017 2975 23075 2981
rect 23017 2972 23029 2975
rect 22511 2944 23029 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 23017 2941 23029 2944
rect 23063 2941 23075 2975
rect 23017 2935 23075 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2972 23719 2975
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23707 2944 24225 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 14182 2904 14188 2916
rect 12728 2876 14188 2904
rect 12161 2867 12219 2873
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14734 2864 14740 2916
rect 14792 2904 14798 2916
rect 16117 2907 16175 2913
rect 16117 2904 16129 2907
rect 14792 2876 16129 2904
rect 14792 2864 14798 2876
rect 16117 2873 16129 2876
rect 16163 2904 16175 2907
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 16163 2876 17509 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 17497 2873 17509 2876
rect 17543 2904 17555 2907
rect 17586 2904 17592 2916
rect 17543 2876 17592 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 17586 2864 17592 2876
rect 17644 2864 17650 2916
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 18288 2876 18521 2904
rect 18288 2864 18294 2876
rect 18509 2873 18521 2876
rect 18555 2904 18567 2907
rect 20438 2904 20444 2916
rect 18555 2876 20444 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 13780 2808 14105 2836
rect 13780 2796 13786 2808
rect 14093 2805 14105 2808
rect 14139 2836 14151 2839
rect 14366 2836 14372 2848
rect 14139 2808 14372 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19061 2839 19119 2845
rect 19061 2836 19073 2839
rect 18748 2808 19073 2836
rect 18748 2796 18754 2808
rect 19061 2805 19073 2808
rect 19107 2805 19119 2839
rect 19978 2836 19984 2848
rect 19939 2808 19984 2836
rect 19061 2799 19119 2805
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 22554 2836 22560 2848
rect 22244 2808 22560 2836
rect 22244 2796 22250 2808
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 23842 2836 23848 2848
rect 23803 2808 23848 2836
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1946 2632 1952 2644
rect 1719 2604 1952 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 3510 2632 3516 2644
rect 2096 2604 2141 2632
rect 3471 2604 3516 2632
rect 2096 2592 2102 2604
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 3878 2564 3884 2576
rect 2915 2536 3884 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 5276 2564 5304 2595
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5592 2604 6285 2632
rect 5592 2592 5598 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 6273 2595 6331 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8352 2604 8585 2632
rect 8352 2592 8358 2604
rect 8573 2601 8585 2604
rect 8619 2632 8631 2635
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8619 2604 9137 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 10744 2604 10793 2632
rect 10744 2592 10750 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 10781 2595 10839 2601
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11333 2635 11391 2641
rect 11333 2632 11345 2635
rect 11020 2604 11345 2632
rect 11020 2592 11026 2604
rect 11333 2601 11345 2604
rect 11379 2601 11391 2635
rect 11333 2595 11391 2601
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 5276 2536 6745 2564
rect 6733 2533 6745 2536
rect 6779 2564 6791 2567
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 6779 2536 8493 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 11348 2564 11376 2595
rect 11422 2592 11428 2644
rect 11480 2632 11486 2644
rect 11974 2632 11980 2644
rect 11480 2604 11525 2632
rect 11935 2604 11980 2632
rect 11480 2592 11486 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 13446 2632 13452 2644
rect 13407 2604 13452 2632
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2632 14062 2644
rect 15102 2632 15108 2644
rect 14056 2604 15108 2632
rect 14056 2592 14062 2604
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 18012 2604 18061 2632
rect 18012 2592 18018 2604
rect 18049 2601 18061 2604
rect 18095 2632 18107 2635
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18095 2604 18797 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20772 2604 20821 2632
rect 20772 2592 20778 2604
rect 20809 2601 20821 2604
rect 20855 2601 20867 2635
rect 20809 2595 20867 2601
rect 22186 2592 22192 2644
rect 22244 2632 22250 2644
rect 22281 2635 22339 2641
rect 22281 2632 22293 2635
rect 22244 2604 22293 2632
rect 22244 2592 22250 2604
rect 22281 2601 22293 2604
rect 22327 2632 22339 2635
rect 23385 2635 23443 2641
rect 23385 2632 23397 2635
rect 22327 2604 23397 2632
rect 22327 2601 22339 2604
rect 22281 2595 22339 2601
rect 23385 2601 23397 2604
rect 23431 2601 23443 2635
rect 23385 2595 23443 2601
rect 12345 2567 12403 2573
rect 12345 2564 12357 2567
rect 11348 2536 12357 2564
rect 8481 2527 8539 2533
rect 12345 2533 12357 2536
rect 12391 2533 12403 2567
rect 12345 2527 12403 2533
rect 12621 2567 12679 2573
rect 12621 2533 12633 2567
rect 12667 2564 12679 2567
rect 13170 2564 13176 2576
rect 12667 2536 13176 2564
rect 12667 2533 12679 2536
rect 12621 2527 12679 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13464 2564 13492 2592
rect 14369 2567 14427 2573
rect 14369 2564 14381 2567
rect 13464 2536 14381 2564
rect 14369 2533 14381 2536
rect 14415 2533 14427 2567
rect 14369 2527 14427 2533
rect 14642 2524 14648 2576
rect 14700 2564 14706 2576
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14700 2536 14933 2564
rect 14700 2524 14706 2536
rect 14921 2533 14933 2536
rect 14967 2564 14979 2567
rect 14967 2536 15976 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 3694 2496 3700 2508
rect 2823 2468 3700 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 3789 2499 3847 2505
rect 3789 2465 3801 2499
rect 3835 2496 3847 2499
rect 5534 2496 5540 2508
rect 3835 2468 5540 2496
rect 3835 2465 3847 2468
rect 3789 2459 3847 2465
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3804 2428 3832 2459
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6086 2496 6092 2508
rect 5767 2468 6092 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 4982 2428 4988 2440
rect 3099 2400 3832 2428
rect 4895 2400 4988 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 4982 2388 4988 2400
rect 5040 2428 5046 2440
rect 5644 2428 5672 2459
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 15948 2505 15976 2536
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 9861 2499 9919 2505
rect 7055 2468 7696 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 5040 2400 5672 2428
rect 5905 2431 5963 2437
rect 5040 2388 5046 2400
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6822 2428 6828 2440
rect 5951 2400 6828 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 4433 2363 4491 2369
rect 4433 2329 4445 2363
rect 4479 2360 4491 2363
rect 5920 2360 5948 2391
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 4479 2332 5948 2360
rect 4479 2329 4491 2332
rect 4433 2323 4491 2329
rect 2406 2292 2412 2304
rect 2367 2264 2412 2292
rect 2406 2252 2412 2264
rect 2464 2252 2470 2304
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 2556 2264 4721 2292
rect 2556 2252 2562 2264
rect 4709 2261 4721 2264
rect 4755 2292 4767 2295
rect 4985 2295 5043 2301
rect 4985 2292 4997 2295
rect 4755 2264 4997 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 4985 2261 4997 2264
rect 5031 2261 5043 2295
rect 5166 2292 5172 2304
rect 5079 2264 5172 2292
rect 4985 2255 5043 2261
rect 5166 2252 5172 2264
rect 5224 2292 5230 2304
rect 6086 2292 6092 2304
rect 5224 2264 6092 2292
rect 5224 2252 5230 2264
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7668 2301 7696 2468
rect 9861 2465 9873 2499
rect 9907 2496 9919 2499
rect 11793 2499 11851 2505
rect 9907 2468 10548 2496
rect 9907 2465 9919 2468
rect 9861 2459 9919 2465
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 8067 2400 8769 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8757 2397 8769 2400
rect 8803 2428 8815 2431
rect 9766 2428 9772 2440
rect 8803 2400 9772 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10520 2437 10548 2468
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 11839 2468 13369 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 13357 2459 13415 2465
rect 15212 2468 15853 2496
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 11609 2431 11667 2437
rect 10551 2400 11560 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 9585 2363 9643 2369
rect 9585 2329 9597 2363
rect 9631 2360 9643 2363
rect 11532 2360 11560 2400
rect 11609 2397 11621 2431
rect 11655 2428 11667 2431
rect 11974 2428 11980 2440
rect 11655 2400 11980 2428
rect 11655 2397 11667 2400
rect 11609 2391 11667 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2428 13691 2431
rect 13722 2428 13728 2440
rect 13679 2400 13728 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 9631 2332 11008 2360
rect 11532 2332 12633 2360
rect 9631 2329 9643 2332
rect 9585 2323 9643 2329
rect 7653 2295 7711 2301
rect 7653 2261 7665 2295
rect 7699 2292 7711 2295
rect 7742 2292 7748 2304
rect 7699 2264 7748 2292
rect 7699 2261 7711 2264
rect 7653 2255 7711 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10980 2301 11008 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 13648 2360 13676 2391
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 12943 2332 13676 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 10965 2295 11023 2301
rect 10965 2261 10977 2295
rect 11011 2292 11023 2295
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11011 2264 11805 2292
rect 11011 2261 11023 2264
rect 10965 2255 11023 2261
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 12986 2292 12992 2304
rect 12947 2264 12992 2292
rect 11793 2255 11851 2261
rect 12986 2252 12992 2264
rect 13044 2252 13050 2304
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 15212 2301 15240 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 16298 2496 16304 2508
rect 15979 2468 16304 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 16298 2456 16304 2468
rect 16356 2456 16362 2508
rect 17034 2496 17040 2508
rect 16995 2468 17040 2496
rect 17034 2456 17040 2468
rect 17092 2496 17098 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17092 2468 17601 2496
rect 17092 2456 17098 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 18690 2496 18696 2508
rect 18651 2468 18696 2496
rect 17589 2459 17647 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19886 2496 19892 2508
rect 19847 2468 19892 2496
rect 19886 2456 19892 2468
rect 19944 2496 19950 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19944 2468 20453 2496
rect 19944 2456 19950 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20441 2459 20499 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21232 2468 21925 2496
rect 21232 2456 21238 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22244 2468 22477 2496
rect 22244 2456 22250 2468
rect 22465 2465 22477 2468
rect 22511 2496 22523 2499
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22511 2468 23029 2496
rect 22511 2465 22523 2468
rect 22465 2459 22523 2465
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 23017 2459 23075 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24084 2468 24593 2496
rect 24084 2456 24090 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 25130 2496 25136 2508
rect 25043 2468 25136 2496
rect 24581 2459 24639 2465
rect 25130 2456 25136 2468
rect 25188 2496 25194 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25188 2468 25697 2496
rect 25188 2456 25194 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 16022 2388 16028 2400
rect 16080 2428 16086 2440
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16080 2400 16497 2428
rect 16080 2388 16086 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17678 2428 17684 2440
rect 16991 2400 17684 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17678 2388 17684 2400
rect 17736 2428 17742 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 17736 2400 18889 2428
rect 17736 2388 17742 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 20772 2400 21373 2428
rect 20772 2388 20778 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 20073 2363 20131 2369
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 21818 2360 21824 2372
rect 20119 2332 21824 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 22649 2363 22707 2369
rect 22649 2329 22661 2363
rect 22695 2360 22707 2363
rect 24118 2360 24124 2372
rect 22695 2332 24124 2360
rect 22695 2329 22707 2332
rect 22649 2323 22707 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 13228 2264 15209 2292
rect 13228 2252 13234 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 15197 2255 15255 2261
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 19705 2295 19763 2301
rect 19705 2261 19717 2295
rect 19751 2292 19763 2295
rect 19978 2292 19984 2304
rect 19751 2264 19984 2292
rect 19751 2261 19763 2264
rect 19705 2255 19763 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 24213 2295 24271 2301
rect 24213 2292 24225 2295
rect 23532 2264 24225 2292
rect 23532 2252 23538 2264
rect 24213 2261 24225 2264
rect 24259 2261 24271 2295
rect 24213 2255 24271 2261
rect 24854 2252 24860 2304
rect 24912 2292 24918 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 24912 2264 25329 2292
rect 24912 2252 24918 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 6546 2088 6552 2100
rect 3200 2060 6552 2088
rect 3200 2048 3206 2060
rect 6546 2048 6552 2060
rect 6604 2048 6610 2100
rect 6546 552 6552 604
rect 6604 592 6610 604
rect 7374 592 7380 604
rect 6604 564 7380 592
rect 6604 552 6610 564
rect 7374 552 7380 564
rect 7432 552 7438 604
rect 9214 552 9220 604
rect 9272 592 9278 604
rect 9398 592 9404 604
rect 9272 564 9404 592
rect 9272 552 9278 564
rect 9398 552 9404 564
rect 9456 552 9462 604
rect 21634 552 21640 604
rect 21692 592 21698 604
rect 23106 592 23112 604
rect 21692 564 23112 592
rect 21692 552 21698 564
rect 23106 552 23112 564
rect 23164 552 23170 604
<< via1 >>
rect 4896 26460 4948 26512
rect 12624 26460 12676 26512
rect 3976 26324 4028 26376
rect 13728 26256 13780 26308
rect 2412 25984 2464 26036
rect 9680 25984 9732 26036
rect 7472 25916 7524 25968
rect 12440 25916 12492 25968
rect 3240 25848 3292 25900
rect 12532 25848 12584 25900
rect 3976 25780 4028 25832
rect 11244 25780 11296 25832
rect 3056 25712 3108 25764
rect 5356 25712 5408 25764
rect 4068 25644 4120 25696
rect 11060 25644 11112 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 4068 25440 4120 25492
rect 11060 25483 11112 25492
rect 11060 25449 11069 25483
rect 11069 25449 11103 25483
rect 11103 25449 11112 25483
rect 11060 25440 11112 25449
rect 7472 25372 7524 25424
rect 2412 25304 2464 25356
rect 4160 25304 4212 25356
rect 6828 25304 6880 25356
rect 7564 25347 7616 25356
rect 7564 25313 7573 25347
rect 7573 25313 7607 25347
rect 7607 25313 7616 25347
rect 7564 25304 7616 25313
rect 7840 25304 7892 25356
rect 10600 25304 10652 25356
rect 1860 25236 1912 25288
rect 1584 25168 1636 25220
rect 8392 25236 8444 25288
rect 12532 25304 12584 25356
rect 13360 25304 13412 25356
rect 13636 25304 13688 25356
rect 15476 25347 15528 25356
rect 15476 25313 15485 25347
rect 15485 25313 15519 25347
rect 15519 25313 15528 25347
rect 15476 25304 15528 25313
rect 24768 25168 24820 25220
rect 2780 25100 2832 25152
rect 5356 25143 5408 25152
rect 5356 25109 5365 25143
rect 5365 25109 5399 25143
rect 5399 25109 5408 25143
rect 5356 25100 5408 25109
rect 5540 25100 5592 25152
rect 7840 25100 7892 25152
rect 8300 25100 8352 25152
rect 13544 25143 13596 25152
rect 13544 25109 13553 25143
rect 13553 25109 13587 25143
rect 13587 25109 13596 25143
rect 13544 25100 13596 25109
rect 26516 25100 26568 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2412 24939 2464 24948
rect 2412 24905 2421 24939
rect 2421 24905 2455 24939
rect 2455 24905 2464 24939
rect 2412 24896 2464 24905
rect 2964 24896 3016 24948
rect 5356 24896 5408 24948
rect 5540 24896 5592 24948
rect 7564 24896 7616 24948
rect 10600 24939 10652 24948
rect 10600 24905 10609 24939
rect 10609 24905 10643 24939
rect 10643 24905 10652 24939
rect 10600 24896 10652 24905
rect 12624 24939 12676 24948
rect 12624 24905 12633 24939
rect 12633 24905 12667 24939
rect 12667 24905 12676 24939
rect 12624 24896 12676 24905
rect 13360 24939 13412 24948
rect 13360 24905 13369 24939
rect 13369 24905 13403 24939
rect 13403 24905 13412 24939
rect 13360 24896 13412 24905
rect 13728 24939 13780 24948
rect 13728 24905 13737 24939
rect 13737 24905 13771 24939
rect 13771 24905 13780 24939
rect 13728 24896 13780 24905
rect 15476 24896 15528 24948
rect 1860 24803 1912 24812
rect 1860 24769 1869 24803
rect 1869 24769 1903 24803
rect 1903 24769 1912 24803
rect 1860 24760 1912 24769
rect 4712 24803 4764 24812
rect 4712 24769 4721 24803
rect 4721 24769 4755 24803
rect 4755 24769 4764 24803
rect 4712 24760 4764 24769
rect 5540 24760 5592 24812
rect 6920 24828 6972 24880
rect 1584 24735 1636 24744
rect 1584 24701 1593 24735
rect 1593 24701 1627 24735
rect 1627 24701 1636 24735
rect 1584 24692 1636 24701
rect 7196 24760 7248 24812
rect 3516 24624 3568 24676
rect 6276 24692 6328 24744
rect 8576 24735 8628 24744
rect 4160 24667 4212 24676
rect 4160 24633 4169 24667
rect 4169 24633 4203 24667
rect 4203 24633 4212 24667
rect 4160 24624 4212 24633
rect 4620 24624 4672 24676
rect 8576 24701 8585 24735
rect 8585 24701 8619 24735
rect 8619 24701 8628 24735
rect 8576 24692 8628 24701
rect 9864 24692 9916 24744
rect 8852 24624 8904 24676
rect 4528 24556 4580 24608
rect 5172 24599 5224 24608
rect 5172 24565 5181 24599
rect 5181 24565 5215 24599
rect 5215 24565 5224 24599
rect 5172 24556 5224 24565
rect 5540 24599 5592 24608
rect 5540 24565 5549 24599
rect 5549 24565 5583 24599
rect 5583 24565 5592 24599
rect 5540 24556 5592 24565
rect 7564 24556 7616 24608
rect 8392 24599 8444 24608
rect 8392 24565 8401 24599
rect 8401 24565 8435 24599
rect 8435 24565 8444 24599
rect 8392 24556 8444 24565
rect 8760 24599 8812 24608
rect 8760 24565 8769 24599
rect 8769 24565 8803 24599
rect 8803 24565 8812 24599
rect 8760 24556 8812 24565
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 12164 24692 12216 24744
rect 13544 24735 13596 24744
rect 13544 24701 13553 24735
rect 13553 24701 13587 24735
rect 13587 24701 13596 24735
rect 13544 24692 13596 24701
rect 14188 24692 14240 24744
rect 15936 24624 15988 24676
rect 12072 24556 12124 24608
rect 13636 24556 13688 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 17040 24599 17092 24608
rect 17040 24565 17049 24599
rect 17049 24565 17083 24599
rect 17083 24565 17092 24599
rect 17040 24556 17092 24565
rect 17776 24556 17828 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 11244 24352 11296 24404
rect 16212 24352 16264 24404
rect 18512 24352 18564 24404
rect 18788 24395 18840 24404
rect 18788 24361 18797 24395
rect 18797 24361 18831 24395
rect 18831 24361 18840 24395
rect 18788 24352 18840 24361
rect 19984 24352 20036 24404
rect 22008 24352 22060 24404
rect 22192 24395 22244 24404
rect 22192 24361 22201 24395
rect 22201 24361 22235 24395
rect 22235 24361 22244 24395
rect 22192 24352 22244 24361
rect 4988 24284 5040 24336
rect 1952 24259 2004 24268
rect 1952 24225 1961 24259
rect 1961 24225 1995 24259
rect 1995 24225 2004 24259
rect 1952 24216 2004 24225
rect 2872 24148 2924 24200
rect 4436 24148 4488 24200
rect 5264 24216 5316 24268
rect 7196 24259 7248 24268
rect 7196 24225 7230 24259
rect 7230 24225 7248 24259
rect 7196 24216 7248 24225
rect 9956 24216 10008 24268
rect 11060 24216 11112 24268
rect 13452 24216 13504 24268
rect 15568 24216 15620 24268
rect 16672 24216 16724 24268
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18144 24216 18196 24268
rect 20076 24216 20128 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 22008 24259 22060 24268
rect 22008 24225 22017 24259
rect 22017 24225 22051 24259
rect 22051 24225 22060 24259
rect 22008 24216 22060 24225
rect 3424 24080 3476 24132
rect 3332 24012 3384 24064
rect 4344 24055 4396 24064
rect 4344 24021 4353 24055
rect 4353 24021 4387 24055
rect 4387 24021 4396 24055
rect 5448 24080 5500 24132
rect 6644 24080 6696 24132
rect 4344 24012 4396 24021
rect 6828 24012 6880 24064
rect 7288 24012 7340 24064
rect 8300 24055 8352 24064
rect 8300 24021 8309 24055
rect 8309 24021 8343 24055
rect 8343 24021 8352 24055
rect 8300 24012 8352 24021
rect 8576 24055 8628 24064
rect 8576 24021 8585 24055
rect 8585 24021 8619 24055
rect 8619 24021 8628 24055
rect 8576 24012 8628 24021
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 17868 24080 17920 24132
rect 10140 24012 10192 24064
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 11704 24012 11756 24064
rect 12716 24055 12768 24064
rect 12716 24021 12725 24055
rect 12725 24021 12759 24055
rect 12759 24021 12768 24055
rect 12716 24012 12768 24021
rect 14004 24012 14056 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2412 23851 2464 23860
rect 2412 23817 2421 23851
rect 2421 23817 2455 23851
rect 2455 23817 2464 23851
rect 2412 23808 2464 23817
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 4896 23808 4948 23860
rect 5448 23808 5500 23860
rect 6276 23851 6328 23860
rect 6276 23817 6285 23851
rect 6285 23817 6319 23851
rect 6319 23817 6328 23851
rect 6276 23808 6328 23817
rect 6644 23851 6696 23860
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 12072 23808 12124 23860
rect 15568 23808 15620 23860
rect 16764 23808 16816 23860
rect 19064 23808 19116 23860
rect 19524 23808 19576 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 23388 23808 23440 23860
rect 25320 23808 25372 23860
rect 2412 23604 2464 23656
rect 4436 23783 4488 23792
rect 4436 23749 4445 23783
rect 4445 23749 4479 23783
rect 4479 23749 4488 23783
rect 4436 23740 4488 23749
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 5540 23672 5592 23724
rect 3424 23647 3476 23656
rect 3424 23613 3433 23647
rect 3433 23613 3467 23647
rect 3467 23613 3476 23647
rect 3424 23604 3476 23613
rect 4160 23604 4212 23656
rect 7748 23647 7800 23656
rect 7748 23613 7757 23647
rect 7757 23613 7791 23647
rect 7791 23613 7800 23647
rect 7748 23604 7800 23613
rect 12716 23672 12768 23724
rect 10140 23647 10192 23656
rect 1860 23579 1912 23588
rect 1860 23545 1869 23579
rect 1869 23545 1903 23579
rect 1903 23545 1912 23579
rect 1860 23536 1912 23545
rect 4712 23536 4764 23588
rect 7196 23536 7248 23588
rect 10140 23613 10149 23647
rect 10149 23613 10183 23647
rect 10183 23613 10192 23647
rect 10140 23604 10192 23613
rect 11704 23604 11756 23656
rect 11888 23647 11940 23656
rect 11888 23613 11897 23647
rect 11897 23613 11931 23647
rect 11931 23613 11940 23647
rect 13728 23672 13780 23724
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 20904 23715 20956 23724
rect 20904 23681 20913 23715
rect 20913 23681 20947 23715
rect 20947 23681 20956 23715
rect 20904 23672 20956 23681
rect 11888 23604 11940 23613
rect 2688 23468 2740 23520
rect 8576 23536 8628 23588
rect 10784 23536 10836 23588
rect 12072 23536 12124 23588
rect 13452 23579 13504 23588
rect 13452 23545 13461 23579
rect 13461 23545 13495 23579
rect 13495 23545 13504 23579
rect 13452 23536 13504 23545
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 19064 23604 19116 23656
rect 20260 23647 20312 23656
rect 20260 23613 20269 23647
rect 20269 23613 20303 23647
rect 20303 23613 20312 23647
rect 20260 23604 20312 23613
rect 21088 23604 21140 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 23480 23604 23532 23656
rect 18144 23536 18196 23588
rect 8208 23468 8260 23520
rect 8392 23468 8444 23520
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 12900 23468 12952 23520
rect 14004 23468 14056 23520
rect 15384 23511 15436 23520
rect 15384 23477 15393 23511
rect 15393 23477 15427 23511
rect 15427 23477 15436 23511
rect 15384 23468 15436 23477
rect 16028 23511 16080 23520
rect 16028 23477 16037 23511
rect 16037 23477 16071 23511
rect 16071 23477 16080 23511
rect 16028 23468 16080 23477
rect 16672 23468 16724 23520
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 20076 23511 20128 23520
rect 20076 23477 20085 23511
rect 20085 23477 20119 23511
rect 20119 23477 20128 23511
rect 20076 23468 20128 23477
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 3424 23307 3476 23316
rect 3424 23273 3433 23307
rect 3433 23273 3467 23307
rect 3467 23273 3476 23307
rect 3424 23264 3476 23273
rect 8300 23264 8352 23316
rect 9128 23307 9180 23316
rect 9128 23273 9137 23307
rect 9137 23273 9171 23307
rect 9171 23273 9180 23307
rect 9128 23264 9180 23273
rect 10784 23307 10836 23316
rect 10784 23273 10793 23307
rect 10793 23273 10827 23307
rect 10827 23273 10836 23307
rect 10784 23264 10836 23273
rect 12716 23264 12768 23316
rect 13728 23264 13780 23316
rect 14096 23264 14148 23316
rect 20628 23264 20680 23316
rect 3240 23196 3292 23248
rect 11888 23196 11940 23248
rect 13912 23196 13964 23248
rect 17500 23196 17552 23248
rect 23388 23196 23440 23248
rect 1768 23171 1820 23180
rect 1768 23137 1777 23171
rect 1777 23137 1811 23171
rect 1811 23137 1820 23171
rect 1768 23128 1820 23137
rect 2688 23128 2740 23180
rect 4344 23171 4396 23180
rect 4344 23137 4378 23171
rect 4378 23137 4396 23171
rect 4344 23128 4396 23137
rect 7288 23171 7340 23180
rect 7288 23137 7297 23171
rect 7297 23137 7331 23171
rect 7331 23137 7340 23171
rect 7288 23128 7340 23137
rect 7380 23128 7432 23180
rect 8392 23128 8444 23180
rect 10324 23128 10376 23180
rect 11796 23128 11848 23180
rect 4068 23103 4120 23112
rect 4068 23069 4077 23103
rect 4077 23069 4111 23103
rect 4111 23069 4120 23103
rect 4068 23060 4120 23069
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 9312 22992 9364 23044
rect 9956 22992 10008 23044
rect 13544 23060 13596 23112
rect 15108 23128 15160 23180
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 16304 23171 16356 23180
rect 16304 23137 16313 23171
rect 16313 23137 16347 23171
rect 16347 23137 16356 23171
rect 16304 23128 16356 23137
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 19156 23171 19208 23180
rect 19156 23137 19165 23171
rect 19165 23137 19199 23171
rect 19199 23137 19208 23171
rect 19156 23128 19208 23137
rect 22376 23171 22428 23180
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 15384 23060 15436 23112
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 2412 22924 2464 22976
rect 3516 22924 3568 22976
rect 3884 22967 3936 22976
rect 3884 22933 3893 22967
rect 3893 22933 3927 22967
rect 3927 22933 3936 22967
rect 3884 22924 3936 22933
rect 5448 22967 5500 22976
rect 5448 22933 5457 22967
rect 5457 22933 5491 22967
rect 5491 22933 5500 22967
rect 5448 22924 5500 22933
rect 9496 22924 9548 22976
rect 12900 22967 12952 22976
rect 12900 22933 12909 22967
rect 12909 22933 12943 22967
rect 12943 22933 12952 22967
rect 12900 22924 12952 22933
rect 13084 22924 13136 22976
rect 20260 22967 20312 22976
rect 20260 22933 20269 22967
rect 20269 22933 20303 22967
rect 20303 22933 20312 22967
rect 20260 22924 20312 22933
rect 21088 22924 21140 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1768 22720 1820 22772
rect 5540 22720 5592 22772
rect 6644 22763 6696 22772
rect 6644 22729 6653 22763
rect 6653 22729 6687 22763
rect 6687 22729 6696 22763
rect 6644 22720 6696 22729
rect 7380 22763 7432 22772
rect 7380 22729 7389 22763
rect 7389 22729 7423 22763
rect 7423 22729 7432 22763
rect 7380 22720 7432 22729
rect 7840 22763 7892 22772
rect 7840 22729 7849 22763
rect 7849 22729 7883 22763
rect 7883 22729 7892 22763
rect 7840 22720 7892 22729
rect 8852 22763 8904 22772
rect 8852 22729 8861 22763
rect 8861 22729 8895 22763
rect 8895 22729 8904 22763
rect 8852 22720 8904 22729
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 9680 22720 9732 22772
rect 9956 22720 10008 22772
rect 10140 22720 10192 22772
rect 11888 22763 11940 22772
rect 11888 22729 11897 22763
rect 11897 22729 11931 22763
rect 11931 22729 11940 22763
rect 11888 22720 11940 22729
rect 12164 22763 12216 22772
rect 12164 22729 12173 22763
rect 12173 22729 12207 22763
rect 12207 22729 12216 22763
rect 12164 22720 12216 22729
rect 13544 22720 13596 22772
rect 13820 22720 13872 22772
rect 15384 22720 15436 22772
rect 19156 22763 19208 22772
rect 19156 22729 19165 22763
rect 19165 22729 19199 22763
rect 19199 22729 19208 22763
rect 19156 22720 19208 22729
rect 22376 22763 22428 22772
rect 22376 22729 22385 22763
rect 22385 22729 22419 22763
rect 22419 22729 22428 22763
rect 22376 22720 22428 22729
rect 2412 22584 2464 22636
rect 3240 22584 3292 22636
rect 3516 22584 3568 22636
rect 3424 22516 3476 22568
rect 3884 22559 3936 22568
rect 3884 22525 3893 22559
rect 3893 22525 3927 22559
rect 3927 22525 3936 22559
rect 3884 22516 3936 22525
rect 6920 22584 6972 22636
rect 8208 22584 8260 22636
rect 10324 22652 10376 22704
rect 11060 22652 11112 22704
rect 12624 22695 12676 22704
rect 12624 22661 12633 22695
rect 12633 22661 12667 22695
rect 12667 22661 12676 22695
rect 12624 22652 12676 22661
rect 11244 22627 11296 22636
rect 11244 22593 11253 22627
rect 11253 22593 11287 22627
rect 11287 22593 11296 22627
rect 11244 22584 11296 22593
rect 5448 22516 5500 22568
rect 9496 22516 9548 22568
rect 10784 22516 10836 22568
rect 11704 22584 11756 22636
rect 16028 22627 16080 22636
rect 12164 22516 12216 22568
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 1400 22448 1452 22500
rect 14096 22516 14148 22568
rect 15752 22559 15804 22568
rect 15752 22525 15761 22559
rect 15761 22525 15795 22559
rect 15795 22525 15804 22559
rect 15752 22516 15804 22525
rect 5264 22423 5316 22432
rect 5264 22389 5273 22423
rect 5273 22389 5307 22423
rect 5307 22389 5316 22423
rect 5264 22380 5316 22389
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 10876 22380 10928 22432
rect 13728 22448 13780 22500
rect 15292 22448 15344 22500
rect 17868 22448 17920 22500
rect 13912 22380 13964 22432
rect 16028 22380 16080 22432
rect 16304 22380 16356 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 4344 22219 4396 22228
rect 4344 22185 4353 22219
rect 4353 22185 4387 22219
rect 4387 22185 4396 22219
rect 4344 22176 4396 22185
rect 9496 22176 9548 22228
rect 13360 22176 13412 22228
rect 13728 22176 13780 22228
rect 2872 22108 2924 22160
rect 3056 22108 3108 22160
rect 5264 22108 5316 22160
rect 2504 21972 2556 22024
rect 4160 22040 4212 22092
rect 6276 22108 6328 22160
rect 7012 22151 7064 22160
rect 7012 22117 7021 22151
rect 7021 22117 7055 22151
rect 7055 22117 7064 22151
rect 7012 22108 7064 22117
rect 7104 22040 7156 22092
rect 7472 22040 7524 22092
rect 7748 22040 7800 22092
rect 9864 22040 9916 22092
rect 11428 22040 11480 22092
rect 12532 22083 12584 22092
rect 12532 22049 12541 22083
rect 12541 22049 12575 22083
rect 12575 22049 12584 22083
rect 12532 22040 12584 22049
rect 13728 22040 13780 22092
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 3424 21972 3476 22024
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 1860 21904 1912 21956
rect 4252 21904 4304 21956
rect 7288 21904 7340 21956
rect 8208 21904 8260 21956
rect 8576 22015 8628 22024
rect 8576 21981 8585 22015
rect 8585 21981 8619 22015
rect 8619 21981 8628 22015
rect 10140 22015 10192 22024
rect 8576 21972 8628 21981
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 11796 22015 11848 22024
rect 8760 21904 8812 21956
rect 1952 21879 2004 21888
rect 1952 21845 1961 21879
rect 1961 21845 1995 21879
rect 1995 21845 2004 21879
rect 1952 21836 2004 21845
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6828 21879 6880 21888
rect 6552 21836 6604 21845
rect 6828 21845 6837 21879
rect 6837 21845 6871 21879
rect 6871 21845 6880 21879
rect 6828 21836 6880 21845
rect 7748 21836 7800 21888
rect 8024 21879 8076 21888
rect 8024 21845 8033 21879
rect 8033 21845 8067 21879
rect 8067 21845 8076 21879
rect 8024 21836 8076 21845
rect 8392 21836 8444 21888
rect 11796 21981 11805 22015
rect 11805 21981 11839 22015
rect 11839 21981 11848 22015
rect 11796 21972 11848 21981
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 13452 21972 13504 22024
rect 15568 22083 15620 22092
rect 15568 22049 15602 22083
rect 15602 22049 15620 22083
rect 15568 22040 15620 22049
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 11244 21947 11296 21956
rect 11244 21913 11253 21947
rect 11253 21913 11287 21947
rect 11287 21913 11296 21947
rect 11244 21904 11296 21913
rect 14004 21904 14056 21956
rect 10876 21879 10928 21888
rect 10876 21845 10885 21879
rect 10885 21845 10919 21879
rect 10919 21845 10928 21879
rect 10876 21836 10928 21845
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 13636 21879 13688 21888
rect 13636 21845 13645 21879
rect 13645 21845 13679 21879
rect 13679 21845 13688 21879
rect 13636 21836 13688 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1400 21675 1452 21684
rect 1400 21641 1409 21675
rect 1409 21641 1443 21675
rect 1443 21641 1452 21675
rect 1400 21632 1452 21641
rect 2504 21675 2556 21684
rect 2504 21641 2513 21675
rect 2513 21641 2547 21675
rect 2547 21641 2556 21675
rect 2504 21632 2556 21641
rect 3056 21632 3108 21684
rect 5264 21632 5316 21684
rect 8484 21632 8536 21684
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 9956 21632 10008 21684
rect 11704 21632 11756 21684
rect 12164 21632 12216 21684
rect 14004 21632 14056 21684
rect 14096 21632 14148 21684
rect 1860 21496 1912 21548
rect 4252 21539 4304 21548
rect 1676 21428 1728 21480
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 6184 21564 6236 21616
rect 10232 21607 10284 21616
rect 10232 21573 10241 21607
rect 10241 21573 10275 21607
rect 10275 21573 10284 21607
rect 10232 21564 10284 21573
rect 4620 21496 4672 21548
rect 6920 21496 6972 21548
rect 11244 21496 11296 21548
rect 2412 21428 2464 21480
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 5448 21428 5500 21480
rect 8024 21428 8076 21480
rect 8208 21428 8260 21480
rect 8392 21471 8444 21480
rect 1492 21360 1544 21412
rect 2504 21360 2556 21412
rect 3332 21360 3384 21412
rect 1400 21292 1452 21344
rect 1952 21292 2004 21344
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 3700 21292 3752 21344
rect 7932 21360 7984 21412
rect 8392 21437 8426 21471
rect 8426 21437 8444 21471
rect 8392 21428 8444 21437
rect 11336 21428 11388 21480
rect 11612 21428 11664 21480
rect 13084 21496 13136 21548
rect 13360 21496 13412 21548
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 15568 21496 15620 21548
rect 12532 21428 12584 21480
rect 12164 21360 12216 21412
rect 16672 21428 16724 21480
rect 4804 21292 4856 21344
rect 6552 21292 6604 21344
rect 9956 21292 10008 21344
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 11428 21335 11480 21344
rect 11428 21301 11437 21335
rect 11437 21301 11471 21335
rect 11471 21301 11480 21335
rect 11428 21292 11480 21301
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 13820 21292 13872 21344
rect 15660 21292 15712 21344
rect 15936 21292 15988 21344
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1676 21088 1728 21140
rect 4160 21088 4212 21140
rect 4896 21131 4948 21140
rect 4896 21097 4905 21131
rect 4905 21097 4939 21131
rect 4939 21097 4948 21131
rect 4896 21088 4948 21097
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 8392 21131 8444 21140
rect 8392 21097 8401 21131
rect 8401 21097 8435 21131
rect 8435 21097 8444 21131
rect 8392 21088 8444 21097
rect 8760 21131 8812 21140
rect 8760 21097 8769 21131
rect 8769 21097 8803 21131
rect 8803 21097 8812 21131
rect 8760 21088 8812 21097
rect 9680 21088 9732 21140
rect 10692 21088 10744 21140
rect 11060 21131 11112 21140
rect 11060 21097 11069 21131
rect 11069 21097 11103 21131
rect 11103 21097 11112 21131
rect 11060 21088 11112 21097
rect 4436 21020 4488 21072
rect 1492 20952 1544 21004
rect 6000 21020 6052 21072
rect 7196 21020 7248 21072
rect 9496 21020 9548 21072
rect 9864 21020 9916 21072
rect 11336 21088 11388 21140
rect 12072 21131 12124 21140
rect 12072 21097 12081 21131
rect 12081 21097 12115 21131
rect 12115 21097 12124 21131
rect 12072 21088 12124 21097
rect 13452 21088 13504 21140
rect 13728 21088 13780 21140
rect 15384 21088 15436 21140
rect 11888 21020 11940 21072
rect 14096 21020 14148 21072
rect 5540 20952 5592 21004
rect 7104 20952 7156 21004
rect 9404 20995 9456 21004
rect 9404 20961 9413 20995
rect 9413 20961 9447 20995
rect 9447 20961 9456 20995
rect 9404 20952 9456 20961
rect 10232 20952 10284 21004
rect 12440 20995 12492 21004
rect 12440 20961 12449 20995
rect 12449 20961 12483 20995
rect 12483 20961 12492 20995
rect 12440 20952 12492 20961
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 2044 20748 2096 20800
rect 2596 20748 2648 20800
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 5448 20748 5500 20800
rect 6552 20791 6604 20800
rect 6552 20757 6561 20791
rect 6561 20757 6595 20791
rect 6595 20757 6604 20791
rect 6552 20748 6604 20757
rect 6828 20748 6880 20800
rect 8208 20816 8260 20868
rect 9496 20816 9548 20868
rect 12624 20927 12676 20936
rect 12624 20893 12633 20927
rect 12633 20893 12667 20927
rect 12667 20893 12676 20927
rect 12624 20884 12676 20893
rect 13820 20884 13872 20936
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 14556 20884 14608 20936
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 15568 20816 15620 20868
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 14740 20748 14792 20800
rect 16396 20748 16448 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2504 20544 2556 20596
rect 3240 20544 3292 20596
rect 6092 20544 6144 20596
rect 7196 20544 7248 20596
rect 9220 20587 9272 20596
rect 9220 20553 9229 20587
rect 9229 20553 9263 20587
rect 9263 20553 9272 20587
rect 9220 20544 9272 20553
rect 9864 20544 9916 20596
rect 12624 20544 12676 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 14096 20587 14148 20596
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 14556 20587 14608 20596
rect 14556 20553 14565 20587
rect 14565 20553 14599 20587
rect 14599 20553 14608 20587
rect 14556 20544 14608 20553
rect 15568 20544 15620 20596
rect 16120 20544 16172 20596
rect 8760 20476 8812 20528
rect 9404 20476 9456 20528
rect 15384 20476 15436 20528
rect 1860 20408 1912 20460
rect 3056 20408 3108 20460
rect 3516 20408 3568 20460
rect 4160 20451 4212 20460
rect 4160 20417 4169 20451
rect 4169 20417 4203 20451
rect 4203 20417 4212 20451
rect 4160 20408 4212 20417
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 4344 20340 4396 20392
rect 1952 20272 2004 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 1768 20204 1820 20256
rect 2596 20204 2648 20256
rect 3056 20247 3108 20256
rect 3056 20213 3065 20247
rect 3065 20213 3099 20247
rect 3099 20213 3108 20247
rect 3056 20204 3108 20213
rect 3608 20247 3660 20256
rect 3608 20213 3617 20247
rect 3617 20213 3651 20247
rect 3651 20213 3660 20247
rect 3608 20204 3660 20213
rect 4252 20204 4304 20256
rect 4436 20204 4488 20256
rect 6828 20383 6880 20392
rect 5448 20272 5500 20324
rect 6092 20272 6144 20324
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 11704 20408 11756 20460
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14691 20451
rect 14691 20417 14700 20451
rect 14648 20408 14700 20417
rect 7104 20383 7156 20392
rect 7104 20349 7138 20383
rect 7138 20349 7156 20383
rect 7104 20340 7156 20349
rect 7288 20272 7340 20324
rect 10232 20340 10284 20392
rect 15844 20383 15896 20392
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 11060 20272 11112 20324
rect 13084 20272 13136 20324
rect 5172 20247 5224 20256
rect 5172 20213 5181 20247
rect 5181 20213 5215 20247
rect 5215 20213 5224 20247
rect 5172 20204 5224 20213
rect 8944 20247 8996 20256
rect 8944 20213 8953 20247
rect 8953 20213 8987 20247
rect 8987 20213 8996 20247
rect 8944 20204 8996 20213
rect 11336 20204 11388 20256
rect 13820 20204 13872 20256
rect 14188 20204 14240 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1952 20000 2004 20052
rect 2688 20000 2740 20052
rect 4068 20000 4120 20052
rect 6000 20000 6052 20052
rect 7380 20000 7432 20052
rect 7932 20043 7984 20052
rect 7932 20009 7941 20043
rect 7941 20009 7975 20043
rect 7975 20009 7984 20043
rect 7932 20000 7984 20009
rect 9680 20043 9732 20052
rect 9680 20009 9689 20043
rect 9689 20009 9723 20043
rect 9723 20009 9732 20043
rect 9680 20000 9732 20009
rect 3884 19932 3936 19984
rect 4160 19932 4212 19984
rect 5172 19932 5224 19984
rect 5540 19932 5592 19984
rect 6552 19975 6604 19984
rect 6552 19941 6561 19975
rect 6561 19941 6595 19975
rect 6595 19941 6604 19975
rect 6552 19932 6604 19941
rect 10324 19932 10376 19984
rect 3792 19864 3844 19916
rect 7656 19864 7708 19916
rect 8392 19864 8444 19916
rect 9680 19864 9732 19916
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 7196 19796 7248 19848
rect 10140 19796 10192 19848
rect 11060 20000 11112 20052
rect 13176 20000 13228 20052
rect 13820 20043 13872 20052
rect 13820 20009 13829 20043
rect 13829 20009 13863 20043
rect 13863 20009 13872 20043
rect 13820 20000 13872 20009
rect 14556 20000 14608 20052
rect 11704 19932 11756 19984
rect 12440 19932 12492 19984
rect 14280 19932 14332 19984
rect 11336 19864 11388 19916
rect 14096 19864 14148 19916
rect 15200 19864 15252 19916
rect 15384 20000 15436 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 15384 19864 15436 19916
rect 13912 19839 13964 19848
rect 13912 19805 13921 19839
rect 13921 19805 13955 19839
rect 13955 19805 13964 19839
rect 13912 19796 13964 19805
rect 3976 19728 4028 19780
rect 5356 19728 5408 19780
rect 10692 19728 10744 19780
rect 10876 19728 10928 19780
rect 1492 19660 1544 19712
rect 2136 19660 2188 19712
rect 5172 19660 5224 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 13084 19728 13136 19780
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 3792 19499 3844 19508
rect 3792 19465 3801 19499
rect 3801 19465 3835 19499
rect 3835 19465 3844 19499
rect 3792 19456 3844 19465
rect 7196 19456 7248 19508
rect 7656 19456 7708 19508
rect 11336 19456 11388 19508
rect 12440 19499 12492 19508
rect 12440 19465 12449 19499
rect 12449 19465 12483 19499
rect 12483 19465 12492 19499
rect 12440 19456 12492 19465
rect 15476 19456 15528 19508
rect 1308 19388 1360 19440
rect 1584 19388 1636 19440
rect 3056 19388 3108 19440
rect 4068 19388 4120 19440
rect 13912 19431 13964 19440
rect 13912 19397 13921 19431
rect 13921 19397 13955 19431
rect 13955 19397 13964 19431
rect 13912 19388 13964 19397
rect 14372 19388 14424 19440
rect 3240 19320 3292 19372
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 1584 19252 1636 19304
rect 2688 19252 2740 19304
rect 3608 19252 3660 19304
rect 4068 19252 4120 19304
rect 6092 19320 6144 19372
rect 6552 19252 6604 19304
rect 7380 19320 7432 19372
rect 7840 19320 7892 19372
rect 7932 19320 7984 19372
rect 9404 19320 9456 19372
rect 10968 19320 11020 19372
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 7288 19252 7340 19304
rect 7564 19252 7616 19304
rect 9680 19252 9732 19304
rect 10324 19252 10376 19304
rect 11152 19252 11204 19304
rect 1676 19227 1728 19236
rect 1676 19193 1685 19227
rect 1685 19193 1719 19227
rect 1719 19193 1728 19227
rect 1676 19184 1728 19193
rect 5172 19184 5224 19236
rect 11336 19227 11388 19236
rect 11336 19193 11345 19227
rect 11345 19193 11379 19227
rect 11379 19193 11388 19227
rect 11336 19184 11388 19193
rect 12164 19252 12216 19304
rect 14280 19320 14332 19372
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 14648 19363 14700 19372
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 15844 19320 15896 19329
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 13636 19184 13688 19236
rect 14188 19184 14240 19236
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 3516 19116 3568 19168
rect 3608 19116 3660 19168
rect 3976 19116 4028 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 7748 19116 7800 19168
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 8208 19116 8260 19125
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 9312 19116 9364 19168
rect 9496 19116 9548 19168
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 12164 19159 12216 19168
rect 12164 19125 12173 19159
rect 12173 19125 12207 19159
rect 12207 19125 12216 19159
rect 12164 19116 12216 19125
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 14004 19159 14056 19168
rect 14004 19125 14013 19159
rect 14013 19125 14047 19159
rect 14047 19125 14056 19159
rect 14004 19116 14056 19125
rect 15384 19159 15436 19168
rect 15384 19125 15393 19159
rect 15393 19125 15427 19159
rect 15427 19125 15436 19159
rect 15384 19116 15436 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2780 18955 2832 18964
rect 2780 18921 2789 18955
rect 2789 18921 2823 18955
rect 2823 18921 2832 18955
rect 2780 18912 2832 18921
rect 3148 18912 3200 18964
rect 3884 18955 3936 18964
rect 3884 18921 3893 18955
rect 3893 18921 3927 18955
rect 3927 18921 3936 18955
rect 3884 18912 3936 18921
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 4712 18955 4764 18964
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 7012 18912 7064 18964
rect 8208 18912 8260 18964
rect 8300 18912 8352 18964
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 13084 18912 13136 18964
rect 13636 18955 13688 18964
rect 13636 18921 13645 18955
rect 13645 18921 13679 18955
rect 13679 18921 13688 18955
rect 13636 18912 13688 18921
rect 13728 18912 13780 18964
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 4528 18776 4580 18828
rect 5632 18776 5684 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 10324 18776 10376 18828
rect 10968 18819 11020 18828
rect 10968 18785 10991 18819
rect 10991 18785 11020 18819
rect 14004 18819 14056 18828
rect 10968 18776 11020 18785
rect 14004 18785 14013 18819
rect 14013 18785 14047 18819
rect 14047 18785 14056 18819
rect 14004 18776 14056 18785
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 3884 18708 3936 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 3516 18640 3568 18692
rect 1952 18572 2004 18624
rect 3332 18572 3384 18624
rect 5172 18572 5224 18624
rect 9404 18708 9456 18760
rect 6552 18572 6604 18624
rect 7196 18615 7248 18624
rect 7196 18581 7205 18615
rect 7205 18581 7239 18615
rect 7239 18581 7248 18615
rect 7196 18572 7248 18581
rect 7840 18572 7892 18624
rect 8300 18572 8352 18624
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 12808 18708 12860 18760
rect 14096 18708 14148 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 14648 18640 14700 18692
rect 16488 18708 16540 18760
rect 10876 18572 10928 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1400 18411 1452 18420
rect 1400 18377 1409 18411
rect 1409 18377 1443 18411
rect 1443 18377 1452 18411
rect 1400 18368 1452 18377
rect 2780 18368 2832 18420
rect 3976 18368 4028 18420
rect 4252 18368 4304 18420
rect 4804 18411 4856 18420
rect 4804 18377 4813 18411
rect 4813 18377 4847 18411
rect 4847 18377 4856 18411
rect 4804 18368 4856 18377
rect 5080 18411 5132 18420
rect 5080 18377 5089 18411
rect 5089 18377 5123 18411
rect 5123 18377 5132 18411
rect 5080 18368 5132 18377
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 9036 18368 9088 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10784 18411 10836 18420
rect 10784 18377 10793 18411
rect 10793 18377 10827 18411
rect 10827 18377 10836 18411
rect 10784 18368 10836 18377
rect 11060 18368 11112 18420
rect 8208 18300 8260 18352
rect 8392 18300 8444 18352
rect 11428 18368 11480 18420
rect 12532 18368 12584 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 2780 18232 2832 18284
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 9036 18232 9088 18284
rect 10324 18232 10376 18284
rect 1400 18164 1452 18216
rect 1860 18164 1912 18216
rect 5080 18164 5132 18216
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 7656 18164 7708 18216
rect 12072 18232 12124 18284
rect 12440 18343 12492 18352
rect 12440 18309 12449 18343
rect 12449 18309 12483 18343
rect 12483 18309 12492 18343
rect 12440 18300 12492 18309
rect 14096 18368 14148 18420
rect 15384 18368 15436 18420
rect 12992 18164 13044 18216
rect 14648 18207 14700 18216
rect 14648 18173 14682 18207
rect 14682 18173 14700 18207
rect 1952 18096 2004 18148
rect 2964 18139 3016 18148
rect 2964 18105 2973 18139
rect 2973 18105 3007 18139
rect 3007 18105 3016 18139
rect 2964 18096 3016 18105
rect 4528 18096 4580 18148
rect 14648 18164 14700 18173
rect 15752 18164 15804 18216
rect 14556 18096 14608 18148
rect 15660 18096 15712 18148
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2228 18028 2280 18080
rect 2504 18028 2556 18080
rect 7196 18028 7248 18080
rect 9404 18028 9456 18080
rect 11336 18028 11388 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 14648 18028 14700 18080
rect 14832 18028 14884 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2872 17824 2924 17876
rect 3516 17824 3568 17876
rect 4160 17824 4212 17876
rect 4528 17824 4580 17876
rect 6552 17824 6604 17876
rect 7840 17824 7892 17876
rect 1400 17756 1452 17808
rect 4068 17756 4120 17808
rect 10968 17824 11020 17876
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 14004 17867 14056 17876
rect 14004 17833 14013 17867
rect 14013 17833 14047 17867
rect 14047 17833 14056 17867
rect 14004 17824 14056 17833
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 14556 17824 14608 17876
rect 2872 17731 2924 17740
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 1860 17552 1912 17604
rect 2504 17552 2556 17604
rect 4712 17688 4764 17740
rect 6092 17688 6144 17740
rect 7656 17731 7708 17740
rect 7656 17697 7690 17731
rect 7690 17697 7708 17731
rect 7656 17688 7708 17697
rect 9588 17688 9640 17740
rect 10784 17688 10836 17740
rect 12072 17688 12124 17740
rect 16580 17824 16632 17876
rect 14832 17688 14884 17740
rect 15844 17688 15896 17740
rect 4896 17663 4948 17672
rect 4896 17629 4905 17663
rect 4905 17629 4939 17663
rect 4939 17629 4948 17663
rect 4896 17620 4948 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 6552 17620 6604 17672
rect 7380 17663 7432 17672
rect 7380 17629 7389 17663
rect 7389 17629 7423 17663
rect 7423 17629 7432 17663
rect 7380 17620 7432 17629
rect 10876 17620 10928 17672
rect 6276 17552 6328 17604
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 2688 17484 2740 17536
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 9404 17527 9456 17536
rect 9404 17493 9413 17527
rect 9413 17493 9447 17527
rect 9447 17493 9456 17527
rect 9404 17484 9456 17493
rect 11336 17527 11388 17536
rect 11336 17493 11345 17527
rect 11345 17493 11379 17527
rect 11379 17493 11388 17527
rect 11336 17484 11388 17493
rect 12164 17484 12216 17536
rect 12900 17484 12952 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1400 17280 1452 17332
rect 2780 17280 2832 17332
rect 3056 17280 3108 17332
rect 4252 17323 4304 17332
rect 4252 17289 4261 17323
rect 4261 17289 4295 17323
rect 4295 17289 4304 17323
rect 4252 17280 4304 17289
rect 4712 17323 4764 17332
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 5080 17280 5132 17332
rect 7840 17280 7892 17332
rect 5356 17212 5408 17264
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 9404 17280 9456 17332
rect 11336 17280 11388 17332
rect 9220 17212 9272 17264
rect 9956 17212 10008 17264
rect 11152 17212 11204 17264
rect 12900 17212 12952 17264
rect 9128 17144 9180 17196
rect 10968 17144 11020 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 16856 17187 16908 17196
rect 2228 17076 2280 17128
rect 4252 17076 4304 17128
rect 4804 17076 4856 17128
rect 848 17008 900 17060
rect 2872 17008 2924 17060
rect 5540 17008 5592 17060
rect 8300 17076 8352 17128
rect 8852 17076 8904 17128
rect 9312 17076 9364 17128
rect 9864 17076 9916 17128
rect 13176 17076 13228 17128
rect 13636 17076 13688 17128
rect 14096 17119 14148 17128
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 16672 17076 16724 17128
rect 9404 17008 9456 17060
rect 9956 17008 10008 17060
rect 11796 17051 11848 17060
rect 11796 17017 11805 17051
rect 11805 17017 11839 17051
rect 11839 17017 11848 17051
rect 11796 17008 11848 17017
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 4804 16940 4856 16992
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 6920 16940 6972 16992
rect 7656 16940 7708 16992
rect 9864 16940 9916 16992
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 15476 16983 15528 16992
rect 12440 16940 12492 16949
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 16580 16940 16632 16992
rect 16764 16940 16816 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 2228 16779 2280 16788
rect 2228 16745 2237 16779
rect 2237 16745 2271 16779
rect 2271 16745 2280 16779
rect 2228 16736 2280 16745
rect 3056 16736 3108 16788
rect 4804 16779 4856 16788
rect 4804 16745 4813 16779
rect 4813 16745 4847 16779
rect 4847 16745 4856 16779
rect 4804 16736 4856 16745
rect 4896 16736 4948 16788
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 7012 16736 7064 16788
rect 7748 16779 7800 16788
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 8208 16736 8260 16788
rect 8300 16736 8352 16788
rect 9956 16736 10008 16788
rect 10784 16736 10836 16788
rect 11244 16779 11296 16788
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 12072 16779 12124 16788
rect 12072 16745 12081 16779
rect 12081 16745 12115 16779
rect 12115 16745 12124 16779
rect 12072 16736 12124 16745
rect 12256 16779 12308 16788
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 12348 16736 12400 16788
rect 12532 16736 12584 16788
rect 14832 16736 14884 16788
rect 15752 16736 15804 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 2688 16668 2740 16720
rect 3332 16668 3384 16720
rect 2228 16600 2280 16652
rect 4804 16600 4856 16652
rect 5632 16668 5684 16720
rect 8852 16711 8904 16720
rect 8852 16677 8861 16711
rect 8861 16677 8895 16711
rect 8895 16677 8904 16711
rect 8852 16668 8904 16677
rect 9680 16668 9732 16720
rect 10048 16668 10100 16720
rect 15936 16668 15988 16720
rect 16396 16668 16448 16720
rect 5172 16600 5224 16652
rect 10232 16643 10284 16652
rect 10232 16609 10241 16643
rect 10241 16609 10275 16643
rect 10275 16609 10284 16643
rect 10232 16600 10284 16609
rect 11336 16600 11388 16652
rect 12532 16600 12584 16652
rect 15476 16600 15528 16652
rect 16856 16600 16908 16652
rect 2964 16532 3016 16584
rect 3700 16532 3752 16584
rect 7840 16575 7892 16584
rect 5264 16464 5316 16516
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 10048 16532 10100 16584
rect 12808 16575 12860 16584
rect 7380 16507 7432 16516
rect 7380 16473 7389 16507
rect 7389 16473 7423 16507
rect 7423 16473 7432 16507
rect 7380 16464 7432 16473
rect 9220 16464 9272 16516
rect 9956 16464 10008 16516
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 15844 16532 15896 16584
rect 17040 16532 17092 16584
rect 11704 16464 11756 16516
rect 12532 16464 12584 16516
rect 7564 16396 7616 16448
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 11980 16396 12032 16448
rect 13728 16396 13780 16448
rect 14096 16396 14148 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2688 16192 2740 16244
rect 4804 16192 4856 16244
rect 5448 16192 5500 16244
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 8576 16235 8628 16244
rect 8576 16201 8585 16235
rect 8585 16201 8619 16235
rect 8619 16201 8628 16235
rect 8576 16192 8628 16201
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 9864 16192 9916 16244
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 11704 16192 11756 16244
rect 12348 16192 12400 16244
rect 15844 16192 15896 16244
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 10232 16124 10284 16176
rect 12164 16124 12216 16176
rect 15936 16124 15988 16176
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 5540 16056 5592 16108
rect 6092 16056 6144 16108
rect 6920 16056 6972 16108
rect 7564 16056 7616 16108
rect 9956 16056 10008 16108
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 12992 16056 13044 16108
rect 13728 16056 13780 16108
rect 16580 16099 16632 16108
rect 16580 16065 16589 16099
rect 16589 16065 16623 16099
rect 16623 16065 16632 16099
rect 16580 16056 16632 16065
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 3884 16031 3936 16040
rect 3884 15997 3893 16031
rect 3893 15997 3927 16031
rect 3927 15997 3936 16031
rect 3884 15988 3936 15997
rect 6000 15988 6052 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 10876 15988 10928 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 2044 15920 2096 15972
rect 7840 15963 7892 15972
rect 7840 15929 7849 15963
rect 7849 15929 7883 15963
rect 7883 15929 7892 15963
rect 7840 15920 7892 15929
rect 10140 15963 10192 15972
rect 10140 15929 10149 15963
rect 10149 15929 10183 15963
rect 10183 15929 10192 15963
rect 10140 15920 10192 15929
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 5172 15852 5224 15904
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7012 15852 7064 15904
rect 13360 15852 13412 15904
rect 14188 15920 14240 15972
rect 15752 15920 15804 15972
rect 16948 15920 17000 15972
rect 16396 15895 16448 15904
rect 16396 15861 16405 15895
rect 16405 15861 16439 15895
rect 16439 15861 16448 15895
rect 16396 15852 16448 15861
rect 16488 15895 16540 15904
rect 16488 15861 16497 15895
rect 16497 15861 16531 15895
rect 16531 15861 16540 15895
rect 17500 15895 17552 15904
rect 16488 15852 16540 15861
rect 17500 15861 17509 15895
rect 17509 15861 17543 15895
rect 17543 15861 17552 15895
rect 17500 15852 17552 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2044 15648 2096 15700
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 2320 15648 2372 15700
rect 3056 15648 3108 15700
rect 4160 15648 4212 15700
rect 5540 15648 5592 15700
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 12808 15648 12860 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 15384 15648 15436 15700
rect 5264 15580 5316 15632
rect 6460 15580 6512 15632
rect 8484 15623 8536 15632
rect 2688 15512 2740 15564
rect 4712 15512 4764 15564
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 6276 15512 6328 15564
rect 6736 15512 6788 15564
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 8484 15589 8493 15623
rect 8493 15589 8527 15623
rect 8527 15589 8536 15623
rect 8484 15580 8536 15589
rect 9036 15623 9088 15632
rect 9036 15589 9045 15623
rect 9045 15589 9079 15623
rect 9079 15589 9088 15623
rect 9036 15580 9088 15589
rect 9588 15580 9640 15632
rect 9956 15623 10008 15632
rect 9956 15589 9965 15623
rect 9965 15589 9999 15623
rect 9999 15589 10008 15623
rect 9956 15580 10008 15589
rect 9496 15512 9548 15564
rect 12072 15512 12124 15564
rect 12900 15512 12952 15564
rect 14556 15512 14608 15564
rect 2044 15444 2096 15496
rect 3240 15444 3292 15496
rect 5080 15444 5132 15496
rect 5264 15444 5316 15496
rect 6460 15444 6512 15496
rect 7196 15444 7248 15496
rect 7656 15444 7708 15496
rect 9864 15444 9916 15496
rect 11060 15444 11112 15496
rect 12532 15444 12584 15496
rect 3884 15419 3936 15428
rect 3884 15385 3893 15419
rect 3893 15385 3927 15419
rect 3927 15385 3936 15419
rect 3884 15376 3936 15385
rect 9588 15376 9640 15428
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 8024 15308 8076 15360
rect 8576 15308 8628 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 13912 15376 13964 15428
rect 16488 15648 16540 15700
rect 17776 15648 17828 15700
rect 16672 15623 16724 15632
rect 16672 15589 16681 15623
rect 16681 15589 16715 15623
rect 16715 15589 16724 15623
rect 16672 15580 16724 15589
rect 21088 15580 21140 15632
rect 15568 15512 15620 15564
rect 15936 15512 15988 15564
rect 17500 15512 17552 15564
rect 17868 15512 17920 15564
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 15568 15376 15620 15428
rect 12992 15308 13044 15360
rect 15384 15308 15436 15360
rect 16488 15308 16540 15360
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 18144 15308 18196 15317
rect 18512 15308 18564 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 3240 15147 3292 15156
rect 3240 15113 3249 15147
rect 3249 15113 3283 15147
rect 3283 15113 3292 15147
rect 3240 15104 3292 15113
rect 5448 15104 5500 15156
rect 5540 15079 5592 15088
rect 5540 15045 5549 15079
rect 5549 15045 5583 15079
rect 5583 15045 5592 15079
rect 5540 15036 5592 15045
rect 6276 15104 6328 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10140 15104 10192 15156
rect 10968 15104 11020 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 13820 15147 13872 15156
rect 12440 15104 12492 15113
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 14464 15104 14516 15156
rect 17684 15104 17736 15156
rect 17960 15104 18012 15156
rect 20904 15147 20956 15156
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 1584 14968 1636 15020
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 12532 15036 12584 15088
rect 10692 14968 10744 14977
rect 13360 14968 13412 15020
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 6920 14900 6972 14952
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 15384 14900 15436 14952
rect 17960 14900 18012 14952
rect 2228 14832 2280 14884
rect 3608 14832 3660 14884
rect 4528 14832 4580 14884
rect 7012 14832 7064 14884
rect 6460 14764 6512 14816
rect 7656 14764 7708 14816
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10968 14832 11020 14884
rect 11152 14764 11204 14816
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 12532 14764 12584 14816
rect 16304 14832 16356 14884
rect 17408 14875 17460 14884
rect 17408 14841 17417 14875
rect 17417 14841 17451 14875
rect 17451 14841 17460 14875
rect 17408 14832 17460 14841
rect 17684 14832 17736 14884
rect 15936 14764 15988 14816
rect 17132 14807 17184 14816
rect 17132 14773 17141 14807
rect 17141 14773 17175 14807
rect 17175 14773 17184 14807
rect 17132 14764 17184 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2688 14560 2740 14612
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 10692 14560 10744 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 1768 14492 1820 14544
rect 2136 14424 2188 14476
rect 2780 14424 2832 14476
rect 4160 14492 4212 14544
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 5448 14467 5500 14476
rect 5448 14433 5482 14467
rect 5482 14433 5500 14467
rect 5448 14424 5500 14433
rect 7656 14535 7708 14544
rect 7656 14501 7690 14535
rect 7690 14501 7708 14535
rect 7656 14492 7708 14501
rect 10784 14492 10836 14544
rect 11520 14492 11572 14544
rect 12992 14492 13044 14544
rect 16580 14492 16632 14544
rect 17132 14492 17184 14544
rect 2228 14356 2280 14408
rect 3700 14356 3752 14408
rect 6920 14356 6972 14408
rect 8944 14424 8996 14476
rect 9496 14467 9548 14476
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 10048 14356 10100 14408
rect 12716 14424 12768 14476
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 15384 14356 15436 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 3976 14288 4028 14340
rect 1400 14220 1452 14272
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 6368 14220 6420 14272
rect 7012 14220 7064 14272
rect 8576 14220 8628 14272
rect 12716 14288 12768 14340
rect 15844 14331 15896 14340
rect 15844 14297 15853 14331
rect 15853 14297 15887 14331
rect 15887 14297 15896 14331
rect 15844 14288 15896 14297
rect 10968 14220 11020 14272
rect 12256 14220 12308 14272
rect 12900 14220 12952 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 16856 14220 16908 14272
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 17960 14220 18012 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2320 14016 2372 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 5540 14016 5592 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 6920 14016 6972 14068
rect 7656 14016 7708 14068
rect 8484 14016 8536 14068
rect 3884 13948 3936 14000
rect 10784 14016 10836 14068
rect 12532 14016 12584 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 15476 14016 15528 14068
rect 16856 14059 16908 14068
rect 16856 14025 16865 14059
rect 16865 14025 16899 14059
rect 16899 14025 16908 14059
rect 16856 14016 16908 14025
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 19340 14016 19392 14068
rect 2596 13880 2648 13932
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 4528 13880 4580 13932
rect 4988 13880 5040 13932
rect 11152 13948 11204 14000
rect 12624 13948 12676 14000
rect 1492 13744 1544 13796
rect 4896 13812 4948 13864
rect 6184 13812 6236 13864
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 12256 13880 12308 13932
rect 12992 13880 13044 13932
rect 10140 13812 10192 13864
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 13544 13812 13596 13864
rect 15384 13812 15436 13864
rect 16488 13812 16540 13864
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24676 13855 24728 13864
rect 24676 13821 24710 13855
rect 24710 13821 24728 13855
rect 24676 13812 24728 13821
rect 6644 13744 6696 13796
rect 7380 13744 7432 13796
rect 12164 13744 12216 13796
rect 17960 13744 18012 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 4988 13719 5040 13728
rect 4988 13685 4997 13719
rect 4997 13685 5031 13719
rect 5031 13685 5040 13719
rect 4988 13676 5040 13685
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 11980 13719 12032 13728
rect 11980 13685 11989 13719
rect 11989 13685 12023 13719
rect 12023 13685 12032 13719
rect 11980 13676 12032 13685
rect 12348 13676 12400 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 6736 13472 6788 13524
rect 7012 13472 7064 13524
rect 7196 13472 7248 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9036 13472 9088 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11980 13472 12032 13524
rect 12808 13472 12860 13524
rect 13544 13472 13596 13524
rect 16396 13472 16448 13524
rect 3056 13404 3108 13456
rect 2688 13268 2740 13320
rect 2412 13243 2464 13252
rect 2412 13209 2421 13243
rect 2421 13209 2455 13243
rect 2455 13209 2464 13243
rect 2412 13200 2464 13209
rect 4804 13336 4856 13388
rect 5540 13336 5592 13388
rect 6920 13336 6972 13388
rect 12256 13404 12308 13456
rect 16580 13404 16632 13456
rect 17592 13404 17644 13456
rect 24400 13447 24452 13456
rect 24400 13413 24409 13447
rect 24409 13413 24443 13447
rect 24443 13413 24452 13447
rect 24400 13404 24452 13413
rect 9680 13336 9732 13388
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 12348 13336 12400 13388
rect 12992 13336 13044 13388
rect 15752 13336 15804 13388
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 4160 13268 4212 13320
rect 4896 13268 4948 13320
rect 6000 13268 6052 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 9404 13268 9456 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10784 13268 10836 13320
rect 16028 13311 16080 13320
rect 8392 13200 8444 13252
rect 9588 13200 9640 13252
rect 11520 13243 11572 13252
rect 11520 13209 11529 13243
rect 11529 13209 11563 13243
rect 11563 13209 11572 13243
rect 11520 13200 11572 13209
rect 12716 13200 12768 13252
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16304 13268 16356 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 4068 13132 4120 13184
rect 9220 13132 9272 13184
rect 11060 13132 11112 13184
rect 16764 13200 16816 13252
rect 13544 13132 13596 13184
rect 13912 13132 13964 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12928 1728 12980
rect 2964 12928 3016 12980
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 4896 12928 4948 12980
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8668 12928 8720 12980
rect 8852 12971 8904 12980
rect 8852 12937 8861 12971
rect 8861 12937 8895 12971
rect 8895 12937 8904 12971
rect 8852 12928 8904 12937
rect 9312 12928 9364 12980
rect 10048 12928 10100 12980
rect 11704 12928 11756 12980
rect 11980 12928 12032 12980
rect 12716 12928 12768 12980
rect 14832 12928 14884 12980
rect 15752 12971 15804 12980
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 16028 12928 16080 12980
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 1492 12724 1544 12776
rect 2044 12656 2096 12708
rect 3148 12656 3200 12708
rect 2596 12588 2648 12640
rect 4528 12860 4580 12912
rect 4988 12792 5040 12844
rect 5264 12724 5316 12776
rect 4804 12656 4856 12708
rect 4160 12588 4212 12640
rect 6644 12860 6696 12912
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 10324 12860 10376 12869
rect 6920 12724 6972 12776
rect 7932 12656 7984 12708
rect 8668 12792 8720 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 10048 12792 10100 12844
rect 12808 12792 12860 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 16396 12860 16448 12912
rect 16488 12860 16540 12912
rect 15568 12792 15620 12801
rect 9220 12767 9272 12776
rect 9220 12733 9254 12767
rect 9254 12733 9272 12767
rect 9220 12724 9272 12733
rect 14556 12724 14608 12776
rect 14740 12724 14792 12776
rect 17132 12724 17184 12776
rect 14096 12656 14148 12708
rect 6368 12588 6420 12640
rect 7012 12588 7064 12640
rect 8944 12588 8996 12640
rect 10784 12588 10836 12640
rect 11060 12588 11112 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2964 12384 3016 12436
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 5540 12384 5592 12436
rect 7012 12384 7064 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 13544 12427 13596 12436
rect 4528 12316 4580 12368
rect 6184 12359 6236 12368
rect 1492 12248 1544 12300
rect 1860 12248 1912 12300
rect 2596 12248 2648 12300
rect 3976 12248 4028 12300
rect 6184 12325 6193 12359
rect 6193 12325 6227 12359
rect 6227 12325 6236 12359
rect 6184 12316 6236 12325
rect 7748 12316 7800 12368
rect 11520 12316 11572 12368
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 14648 12384 14700 12436
rect 16304 12427 16356 12436
rect 16304 12393 16313 12427
rect 16313 12393 16347 12427
rect 16347 12393 16356 12427
rect 16304 12384 16356 12393
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 18604 12384 18656 12436
rect 12992 12316 13044 12368
rect 6828 12248 6880 12300
rect 8208 12248 8260 12300
rect 10692 12248 10744 12300
rect 16672 12316 16724 12368
rect 4068 12180 4120 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 7380 12223 7432 12232
rect 6276 12180 6328 12189
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 5540 12112 5592 12164
rect 10508 12112 10560 12164
rect 2872 12044 2924 12096
rect 4804 12044 4856 12096
rect 9220 12044 9272 12096
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9680 12044 9732 12096
rect 10600 12044 10652 12096
rect 14556 12180 14608 12232
rect 12256 12044 12308 12096
rect 13544 12112 13596 12164
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 17868 12180 17920 12232
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 14280 12087 14332 12096
rect 13912 12044 13964 12053
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 14740 12044 14792 12096
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2780 11840 2832 11892
rect 4712 11840 4764 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 6828 11840 6880 11892
rect 7564 11840 7616 11892
rect 7840 11840 7892 11892
rect 10140 11840 10192 11892
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 14648 11840 14700 11892
rect 16028 11840 16080 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 17500 11840 17552 11892
rect 3148 11815 3200 11824
rect 3148 11781 3157 11815
rect 3157 11781 3191 11815
rect 3191 11781 3200 11815
rect 3148 11772 3200 11781
rect 3976 11815 4028 11824
rect 3976 11781 3985 11815
rect 3985 11781 4019 11815
rect 4019 11781 4028 11815
rect 3976 11772 4028 11781
rect 8208 11815 8260 11824
rect 8208 11781 8217 11815
rect 8217 11781 8251 11815
rect 8251 11781 8260 11815
rect 8208 11772 8260 11781
rect 10048 11772 10100 11824
rect 10324 11772 10376 11824
rect 13912 11772 13964 11824
rect 1492 11704 1544 11756
rect 3884 11704 3936 11756
rect 4804 11704 4856 11756
rect 9404 11704 9456 11756
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 7380 11636 7432 11688
rect 8760 11636 8812 11688
rect 10508 11704 10560 11756
rect 10140 11636 10192 11688
rect 10876 11636 10928 11688
rect 11796 11636 11848 11688
rect 2320 11568 2372 11620
rect 7472 11568 7524 11620
rect 9404 11568 9456 11620
rect 9772 11611 9824 11620
rect 9772 11577 9781 11611
rect 9781 11577 9815 11611
rect 9815 11577 9824 11611
rect 9772 11568 9824 11577
rect 10048 11568 10100 11620
rect 12348 11636 12400 11688
rect 12992 11679 13044 11688
rect 12992 11645 13026 11679
rect 13026 11645 13044 11679
rect 12992 11636 13044 11645
rect 15200 11611 15252 11620
rect 15200 11577 15209 11611
rect 15209 11577 15243 11611
rect 15243 11577 15252 11611
rect 15200 11568 15252 11577
rect 15476 11568 15528 11620
rect 3056 11500 3108 11552
rect 4252 11500 4304 11552
rect 6092 11500 6144 11552
rect 10140 11500 10192 11552
rect 10692 11500 10744 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11520 11500 11572 11552
rect 15108 11500 15160 11552
rect 16672 11500 16724 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 6000 11296 6052 11348
rect 8208 11296 8260 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 11152 11296 11204 11348
rect 13452 11296 13504 11348
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 17316 11296 17368 11348
rect 1584 11228 1636 11280
rect 2504 11228 2556 11280
rect 3976 11228 4028 11280
rect 4436 11271 4488 11280
rect 4436 11237 4445 11271
rect 4445 11237 4479 11271
rect 4479 11237 4488 11271
rect 4436 11228 4488 11237
rect 4712 11228 4764 11280
rect 8484 11271 8536 11280
rect 8484 11237 8493 11271
rect 8493 11237 8527 11271
rect 8527 11237 8536 11271
rect 8484 11228 8536 11237
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 3792 11160 3844 11212
rect 4252 11160 4304 11212
rect 5540 11160 5592 11212
rect 6368 11160 6420 11212
rect 7748 11160 7800 11212
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 2412 11024 2464 11076
rect 2504 10956 2556 11008
rect 2688 11024 2740 11076
rect 4804 11092 4856 11144
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 4344 10956 4396 11008
rect 7380 11024 7432 11076
rect 7840 11067 7892 11076
rect 6000 10956 6052 11008
rect 7472 10956 7524 11008
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 9588 11160 9640 11212
rect 10324 11160 10376 11212
rect 9864 11092 9916 11144
rect 11520 11092 11572 11144
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 9404 10956 9456 11008
rect 10968 11024 11020 11076
rect 13268 11228 13320 11280
rect 14280 11228 14332 11280
rect 16580 11228 16632 11280
rect 16764 11271 16816 11280
rect 16764 11237 16773 11271
rect 16773 11237 16807 11271
rect 16807 11237 16816 11271
rect 16764 11228 16816 11237
rect 14004 11160 14056 11212
rect 15384 11160 15436 11212
rect 15568 11160 15620 11212
rect 17592 11160 17644 11212
rect 13360 11092 13412 11144
rect 13544 11092 13596 11144
rect 14096 11092 14148 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 16212 11024 16264 11076
rect 11152 10956 11204 11008
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 14004 10956 14056 11008
rect 14280 10956 14332 11008
rect 16120 10956 16172 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1400 10795 1452 10804
rect 1400 10761 1409 10795
rect 1409 10761 1443 10795
rect 1443 10761 1452 10795
rect 1400 10752 1452 10761
rect 2780 10752 2832 10804
rect 2964 10752 3016 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 6276 10752 6328 10804
rect 7380 10752 7432 10804
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 12072 10752 12124 10804
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 5448 10684 5500 10736
rect 7748 10684 7800 10736
rect 9956 10684 10008 10736
rect 12808 10684 12860 10736
rect 17316 10752 17368 10804
rect 2780 10548 2832 10600
rect 6092 10616 6144 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 9772 10616 9824 10668
rect 11428 10659 11480 10668
rect 4344 10548 4396 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 8576 10548 8628 10600
rect 11428 10625 11437 10659
rect 11437 10625 11471 10659
rect 11471 10625 11480 10659
rect 11428 10616 11480 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17500 10616 17552 10668
rect 12532 10548 12584 10600
rect 14372 10548 14424 10600
rect 15200 10548 15252 10600
rect 15384 10548 15436 10600
rect 2688 10480 2740 10532
rect 12072 10480 12124 10532
rect 13820 10480 13872 10532
rect 15016 10523 15068 10532
rect 15016 10489 15025 10523
rect 15025 10489 15059 10523
rect 15059 10489 15068 10523
rect 15016 10480 15068 10489
rect 16120 10480 16172 10532
rect 2228 10412 2280 10464
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 4620 10412 4672 10464
rect 4712 10412 4764 10464
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 9864 10412 9916 10464
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 14096 10412 14148 10464
rect 14280 10412 14332 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 17592 10455 17644 10464
rect 17592 10421 17601 10455
rect 17601 10421 17635 10455
rect 17635 10421 17644 10455
rect 17592 10412 17644 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2688 10208 2740 10260
rect 3516 10208 3568 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 8576 10208 8628 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 11428 10251 11480 10260
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 11796 10251 11848 10260
rect 11796 10217 11805 10251
rect 11805 10217 11839 10251
rect 11839 10217 11848 10251
rect 11796 10208 11848 10217
rect 15568 10208 15620 10260
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 17868 10208 17920 10260
rect 2228 10140 2280 10192
rect 3884 10183 3936 10192
rect 3884 10149 3893 10183
rect 3893 10149 3927 10183
rect 3927 10149 3936 10183
rect 3884 10140 3936 10149
rect 4528 10140 4580 10192
rect 4988 10140 5040 10192
rect 4068 10072 4120 10124
rect 5632 10115 5684 10124
rect 5632 10081 5641 10115
rect 5641 10081 5675 10115
rect 5675 10081 5684 10115
rect 5632 10072 5684 10081
rect 6000 10072 6052 10124
rect 6828 10140 6880 10192
rect 8024 10140 8076 10192
rect 13728 10140 13780 10192
rect 14096 10140 14148 10192
rect 14648 10140 14700 10192
rect 6368 10115 6420 10124
rect 6368 10081 6402 10115
rect 6402 10081 6420 10115
rect 6368 10072 6420 10081
rect 7748 10072 7800 10124
rect 8484 10072 8536 10124
rect 9772 10072 9824 10124
rect 9956 10115 10008 10124
rect 9956 10081 9990 10115
rect 9990 10081 10008 10115
rect 9956 10072 10008 10081
rect 11980 10072 12032 10124
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 2136 10004 2188 10056
rect 3148 10004 3200 10056
rect 4436 10004 4488 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 12348 10072 12400 10124
rect 12992 10072 13044 10124
rect 9680 10004 9732 10013
rect 5264 9868 5316 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11152 9868 11204 9920
rect 15384 10004 15436 10056
rect 16028 10140 16080 10192
rect 15568 10072 15620 10124
rect 16488 10072 16540 10124
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 17592 9936 17644 9988
rect 13452 9868 13504 9920
rect 13820 9868 13872 9920
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 6736 9664 6788 9716
rect 7196 9664 7248 9716
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 14556 9664 14608 9716
rect 16948 9664 17000 9716
rect 2688 9639 2740 9648
rect 2688 9605 2697 9639
rect 2697 9605 2731 9639
rect 2731 9605 2740 9639
rect 2688 9596 2740 9605
rect 4160 9596 4212 9648
rect 6552 9596 6604 9648
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 4620 9528 4672 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2780 9503 2832 9512
rect 2780 9469 2796 9503
rect 2796 9469 2830 9503
rect 2830 9469 2832 9503
rect 3056 9503 3108 9512
rect 2780 9460 2832 9469
rect 3056 9469 3090 9503
rect 3090 9469 3108 9503
rect 3056 9460 3108 9469
rect 3424 9460 3476 9512
rect 6920 9460 6972 9512
rect 7196 9460 7248 9512
rect 11704 9596 11756 9648
rect 12256 9639 12308 9648
rect 12256 9605 12265 9639
rect 12265 9605 12299 9639
rect 12299 9605 12308 9639
rect 12256 9596 12308 9605
rect 3608 9392 3660 9444
rect 1676 9324 1728 9376
rect 3148 9324 3200 9376
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 4528 9324 4580 9376
rect 5264 9324 5316 9376
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 6368 9392 6420 9444
rect 7104 9392 7156 9444
rect 9036 9460 9088 9512
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 12532 9528 12584 9580
rect 15476 9596 15528 9648
rect 10968 9460 11020 9512
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 16580 9596 16632 9648
rect 18052 9596 18104 9648
rect 18512 9664 18564 9716
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 18236 9528 18288 9580
rect 5448 9324 5500 9333
rect 7012 9324 7064 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 8024 9324 8076 9376
rect 9936 9324 9988 9376
rect 11060 9324 11112 9376
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 16672 9324 16724 9376
rect 17500 9324 17552 9376
rect 17868 9324 17920 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1952 9120 2004 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 1676 9095 1728 9104
rect 1676 9061 1710 9095
rect 1710 9061 1728 9095
rect 1676 9052 1728 9061
rect 3056 9052 3108 9104
rect 4620 9120 4672 9172
rect 4896 9052 4948 9104
rect 7656 9120 7708 9172
rect 8024 9120 8076 9172
rect 7196 9052 7248 9104
rect 9772 9120 9824 9172
rect 12440 9120 12492 9172
rect 12900 9163 12952 9172
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 16304 9120 16356 9172
rect 16948 9120 17000 9172
rect 1492 8984 1544 9036
rect 2780 8984 2832 9036
rect 4804 8984 4856 9036
rect 5908 8984 5960 9036
rect 6460 8984 6512 9036
rect 7012 8984 7064 9036
rect 8024 8984 8076 9036
rect 10416 9052 10468 9104
rect 11152 9052 11204 9104
rect 13544 9052 13596 9104
rect 14188 9095 14240 9104
rect 14188 9061 14197 9095
rect 14197 9061 14231 9095
rect 14231 9061 14240 9095
rect 14188 9052 14240 9061
rect 10784 9027 10836 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 6920 8916 6972 8968
rect 7932 8916 7984 8968
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 9128 8916 9180 8968
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 12440 8984 12492 9036
rect 12992 8984 13044 9036
rect 15292 8984 15344 9036
rect 16028 8984 16080 9036
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 13452 8916 13504 8968
rect 15384 8916 15436 8968
rect 15936 8959 15988 8968
rect 10324 8848 10376 8900
rect 11980 8848 12032 8900
rect 14280 8848 14332 8900
rect 5448 8780 5500 8832
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 9956 8780 10008 8832
rect 10232 8780 10284 8832
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 11796 8780 11848 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 15844 8780 15896 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 17500 8780 17552 8832
rect 17868 8780 17920 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1860 8576 1912 8628
rect 4896 8576 4948 8628
rect 6184 8576 6236 8628
rect 8024 8619 8076 8628
rect 4068 8551 4120 8560
rect 4068 8517 4077 8551
rect 4077 8517 4111 8551
rect 4111 8517 4120 8551
rect 4068 8508 4120 8517
rect 1492 8440 1544 8492
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9036 8576 9088 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 11796 8576 11848 8628
rect 12900 8576 12952 8628
rect 14556 8576 14608 8628
rect 16396 8576 16448 8628
rect 9312 8508 9364 8560
rect 4620 8440 4672 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8024 8440 8076 8492
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 1952 8372 2004 8424
rect 4436 8415 4488 8424
rect 2780 8304 2832 8356
rect 4068 8304 4120 8356
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 11244 8440 11296 8492
rect 11704 8440 11756 8492
rect 13268 8508 13320 8560
rect 15384 8508 15436 8560
rect 16028 8508 16080 8560
rect 14188 8483 14240 8492
rect 4804 8304 4856 8356
rect 5448 8304 5500 8356
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 4252 8236 4304 8288
rect 6552 8236 6604 8288
rect 6828 8279 6880 8288
rect 6828 8245 6837 8279
rect 6837 8245 6871 8279
rect 6871 8245 6880 8279
rect 6828 8236 6880 8245
rect 9128 8236 9180 8288
rect 9496 8236 9548 8288
rect 9680 8304 9732 8356
rect 10968 8304 11020 8356
rect 11336 8304 11388 8356
rect 12164 8347 12216 8356
rect 12164 8313 12173 8347
rect 12173 8313 12207 8347
rect 12207 8313 12216 8347
rect 12164 8304 12216 8313
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 16396 8372 16448 8424
rect 17500 8415 17552 8424
rect 17500 8381 17509 8415
rect 17509 8381 17543 8415
rect 17543 8381 17552 8415
rect 17500 8372 17552 8381
rect 13544 8304 13596 8356
rect 14556 8304 14608 8356
rect 15292 8304 15344 8356
rect 16488 8304 16540 8356
rect 17868 8347 17920 8356
rect 17868 8313 17877 8347
rect 17877 8313 17911 8347
rect 17911 8313 17920 8347
rect 17868 8304 17920 8313
rect 12072 8236 12124 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 16396 8279 16448 8288
rect 16396 8245 16405 8279
rect 16405 8245 16439 8279
rect 16439 8245 16448 8279
rect 16396 8236 16448 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 2688 8032 2740 8084
rect 3148 8032 3200 8084
rect 4620 8032 4672 8084
rect 5540 8075 5592 8084
rect 2872 7964 2924 8016
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6828 8032 6880 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 4988 7964 5040 8016
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 6184 7896 6236 7948
rect 6552 7964 6604 8016
rect 7380 8032 7432 8084
rect 7932 8032 7984 8084
rect 8576 8032 8628 8084
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 10140 8032 10192 8084
rect 12164 8032 12216 8084
rect 12900 8032 12952 8084
rect 13636 8032 13688 8084
rect 13728 8032 13780 8084
rect 13912 8032 13964 8084
rect 14372 8032 14424 8084
rect 15292 8075 15344 8084
rect 15292 8041 15301 8075
rect 15301 8041 15335 8075
rect 15335 8041 15344 8075
rect 15292 8032 15344 8041
rect 15936 8032 15988 8084
rect 8760 7964 8812 8016
rect 16672 7964 16724 8016
rect 18972 8007 19024 8016
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 10784 7896 10836 7948
rect 10968 7939 11020 7948
rect 10968 7905 10991 7939
rect 10991 7905 11020 7939
rect 10968 7896 11020 7905
rect 12440 7896 12492 7948
rect 13360 7896 13412 7948
rect 13636 7896 13688 7948
rect 13820 7896 13872 7948
rect 18972 7973 18981 8007
rect 18981 7973 19015 8007
rect 19015 7973 19024 8007
rect 18972 7964 19024 7973
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 3148 7828 3200 7880
rect 5172 7828 5224 7880
rect 7196 7828 7248 7880
rect 13452 7828 13504 7880
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 6092 7760 6144 7812
rect 7380 7760 7432 7812
rect 11980 7760 12032 7812
rect 14648 7760 14700 7812
rect 17776 7828 17828 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5448 7692 5500 7744
rect 6460 7692 6512 7744
rect 6736 7735 6788 7744
rect 6736 7701 6745 7735
rect 6745 7701 6779 7735
rect 6779 7701 6788 7735
rect 6736 7692 6788 7701
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 13452 7692 13504 7744
rect 13912 7692 13964 7744
rect 14096 7692 14148 7744
rect 14188 7692 14240 7744
rect 17960 7692 18012 7744
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 1768 7420 1820 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 5356 7420 5408 7472
rect 5632 7420 5684 7472
rect 6552 7488 6604 7540
rect 7104 7488 7156 7540
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 11612 7488 11664 7540
rect 12256 7488 12308 7540
rect 13360 7488 13412 7540
rect 16396 7488 16448 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 18604 7488 18656 7540
rect 18972 7488 19024 7540
rect 10692 7420 10744 7472
rect 15476 7463 15528 7472
rect 15476 7429 15485 7463
rect 15485 7429 15519 7463
rect 15519 7429 15528 7463
rect 15476 7420 15528 7429
rect 3792 7352 3844 7404
rect 1676 7284 1728 7336
rect 2780 7284 2832 7336
rect 3700 7284 3752 7336
rect 6000 7352 6052 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 8576 7352 8628 7404
rect 11336 7395 11388 7404
rect 7288 7284 7340 7336
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 9496 7284 9548 7336
rect 9680 7284 9732 7336
rect 11980 7284 12032 7336
rect 3884 7216 3936 7268
rect 6276 7216 6328 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 4896 7148 4948 7200
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 6920 7148 6972 7200
rect 8944 7259 8996 7268
rect 8944 7225 8978 7259
rect 8978 7225 8996 7259
rect 8944 7216 8996 7225
rect 9956 7216 10008 7268
rect 11336 7216 11388 7268
rect 12072 7216 12124 7268
rect 15752 7352 15804 7404
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 17960 7352 18012 7404
rect 16396 7284 16448 7336
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 18052 7284 18104 7336
rect 18236 7284 18288 7336
rect 18512 7284 18564 7336
rect 13452 7216 13504 7268
rect 10140 7148 10192 7200
rect 11244 7148 11296 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 15200 7148 15252 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 18604 7148 18656 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3056 6944 3108 6996
rect 5172 6944 5224 6996
rect 6092 6944 6144 6996
rect 7196 6944 7248 6996
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 13544 6944 13596 6996
rect 13728 6987 13780 6996
rect 13728 6953 13737 6987
rect 13737 6953 13771 6987
rect 13771 6953 13780 6987
rect 13728 6944 13780 6953
rect 18880 6944 18932 6996
rect 2044 6876 2096 6928
rect 3792 6876 3844 6928
rect 1400 6808 1452 6860
rect 2872 6808 2924 6860
rect 4988 6876 5040 6928
rect 7380 6876 7432 6928
rect 12532 6876 12584 6928
rect 16120 6876 16172 6928
rect 4896 6808 4948 6860
rect 6000 6808 6052 6860
rect 8576 6808 8628 6860
rect 9772 6808 9824 6860
rect 5908 6672 5960 6724
rect 6276 6672 6328 6724
rect 2320 6604 2372 6656
rect 5540 6604 5592 6656
rect 7288 6604 7340 6656
rect 8024 6604 8076 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 12072 6783 12124 6792
rect 11060 6715 11112 6724
rect 11060 6681 11069 6715
rect 11069 6681 11103 6715
rect 11103 6681 11112 6715
rect 11060 6672 11112 6681
rect 9036 6604 9088 6613
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 14464 6740 14516 6792
rect 14740 6740 14792 6792
rect 15292 6740 15344 6792
rect 19432 6808 19484 6860
rect 19156 6740 19208 6792
rect 15200 6672 15252 6724
rect 19524 6715 19576 6724
rect 19524 6681 19533 6715
rect 19533 6681 19567 6715
rect 19567 6681 19576 6715
rect 19524 6672 19576 6681
rect 20444 6672 20496 6724
rect 11520 6604 11572 6656
rect 11612 6604 11664 6656
rect 11980 6604 12032 6656
rect 13636 6604 13688 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 15568 6604 15620 6656
rect 16304 6604 16356 6656
rect 16672 6604 16724 6656
rect 18512 6604 18564 6656
rect 20260 6604 20312 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3976 6400 4028 6452
rect 4896 6400 4948 6452
rect 6092 6400 6144 6452
rect 1400 6264 1452 6316
rect 2780 6264 2832 6316
rect 6000 6264 6052 6316
rect 1768 6171 1820 6180
rect 1768 6137 1802 6171
rect 1802 6137 1820 6171
rect 1768 6128 1820 6137
rect 2044 6060 2096 6112
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 4160 6060 4212 6112
rect 7380 6400 7432 6452
rect 7656 6400 7708 6452
rect 11704 6400 11756 6452
rect 15476 6400 15528 6452
rect 16764 6400 16816 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 9772 6332 9824 6384
rect 8576 6264 8628 6316
rect 18604 6307 18656 6316
rect 8024 6128 8076 6180
rect 10140 6128 10192 6180
rect 12072 6196 12124 6248
rect 13268 6196 13320 6248
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 5632 6103 5684 6112
rect 4988 6060 5040 6069
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7380 6060 7432 6112
rect 10968 6060 11020 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11428 6103 11480 6112
rect 11428 6069 11437 6103
rect 11437 6069 11471 6103
rect 11471 6069 11480 6103
rect 11428 6060 11480 6069
rect 12808 6060 12860 6112
rect 14188 6128 14240 6180
rect 15292 6128 15344 6180
rect 16212 6196 16264 6248
rect 17868 6196 17920 6248
rect 16028 6128 16080 6180
rect 17960 6128 18012 6180
rect 19156 6128 19208 6180
rect 20628 6128 20680 6180
rect 13544 6060 13596 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 15476 6060 15528 6112
rect 15936 6060 15988 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 20720 6060 20772 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 4068 5856 4120 5908
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 9036 5856 9088 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 3792 5788 3844 5840
rect 4436 5788 4488 5840
rect 5264 5788 5316 5840
rect 6092 5788 6144 5840
rect 10692 5856 10744 5908
rect 11980 5856 12032 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 14740 5856 14792 5908
rect 11060 5788 11112 5840
rect 11796 5788 11848 5840
rect 15568 5856 15620 5908
rect 15936 5856 15988 5908
rect 16488 5856 16540 5908
rect 16764 5899 16816 5908
rect 16764 5865 16773 5899
rect 16773 5865 16807 5899
rect 16807 5865 16816 5899
rect 16764 5856 16816 5865
rect 19340 5899 19392 5908
rect 19340 5865 19349 5899
rect 19349 5865 19383 5899
rect 19383 5865 19392 5899
rect 19340 5856 19392 5865
rect 18236 5788 18288 5840
rect 18696 5831 18748 5840
rect 18696 5797 18705 5831
rect 18705 5797 18739 5831
rect 18739 5797 18748 5831
rect 18696 5788 18748 5797
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 5080 5720 5132 5772
rect 6920 5720 6972 5772
rect 11336 5720 11388 5772
rect 13360 5763 13412 5772
rect 13360 5729 13369 5763
rect 13369 5729 13403 5763
rect 13403 5729 13412 5763
rect 13360 5720 13412 5729
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 7012 5652 7064 5704
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 9772 5652 9824 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 12348 5652 12400 5704
rect 12808 5652 12860 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14096 5652 14148 5704
rect 15844 5652 15896 5704
rect 16672 5652 16724 5704
rect 17316 5652 17368 5704
rect 1768 5584 1820 5636
rect 3056 5584 3108 5636
rect 9680 5627 9732 5636
rect 9680 5593 9689 5627
rect 9689 5593 9723 5627
rect 9723 5593 9732 5627
rect 9680 5584 9732 5593
rect 12900 5627 12952 5636
rect 12900 5593 12909 5627
rect 12909 5593 12943 5627
rect 12943 5593 12952 5627
rect 12900 5584 12952 5593
rect 13636 5584 13688 5636
rect 16028 5584 16080 5636
rect 16580 5584 16632 5636
rect 17592 5584 17644 5636
rect 18604 5652 18656 5704
rect 19156 5652 19208 5704
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 23480 5652 23532 5704
rect 18880 5627 18932 5636
rect 18880 5593 18889 5627
rect 18889 5593 18923 5627
rect 18923 5593 18932 5627
rect 18880 5584 18932 5593
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 10692 5516 10744 5568
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 12440 5516 12492 5525
rect 13820 5516 13872 5568
rect 14188 5516 14240 5568
rect 16304 5516 16356 5568
rect 19984 5559 20036 5568
rect 19984 5525 19993 5559
rect 19993 5525 20027 5559
rect 20027 5525 20036 5559
rect 19984 5516 20036 5525
rect 20444 5516 20496 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2596 5312 2648 5364
rect 5264 5355 5316 5364
rect 5264 5321 5273 5355
rect 5273 5321 5307 5355
rect 5307 5321 5316 5355
rect 5264 5312 5316 5321
rect 5356 5312 5408 5364
rect 6736 5312 6788 5364
rect 8944 5312 8996 5364
rect 2780 5244 2832 5296
rect 6184 5287 6236 5296
rect 6184 5253 6193 5287
rect 6193 5253 6227 5287
rect 6227 5253 6236 5287
rect 6184 5244 6236 5253
rect 9588 5312 9640 5364
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12072 5312 12124 5364
rect 12348 5312 12400 5364
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 13360 5312 13412 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 15936 5312 15988 5364
rect 17960 5312 18012 5364
rect 19248 5312 19300 5364
rect 19340 5312 19392 5364
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 4436 5176 4488 5228
rect 9312 5176 9364 5228
rect 10692 5176 10744 5228
rect 3976 5040 4028 5092
rect 1584 4972 1636 5024
rect 3792 5015 3844 5024
rect 3792 4981 3801 5015
rect 3801 4981 3835 5015
rect 3835 4981 3844 5015
rect 8576 5108 8628 5160
rect 9496 5108 9548 5160
rect 10600 5108 10652 5160
rect 6092 5040 6144 5092
rect 6552 5083 6604 5092
rect 6552 5049 6561 5083
rect 6561 5049 6595 5083
rect 6595 5049 6604 5083
rect 6552 5040 6604 5049
rect 4436 5015 4488 5024
rect 3792 4972 3844 4981
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 9404 4972 9456 5024
rect 10968 4972 11020 5024
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 12440 5176 12492 5228
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 14004 5176 14056 5228
rect 14924 5176 14976 5228
rect 15384 5176 15436 5228
rect 16488 5176 16540 5228
rect 17592 5176 17644 5228
rect 19340 5176 19392 5228
rect 11428 5108 11480 5160
rect 13728 5108 13780 5160
rect 12532 4972 12584 5024
rect 12716 4972 12768 5024
rect 13360 4972 13412 5024
rect 14096 5108 14148 5160
rect 14832 5151 14884 5160
rect 14832 5117 14841 5151
rect 14841 5117 14875 5151
rect 14875 5117 14884 5151
rect 14832 5108 14884 5117
rect 18236 5108 18288 5160
rect 18696 5108 18748 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 23480 5108 23532 5160
rect 15568 5040 15620 5092
rect 16580 5040 16632 5092
rect 20536 5083 20588 5092
rect 20536 5049 20545 5083
rect 20545 5049 20579 5083
rect 20579 5049 20588 5083
rect 20536 5040 20588 5049
rect 15384 4972 15436 5024
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 17684 5015 17736 5024
rect 17684 4981 17693 5015
rect 17693 4981 17727 5015
rect 17727 4981 17736 5015
rect 17684 4972 17736 4981
rect 25320 4972 25372 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1860 4811 1912 4820
rect 1860 4777 1869 4811
rect 1869 4777 1903 4811
rect 1903 4777 1912 4811
rect 1860 4768 1912 4777
rect 2228 4768 2280 4820
rect 2688 4768 2740 4820
rect 2780 4768 2832 4820
rect 5540 4768 5592 4820
rect 3056 4700 3108 4752
rect 4344 4743 4396 4752
rect 4344 4709 4353 4743
rect 4353 4709 4387 4743
rect 4387 4709 4396 4743
rect 4344 4700 4396 4709
rect 6000 4768 6052 4820
rect 6828 4768 6880 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7564 4768 7616 4820
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 9588 4768 9640 4820
rect 9864 4768 9916 4820
rect 11152 4768 11204 4820
rect 11428 4811 11480 4820
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 12164 4768 12216 4820
rect 13544 4768 13596 4820
rect 13728 4768 13780 4820
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14740 4768 14792 4820
rect 15292 4768 15344 4820
rect 16120 4768 16172 4820
rect 16396 4768 16448 4820
rect 17592 4768 17644 4820
rect 17868 4768 17920 4820
rect 19156 4811 19208 4820
rect 19156 4777 19165 4811
rect 19165 4777 19199 4811
rect 19199 4777 19208 4811
rect 19156 4768 19208 4777
rect 20076 4811 20128 4820
rect 20076 4777 20085 4811
rect 20085 4777 20119 4811
rect 20119 4777 20128 4811
rect 20076 4768 20128 4777
rect 22100 4811 22152 4820
rect 22100 4777 22109 4811
rect 22109 4777 22143 4811
rect 22143 4777 22152 4811
rect 22100 4768 22152 4777
rect 22560 4768 22612 4820
rect 6184 4700 6236 4752
rect 6920 4743 6972 4752
rect 6920 4709 6929 4743
rect 6929 4709 6963 4743
rect 6963 4709 6972 4743
rect 6920 4700 6972 4709
rect 9956 4700 10008 4752
rect 10140 4700 10192 4752
rect 11336 4743 11388 4752
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 11704 4700 11756 4752
rect 1492 4632 1544 4684
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 4068 4675 4120 4684
rect 4068 4641 4087 4675
rect 4087 4641 4120 4675
rect 4068 4632 4120 4641
rect 7840 4632 7892 4684
rect 8300 4632 8352 4684
rect 2320 4564 2372 4616
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 9496 4564 9548 4616
rect 9956 4564 10008 4616
rect 5540 4496 5592 4548
rect 9404 4496 9456 4548
rect 10692 4564 10744 4616
rect 14924 4632 14976 4684
rect 16120 4632 16172 4684
rect 17960 4632 18012 4684
rect 11796 4496 11848 4548
rect 13820 4564 13872 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 18236 4607 18288 4616
rect 14188 4496 14240 4548
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 19432 4700 19484 4752
rect 19524 4632 19576 4684
rect 20536 4632 20588 4684
rect 20996 4632 21048 4684
rect 22100 4632 22152 4684
rect 20076 4564 20128 4616
rect 20720 4496 20772 4548
rect 2136 4428 2188 4480
rect 3700 4471 3752 4480
rect 3700 4437 3709 4471
rect 3709 4437 3743 4471
rect 3743 4437 3752 4471
rect 3700 4428 3752 4437
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 6460 4471 6512 4480
rect 6460 4437 6469 4471
rect 6469 4437 6503 4471
rect 6503 4437 6512 4471
rect 6460 4428 6512 4437
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 12900 4428 12952 4480
rect 14372 4428 14424 4480
rect 14740 4428 14792 4480
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 21640 4428 21692 4480
rect 21824 4471 21876 4480
rect 21824 4437 21833 4471
rect 21833 4437 21867 4471
rect 21867 4437 21876 4471
rect 21824 4428 21876 4437
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2228 4224 2280 4276
rect 1400 4088 1452 4140
rect 1768 4088 1820 4140
rect 3792 4224 3844 4276
rect 7288 4224 7340 4276
rect 7932 4224 7984 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 14004 4267 14056 4276
rect 14004 4233 14013 4267
rect 14013 4233 14047 4267
rect 14047 4233 14056 4267
rect 14004 4224 14056 4233
rect 19340 4224 19392 4276
rect 19524 4224 19576 4276
rect 20996 4267 21048 4276
rect 20996 4233 21005 4267
rect 21005 4233 21039 4267
rect 21039 4233 21048 4267
rect 20996 4224 21048 4233
rect 3332 4199 3384 4208
rect 3332 4165 3341 4199
rect 3341 4165 3375 4199
rect 3375 4165 3384 4199
rect 3332 4156 3384 4165
rect 6092 4156 6144 4208
rect 5540 4088 5592 4140
rect 7564 4156 7616 4208
rect 7656 4156 7708 4208
rect 8024 4088 8076 4140
rect 8300 4199 8352 4208
rect 8300 4165 8309 4199
rect 8309 4165 8343 4199
rect 8343 4165 8352 4199
rect 8300 4156 8352 4165
rect 9036 4156 9088 4208
rect 9128 4156 9180 4208
rect 9772 4088 9824 4140
rect 11704 4156 11756 4208
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 12900 4088 12952 4140
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 3240 3952 3292 4004
rect 2320 3884 2372 3936
rect 3792 3884 3844 3936
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4896 3884 4948 3936
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 5356 4020 5408 4072
rect 5724 3952 5776 4004
rect 6460 3952 6512 4004
rect 8392 4020 8444 4072
rect 9588 4020 9640 4072
rect 11244 4020 11296 4072
rect 13636 4020 13688 4072
rect 14188 4020 14240 4072
rect 15292 4020 15344 4072
rect 16580 4020 16632 4072
rect 18236 4156 18288 4208
rect 20168 4156 20220 4208
rect 6092 3884 6144 3936
rect 6276 3884 6328 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 8300 3952 8352 4004
rect 8484 3952 8536 4004
rect 7288 3884 7340 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9680 3884 9732 3936
rect 9956 3884 10008 3936
rect 10876 3884 10928 3936
rect 11520 3884 11572 3936
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 12716 3952 12768 4004
rect 13820 3952 13872 4004
rect 14372 3952 14424 4004
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 13544 3884 13596 3936
rect 16764 3995 16816 4004
rect 16120 3884 16172 3936
rect 16764 3961 16773 3995
rect 16773 3961 16807 3995
rect 16807 3961 16816 3995
rect 16764 3952 16816 3961
rect 19248 4088 19300 4140
rect 18052 4020 18104 4072
rect 18788 4020 18840 4072
rect 19340 4020 19392 4072
rect 19984 4063 20036 4072
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 21180 4063 21232 4072
rect 21180 4029 21189 4063
rect 21189 4029 21223 4063
rect 21223 4029 21232 4063
rect 21180 4020 21232 4029
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 18144 3952 18196 4004
rect 18328 3884 18380 3936
rect 20352 3952 20404 4004
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 22376 3952 22428 4004
rect 22100 3927 22152 3936
rect 22100 3893 22109 3927
rect 22109 3893 22143 3927
rect 22143 3893 22152 3927
rect 22468 3927 22520 3936
rect 22100 3884 22152 3893
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 22468 3884 22520 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 2780 3680 2832 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 6000 3680 6052 3732
rect 6184 3723 6236 3732
rect 6184 3689 6193 3723
rect 6193 3689 6227 3723
rect 6227 3689 6236 3723
rect 6184 3680 6236 3689
rect 7748 3680 7800 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 11336 3680 11388 3732
rect 4068 3612 4120 3664
rect 5540 3612 5592 3664
rect 7840 3612 7892 3664
rect 12440 3680 12492 3732
rect 12532 3680 12584 3732
rect 13636 3680 13688 3732
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 16028 3723 16080 3732
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 17132 3723 17184 3732
rect 17132 3689 17141 3723
rect 17141 3689 17175 3723
rect 17175 3689 17184 3723
rect 17132 3680 17184 3689
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 17960 3680 18012 3732
rect 21456 3723 21508 3732
rect 21456 3689 21465 3723
rect 21465 3689 21499 3723
rect 21499 3689 21508 3723
rect 21456 3680 21508 3689
rect 21824 3723 21876 3732
rect 21824 3689 21833 3723
rect 21833 3689 21867 3723
rect 21867 3689 21876 3723
rect 21824 3680 21876 3689
rect 22560 3723 22612 3732
rect 22560 3689 22569 3723
rect 22569 3689 22603 3723
rect 22603 3689 22612 3723
rect 22560 3680 22612 3689
rect 23664 3723 23716 3732
rect 23664 3689 23673 3723
rect 23673 3689 23707 3723
rect 23707 3689 23716 3723
rect 23664 3680 23716 3689
rect 12072 3612 12124 3664
rect 13728 3655 13780 3664
rect 13728 3621 13737 3655
rect 13737 3621 13771 3655
rect 13771 3621 13780 3655
rect 13728 3612 13780 3621
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 16580 3612 16632 3664
rect 18972 3612 19024 3664
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 2044 3587 2096 3596
rect 2044 3553 2078 3587
rect 2078 3553 2096 3587
rect 2044 3544 2096 3553
rect 2872 3544 2924 3596
rect 8392 3544 8444 3596
rect 8668 3544 8720 3596
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 11980 3544 12032 3596
rect 12808 3544 12860 3596
rect 14004 3544 14056 3596
rect 14556 3544 14608 3596
rect 17408 3544 17460 3596
rect 17592 3587 17644 3596
rect 17592 3553 17601 3587
rect 17601 3553 17635 3587
rect 17635 3553 17644 3587
rect 17592 3544 17644 3553
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 22008 3587 22060 3596
rect 22008 3553 22017 3587
rect 22017 3553 22051 3587
rect 22051 3553 22060 3587
rect 22008 3544 22060 3553
rect 23112 3587 23164 3596
rect 23112 3553 23121 3587
rect 23121 3553 23155 3587
rect 23155 3553 23164 3587
rect 23112 3544 23164 3553
rect 3332 3476 3384 3528
rect 1768 3340 1820 3392
rect 4436 3340 4488 3392
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 13636 3476 13688 3528
rect 14280 3476 14332 3528
rect 16396 3476 16448 3528
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 20168 3476 20220 3528
rect 12440 3408 12492 3460
rect 6000 3340 6052 3392
rect 8944 3340 8996 3392
rect 11336 3340 11388 3392
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 16580 3383 16632 3392
rect 16580 3349 16589 3383
rect 16589 3349 16623 3383
rect 16623 3349 16632 3383
rect 16580 3340 16632 3349
rect 18880 3408 18932 3460
rect 20812 3408 20864 3460
rect 19432 3340 19484 3392
rect 20444 3383 20496 3392
rect 20444 3349 20453 3383
rect 20453 3349 20487 3383
rect 20487 3349 20496 3383
rect 20444 3340 20496 3349
rect 21088 3383 21140 3392
rect 21088 3349 21097 3383
rect 21097 3349 21131 3383
rect 21131 3349 21140 3383
rect 21088 3340 21140 3349
rect 23296 3383 23348 3392
rect 23296 3349 23305 3383
rect 23305 3349 23339 3383
rect 23339 3349 23348 3383
rect 23296 3340 23348 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1400 3179 1452 3188
rect 1400 3145 1409 3179
rect 1409 3145 1443 3179
rect 1443 3145 1452 3179
rect 1400 3136 1452 3145
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 5540 3136 5592 3188
rect 8484 3136 8536 3188
rect 9680 3136 9732 3188
rect 2136 3000 2188 3052
rect 8024 3111 8076 3120
rect 8024 3077 8033 3111
rect 8033 3077 8067 3111
rect 8067 3077 8076 3111
rect 8024 3068 8076 3077
rect 8392 3111 8444 3120
rect 8392 3077 8401 3111
rect 8401 3077 8435 3111
rect 8435 3077 8444 3111
rect 8392 3068 8444 3077
rect 9864 3068 9916 3120
rect 3516 3000 3568 3052
rect 3792 3000 3844 3052
rect 4436 3000 4488 3052
rect 6920 3000 6972 3052
rect 1676 2932 1728 2984
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 3976 2932 4028 2984
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 3792 2864 3844 2916
rect 4896 2864 4948 2916
rect 6000 2864 6052 2916
rect 6552 2907 6604 2916
rect 6552 2873 6561 2907
rect 6561 2873 6595 2907
rect 6595 2873 6604 2907
rect 6552 2864 6604 2873
rect 9496 2864 9548 2916
rect 10692 3068 10744 3120
rect 11060 3000 11112 3052
rect 11980 3136 12032 3188
rect 13728 3136 13780 3188
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 15476 3136 15528 3188
rect 16028 3136 16080 3188
rect 17500 3136 17552 3188
rect 18420 3136 18472 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 20076 3136 20128 3188
rect 20904 3179 20956 3188
rect 20904 3145 20913 3179
rect 20913 3145 20947 3179
rect 20947 3145 20956 3179
rect 20904 3136 20956 3145
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 23112 3136 23164 3188
rect 23388 3179 23440 3188
rect 23388 3145 23397 3179
rect 23397 3145 23431 3179
rect 23431 3145 23440 3179
rect 23388 3136 23440 3145
rect 15108 3068 15160 3120
rect 15936 3068 15988 3120
rect 11980 3000 12032 3052
rect 11152 2932 11204 2984
rect 16120 3000 16172 3052
rect 17408 3000 17460 3052
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 2964 2839 3016 2848
rect 2964 2805 2973 2839
rect 2973 2805 3007 2839
rect 3007 2805 3016 2839
rect 2964 2796 3016 2805
rect 8116 2796 8168 2848
rect 8392 2796 8444 2848
rect 9772 2796 9824 2848
rect 10692 2796 10744 2848
rect 10968 2796 11020 2848
rect 11336 2864 11388 2916
rect 11980 2864 12032 2916
rect 15568 2932 15620 2984
rect 20628 3068 20680 3120
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 23664 3068 23716 3120
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 21364 2932 21416 2984
rect 22192 2932 22244 2984
rect 23572 2932 23624 2984
rect 14188 2864 14240 2916
rect 14740 2864 14792 2916
rect 17592 2864 17644 2916
rect 18236 2864 18288 2916
rect 20444 2864 20496 2916
rect 13728 2796 13780 2848
rect 14372 2796 14424 2848
rect 18696 2796 18748 2848
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 22192 2796 22244 2848
rect 22560 2796 22612 2848
rect 23848 2839 23900 2848
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1952 2592 2004 2644
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 3516 2635 3568 2644
rect 2044 2592 2096 2601
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 3884 2524 3936 2576
rect 5540 2592 5592 2644
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8300 2592 8352 2644
rect 10692 2592 10744 2644
rect 10968 2592 11020 2644
rect 11428 2635 11480 2644
rect 11428 2601 11437 2635
rect 11437 2601 11471 2635
rect 11471 2601 11480 2635
rect 11980 2635 12032 2644
rect 11428 2592 11480 2601
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 15108 2592 15160 2644
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 17960 2592 18012 2644
rect 20720 2592 20772 2644
rect 22192 2592 22244 2644
rect 13176 2524 13228 2576
rect 14648 2524 14700 2576
rect 3700 2456 3752 2508
rect 5540 2456 5592 2508
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 6092 2456 6144 2508
rect 4988 2388 5040 2397
rect 6828 2388 6880 2440
rect 2412 2295 2464 2304
rect 2412 2261 2421 2295
rect 2421 2261 2455 2295
rect 2455 2261 2464 2295
rect 2412 2252 2464 2261
rect 2504 2252 2556 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 6092 2252 6144 2304
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 9772 2388 9824 2440
rect 11980 2388 12032 2440
rect 7748 2252 7800 2304
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 13728 2388 13780 2440
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 13176 2252 13228 2304
rect 16304 2456 16356 2508
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22192 2456 22244 2508
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 17684 2388 17736 2440
rect 20720 2388 20772 2440
rect 21824 2320 21876 2372
rect 24124 2320 24176 2372
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 19984 2252 20036 2304
rect 23480 2252 23532 2304
rect 24860 2252 24912 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 3148 2048 3200 2100
rect 6552 2048 6604 2100
rect 6552 552 6604 604
rect 7380 552 7432 604
rect 9220 552 9272 604
rect 9404 552 9456 604
rect 21640 552 21692 604
rect 23112 552 23164 604
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 3974 27704 4030 27713
rect 3974 27639 4030 27648
rect 308 20369 336 27520
rect 294 20360 350 20369
rect 294 20295 350 20304
rect 860 17066 888 27520
rect 1412 27418 1440 27520
rect 1412 27390 1532 27418
rect 1400 22500 1452 22506
rect 1400 22442 1452 22448
rect 1412 21690 1440 22442
rect 1400 21684 1452 21690
rect 1400 21626 1452 21632
rect 1504 21418 1532 27390
rect 1860 25288 1912 25294
rect 1860 25230 1912 25236
rect 1584 25220 1636 25226
rect 1584 25162 1636 25168
rect 1596 24750 1624 25162
rect 1872 24818 1900 25230
rect 1860 24812 1912 24818
rect 1860 24754 1912 24760
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1964 24562 1992 27520
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2424 25362 2452 25978
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2424 24954 2452 25298
rect 2412 24948 2464 24954
rect 2412 24890 2464 24896
rect 1596 24534 1992 24562
rect 1492 21412 1544 21418
rect 1492 21354 1544 21360
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1308 19440 1360 19446
rect 1308 19382 1360 19388
rect 1320 17218 1348 19382
rect 1412 18426 1440 21286
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1504 19718 1532 20946
rect 1596 20346 1624 24534
rect 1950 24304 2006 24313
rect 1950 24239 1952 24248
rect 2004 24239 2006 24248
rect 1952 24210 2004 24216
rect 2516 24177 2544 27520
rect 3056 25764 3108 25770
rect 3056 25706 3108 25712
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2502 24168 2558 24177
rect 2502 24103 2558 24112
rect 2410 23896 2466 23905
rect 2410 23831 2412 23840
rect 2464 23831 2466 23840
rect 2412 23802 2464 23808
rect 2424 23662 2452 23802
rect 2412 23656 2464 23662
rect 1858 23624 1914 23633
rect 2412 23598 2464 23604
rect 1858 23559 1860 23568
rect 1912 23559 1914 23568
rect 1860 23530 1912 23536
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2700 23186 2728 23462
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1688 21486 1716 22918
rect 1780 22778 1808 23122
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 2424 22642 2452 22918
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2424 21978 2452 22578
rect 1860 21956 1912 21962
rect 1860 21898 1912 21904
rect 2332 21950 2452 21978
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 1872 21554 1900 21898
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1688 21146 1716 21422
rect 1964 21350 1992 21830
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1872 20466 1900 20878
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1950 20360 2006 20369
rect 1596 20318 1900 20346
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1412 17814 1440 18158
rect 1400 17808 1452 17814
rect 1400 17750 1452 17756
rect 1412 17338 1440 17750
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1320 17190 1440 17218
rect 848 17060 900 17066
rect 848 17002 900 17008
rect 1412 15178 1440 17190
rect 1320 15150 1440 15178
rect 1320 13161 1348 15150
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1306 13152 1362 13161
rect 1306 13087 1362 13096
rect 1412 12782 1440 14214
rect 1504 13802 1532 19654
rect 1596 19446 1624 20198
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 17649 1624 19246
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1688 18601 1716 19178
rect 1674 18592 1730 18601
rect 1674 18527 1730 18536
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1582 17640 1638 17649
rect 1582 17575 1638 17584
rect 1596 16794 1624 17575
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15026 1624 15982
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1492 13796 1544 13802
rect 1492 13738 1544 13744
rect 1688 12986 1716 17711
rect 1780 14550 1808 20198
rect 1872 18222 1900 20318
rect 1950 20295 1952 20304
rect 2004 20295 2006 20304
rect 1952 20266 2004 20272
rect 1964 20058 1992 20266
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1964 18154 1992 18566
rect 2056 18290 2084 20742
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1872 17610 1900 18022
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1766 14240 1822 14249
rect 1766 14175 1822 14184
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1780 12866 1808 14175
rect 1688 12838 1808 12866
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 12306 1532 12718
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 11762 1532 12242
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1412 9518 1440 10746
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1504 9042 1532 11698
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8498 1532 8978
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 294 6352 350 6361
rect 1412 6322 1440 6802
rect 294 6287 350 6296
rect 1400 6316 1452 6322
rect 308 480 336 6287
rect 1400 6258 1452 6264
rect 1412 4146 1440 6258
rect 1504 4690 1532 7142
rect 1596 5030 1624 11222
rect 1688 9586 1716 12838
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11354 1900 12242
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1964 10792 1992 18090
rect 2056 17542 2084 18226
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2042 17096 2098 17105
rect 2042 17031 2098 17040
rect 2056 15978 2084 17031
rect 2044 15972 2096 15978
rect 2044 15914 2096 15920
rect 2056 15706 2084 15914
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2056 15502 2084 15642
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2148 14482 2176 19654
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2240 17134 2268 18022
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2240 16794 2268 17070
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2240 15706 2268 16594
rect 2332 15706 2360 21950
rect 2516 21690 2544 21966
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2686 21448 2742 21457
rect 2424 17105 2452 21422
rect 2504 21412 2556 21418
rect 2686 21383 2742 21392
rect 2504 21354 2556 21360
rect 2516 20890 2544 21354
rect 2516 20862 2636 20890
rect 2608 20806 2636 20862
rect 2596 20800 2648 20806
rect 2596 20742 2648 20748
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 2516 18086 2544 20538
rect 2608 20262 2636 20742
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2410 17096 2466 17105
rect 2410 17031 2466 17040
rect 2410 16960 2466 16969
rect 2410 16895 2466 16904
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2240 15042 2268 15642
rect 2240 15014 2360 15042
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 14618 2268 14826
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2240 14414 2268 14554
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2332 14074 2360 15014
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13025 2360 13670
rect 2424 13258 2452 16895
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2318 13016 2374 13025
rect 2318 12951 2374 12960
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1872 10764 1992 10792
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9110 1716 9318
rect 1676 9104 1728 9110
rect 1872 9081 1900 10764
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1964 10266 1992 10610
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1964 9178 1992 10202
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1858 9072 1914 9081
rect 1676 9046 1728 9052
rect 1780 9030 1858 9058
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7342 1716 7686
rect 1780 7478 1808 9030
rect 1858 9007 1914 9016
rect 1964 8650 1992 9114
rect 1872 8634 1992 8650
rect 1860 8628 1992 8634
rect 1912 8622 1992 8628
rect 1860 8570 1912 8576
rect 1964 8430 1992 8622
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2056 8378 2084 12650
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2240 10198 2268 10406
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 8537 2176 9998
rect 2134 8528 2190 8537
rect 2134 8463 2190 8472
rect 2056 8350 2176 8378
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 2056 7410 2084 7686
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 2056 6934 2084 7346
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1780 5642 1808 6122
rect 2056 6118 2084 6870
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5914 2084 6054
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2148 5817 2176 8350
rect 2240 8090 2268 10134
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2332 6662 2360 11562
rect 2516 11286 2544 17546
rect 2608 16561 2636 20198
rect 2700 20058 2728 21383
rect 2792 21321 2820 25094
rect 2964 24948 3016 24954
rect 2964 24890 3016 24896
rect 2872 24200 2924 24206
rect 2872 24142 2924 24148
rect 2884 23866 2912 24142
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 2884 21350 2912 22102
rect 2976 21865 3004 24890
rect 3068 22166 3096 25706
rect 3056 22160 3108 22166
rect 3056 22102 3108 22108
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 2962 21856 3018 21865
rect 2962 21791 3018 21800
rect 3068 21690 3096 21966
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 2872 21344 2924 21350
rect 2778 21312 2834 21321
rect 2872 21286 2924 21292
rect 2778 21247 2834 21256
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 3068 20262 3096 20402
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2700 19310 2728 19994
rect 3068 19854 3096 20198
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 19009 2728 19110
rect 2686 19000 2742 19009
rect 2686 18935 2742 18944
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2792 18426 2820 18906
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 16946 2728 17478
rect 2792 17338 2820 18226
rect 2884 17882 2912 18702
rect 3068 18290 3096 19382
rect 3160 18970 3188 27520
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 3252 23254 3280 25842
rect 3514 24712 3570 24721
rect 3514 24647 3516 24656
rect 3568 24647 3570 24656
rect 3516 24618 3568 24624
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3240 23248 3292 23254
rect 3240 23190 3292 23196
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3252 20602 3280 22578
rect 3344 21418 3372 24006
rect 3436 23662 3464 24074
rect 3516 23724 3568 23730
rect 3712 23712 3740 27520
rect 3988 26382 4016 27639
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3988 25401 4016 25774
rect 4080 25702 4108 25871
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 3974 25392 4030 25401
rect 3974 25327 4030 25336
rect 4080 24857 4108 25434
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4066 24848 4122 24857
rect 4066 24783 4122 24792
rect 4172 24682 4200 25298
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 3712 23684 3832 23712
rect 3516 23666 3568 23672
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3436 23322 3464 23598
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3528 22982 3556 23666
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22642 3556 22918
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 3436 22030 3464 22510
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3332 21412 3384 21418
rect 3332 21354 3384 21360
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3528 20466 3556 20742
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3160 18193 3188 18906
rect 3252 18737 3280 19314
rect 3238 18728 3294 18737
rect 3238 18663 3294 18672
rect 3344 18630 3372 19314
rect 3620 19310 3648 20198
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3528 18698 3556 19110
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3146 18184 3202 18193
rect 2964 18148 3016 18154
rect 3146 18119 3202 18128
rect 2964 18090 3016 18096
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 17066 2912 17682
rect 2976 17678 3004 18090
rect 3528 17882 3556 18634
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2976 17354 3004 17614
rect 2976 17338 3096 17354
rect 2976 17332 3108 17338
rect 2976 17326 3056 17332
rect 3056 17274 3108 17280
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2700 16918 2912 16946
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2594 16552 2650 16561
rect 2594 16487 2650 16496
rect 2700 16250 2728 16662
rect 2884 16538 2912 16918
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 2964 16584 3016 16590
rect 2884 16532 2964 16538
rect 2884 16526 3016 16532
rect 2884 16510 3004 16526
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3068 15706 3096 16730
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3344 16153 3372 16662
rect 3330 16144 3386 16153
rect 3330 16079 3332 16088
rect 3384 16079 3386 16088
rect 3332 16050 3384 16056
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2594 15328 2650 15337
rect 2594 15263 2650 15272
rect 2608 13938 2636 15263
rect 2700 14618 2728 15506
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3514 15464 3570 15473
rect 3252 15162 3280 15438
rect 3514 15399 3570 15408
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2792 14482 2820 14554
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13462 3096 13874
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12306 2636 12582
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2700 11914 2728 13262
rect 2976 12986 3004 13262
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2976 12442 3004 12922
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2700 11898 2820 11914
rect 2700 11892 2832 11898
rect 2700 11886 2780 11892
rect 2780 11834 2832 11840
rect 2504 11280 2556 11286
rect 2410 11248 2466 11257
rect 2504 11222 2556 11228
rect 2410 11183 2412 11192
rect 2464 11183 2466 11192
rect 2412 11154 2464 11160
rect 2504 11144 2556 11150
rect 2502 11112 2504 11121
rect 2556 11112 2558 11121
rect 2412 11076 2464 11082
rect 2502 11047 2558 11056
rect 2688 11076 2740 11082
rect 2412 11018 2464 11024
rect 2688 11018 2740 11024
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2134 5808 2190 5817
rect 2134 5743 2190 5752
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1584 5024 1636 5030
rect 1582 4992 1584 5001
rect 1636 4992 1638 5001
rect 1582 4927 1638 4936
rect 1872 4826 1900 5063
rect 2240 4826 2268 5510
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 1674 4584 1730 4593
rect 1674 4519 1730 4528
rect 1490 4312 1546 4321
rect 1490 4247 1546 4256
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 846 3632 902 3641
rect 846 3567 902 3576
rect 860 480 888 3567
rect 1412 3194 1440 3839
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1504 3074 1532 4247
rect 1688 3738 1716 4519
rect 2136 4480 2188 4486
rect 1858 4448 1914 4457
rect 2136 4422 2188 4428
rect 1858 4383 1914 4392
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1412 3046 1532 3074
rect 1412 480 1440 3046
rect 1688 2990 1716 3674
rect 1780 3602 1808 4082
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3398 1808 3538
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1872 3074 1900 4383
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1780 3046 1900 3074
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1780 2836 1808 3046
rect 1872 2854 1900 2919
rect 1860 2848 1912 2854
rect 1780 2808 1860 2836
rect 1912 2808 1992 2836
rect 1860 2790 1912 2796
rect 1964 2650 1992 2808
rect 2056 2650 2084 3538
rect 2148 3097 2176 4422
rect 2240 4282 2268 4626
rect 2332 4622 2360 6598
rect 2424 4729 2452 11018
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 10470 2544 10950
rect 2700 10538 2728 11018
rect 2884 10826 2912 12038
rect 2792 10810 2912 10826
rect 2976 10810 3004 12378
rect 3160 11830 3188 12650
rect 3252 12345 3280 14311
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3238 12336 3294 12345
rect 3238 12271 3294 12280
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2780 10804 2912 10810
rect 2832 10798 2912 10804
rect 2964 10804 3016 10810
rect 2780 10746 2832 10752
rect 2964 10746 3016 10752
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2410 4720 2466 4729
rect 2410 4655 2466 4664
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2332 3942 2360 4558
rect 2516 4434 2544 10406
rect 2700 10266 2728 10474
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 9648 2740 9654
rect 2686 9616 2688 9625
rect 2740 9616 2742 9625
rect 2686 9551 2742 9560
rect 2792 9518 2820 10542
rect 3068 10248 3096 11494
rect 3436 11393 3464 14214
rect 3528 13297 3556 15399
rect 3620 14890 3648 19110
rect 3712 18329 3740 21286
rect 3804 19922 3832 23684
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 3974 23488 4030 23497
rect 4172 23474 4200 23598
rect 3974 23423 4030 23432
rect 4080 23446 4200 23474
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3896 22574 3924 22918
rect 3988 22681 4016 23423
rect 4080 23118 4108 23446
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 3974 22672 4030 22681
rect 3974 22607 4030 22616
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 4264 22216 4292 27520
rect 4816 24834 4844 27520
rect 4894 26616 4950 26625
rect 4894 26551 4950 26560
rect 4908 26518 4936 26551
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 5368 25770 5396 27520
rect 5356 25764 5408 25770
rect 5356 25706 5408 25712
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5368 24954 5396 25094
rect 5552 24954 5580 25094
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 5540 24948 5592 24954
rect 5540 24890 5592 24896
rect 4712 24812 4764 24818
rect 4816 24806 5120 24834
rect 5552 24818 5580 24890
rect 6012 24834 6040 27520
rect 4712 24754 4764 24760
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4356 23186 4384 24006
rect 4448 23798 4476 24142
rect 4436 23792 4488 23798
rect 4436 23734 4488 23740
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4356 22234 4384 23122
rect 4434 23080 4490 23089
rect 4434 23015 4490 23024
rect 4080 22188 4292 22216
rect 4344 22228 4396 22234
rect 4080 20398 4108 22188
rect 4344 22170 4396 22176
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4172 21486 4200 22034
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4264 21554 4292 21898
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4172 21146 4200 21422
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4448 21078 4476 23015
rect 4540 22001 4568 24550
rect 4526 21992 4582 22001
rect 4526 21927 4582 21936
rect 4632 21554 4660 24618
rect 4724 23594 4752 24754
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4896 23860 4948 23866
rect 5000 23848 5028 24278
rect 4948 23820 5028 23848
rect 4896 23802 4948 23808
rect 4712 23588 4764 23594
rect 4712 23530 4764 23536
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4816 21350 4844 21966
rect 4894 21448 4950 21457
rect 4894 21383 4950 21392
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4908 21146 4936 21383
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4436 21072 4488 21078
rect 4436 21014 4488 21020
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4080 20058 4108 20334
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4172 19990 4200 20402
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3804 19514 3832 19858
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3804 19281 3832 19450
rect 3790 19272 3846 19281
rect 3790 19207 3846 19216
rect 3896 18970 3924 19926
rect 4068 19848 4120 19854
rect 4264 19825 4292 20198
rect 4068 19790 4120 19796
rect 4250 19816 4306 19825
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 3988 19174 4016 19722
rect 4080 19446 4108 19790
rect 4250 19751 4306 19760
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4068 19304 4120 19310
rect 4120 19264 4200 19292
rect 4068 19246 4120 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3896 18766 3924 18906
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3896 18408 3924 18702
rect 3976 18420 4028 18426
rect 3896 18380 3976 18408
rect 3976 18362 4028 18368
rect 3698 18320 3754 18329
rect 3698 18255 3754 18264
rect 3712 16674 3740 18255
rect 4172 17882 4200 19264
rect 4250 19136 4306 19145
rect 4250 19071 4306 19080
rect 4264 18970 4292 19071
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3974 17232 4030 17241
rect 3974 17167 4030 17176
rect 3712 16646 3832 16674
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3712 15910 3740 16526
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15065 3740 15846
rect 3698 15056 3754 15065
rect 3698 14991 3754 15000
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3712 14414 3740 14991
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3606 13696 3662 13705
rect 3606 13631 3662 13640
rect 3514 13288 3570 13297
rect 3514 13223 3570 13232
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3422 11384 3478 11393
rect 3422 11319 3478 11328
rect 3528 11121 3556 13126
rect 3514 11112 3570 11121
rect 3514 11047 3570 11056
rect 2976 10220 3096 10248
rect 3516 10260 3568 10266
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 9042 2820 9454
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8480 2820 8978
rect 2792 8452 2912 8480
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 8106 2820 8298
rect 2700 8090 2820 8106
rect 2688 8084 2820 8090
rect 2740 8078 2820 8084
rect 2688 8026 2740 8032
rect 2884 8022 2912 8452
rect 2872 8016 2924 8022
rect 2686 7984 2742 7993
rect 2872 7958 2924 7964
rect 2686 7919 2688 7928
rect 2740 7919 2742 7928
rect 2688 7890 2740 7896
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2792 6322 2820 7278
rect 2884 6866 2912 7958
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2608 5370 2636 5714
rect 2884 5710 2912 6054
rect 2688 5704 2740 5710
rect 2872 5704 2924 5710
rect 2740 5664 2820 5692
rect 2688 5646 2740 5652
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2792 5302 2820 5664
rect 2872 5646 2924 5652
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2792 4826 2820 5238
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2700 4570 2728 4762
rect 2700 4542 2912 4570
rect 2516 4406 2728 4434
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2700 3618 2728 4406
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2792 3618 2820 3674
rect 2700 3590 2820 3618
rect 2884 3602 2912 4542
rect 2976 3777 3004 10220
rect 3516 10202 3568 10208
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3054 9616 3110 9625
rect 3054 9551 3110 9560
rect 3068 9518 3096 9551
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 9110 3096 9454
rect 3160 9382 3188 9998
rect 3424 9512 3476 9518
rect 3422 9480 3424 9489
rect 3476 9480 3478 9489
rect 3422 9415 3478 9424
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9178 3188 9318
rect 3528 9178 3556 10202
rect 3620 9450 3648 13631
rect 3698 13152 3754 13161
rect 3698 13087 3754 13096
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3160 8090 3188 9114
rect 3606 8392 3662 8401
rect 3606 8327 3662 8336
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3514 8256 3570 8265
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3160 7886 3188 8026
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 7002 3096 7142
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3146 6896 3202 6905
rect 3146 6831 3202 6840
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 5234 3096 5578
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 4758 3096 5170
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3160 4604 3188 6831
rect 3068 4576 3188 4604
rect 2962 3768 3018 3777
rect 2962 3703 3018 3712
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2976 3482 3004 3703
rect 2884 3454 3004 3482
rect 2134 3088 2190 3097
rect 2134 3023 2136 3032
rect 2188 3023 2190 3032
rect 2136 2994 2188 3000
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2412 2304 2464 2310
rect 1950 2272 2006 2281
rect 2412 2246 2464 2252
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 1950 2207 2006 2216
rect 1964 480 1992 2207
rect 2424 1737 2452 2246
rect 2410 1728 2466 1737
rect 2410 1663 2466 1672
rect 2516 480 2544 2246
rect 2884 649 2912 3454
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 2976 513 3004 2790
rect 3068 1465 3096 4576
rect 3252 4010 3280 8230
rect 3514 8191 3570 8200
rect 3332 4208 3384 4214
rect 3332 4150 3384 4156
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3344 3534 3372 4150
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3528 3233 3556 8191
rect 3620 5545 3648 8327
rect 3712 7342 3740 13087
rect 3804 11218 3832 16646
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3896 15434 3924 15982
rect 3884 15428 3936 15434
rect 3884 15370 3936 15376
rect 3988 14346 4016 17167
rect 4080 16776 4108 17750
rect 4264 17338 4292 18362
rect 4356 17785 4384 20334
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4342 17776 4398 17785
rect 4342 17711 4398 17720
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4080 16748 4200 16776
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 4080 14929 4108 16623
rect 4172 15706 4200 16748
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4160 14952 4212 14958
rect 4066 14920 4122 14929
rect 4160 14894 4212 14900
rect 4066 14855 4122 14864
rect 4172 14550 4200 14894
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 4080 14249 4108 14418
rect 4066 14240 4122 14249
rect 4066 14175 4122 14184
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3896 13308 3924 13942
rect 4160 13320 4212 13326
rect 3896 13280 4160 13308
rect 3896 12442 3924 13280
rect 4160 13262 4212 13268
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 12442 4108 13126
rect 4158 13016 4214 13025
rect 4158 12951 4214 12960
rect 4172 12646 4200 12951
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3988 11830 4016 12242
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3896 10198 3924 11698
rect 3988 11286 4016 11766
rect 4080 11354 4108 12174
rect 4264 11558 4292 17070
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 12481 4384 13670
rect 4342 12472 4398 12481
rect 4342 12407 4398 12416
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4448 11286 4476 20198
rect 5000 19009 5028 23820
rect 4710 19000 4766 19009
rect 4710 18935 4712 18944
rect 4764 18935 4766 18944
rect 4986 19000 5042 19009
rect 4986 18935 5042 18944
rect 4712 18906 4764 18912
rect 5000 18850 5028 18935
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4908 18822 5028 18850
rect 4540 18154 4568 18770
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18426 4844 18702
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4908 18306 4936 18822
rect 5092 18714 5120 24806
rect 5540 24812 5592 24818
rect 6012 24806 6408 24834
rect 5540 24754 5592 24760
rect 6276 24744 6328 24750
rect 6276 24686 6328 24692
rect 5172 24608 5224 24614
rect 5540 24608 5592 24614
rect 5172 24550 5224 24556
rect 5262 24576 5318 24585
rect 5184 23905 5212 24550
rect 5540 24550 5592 24556
rect 5262 24511 5318 24520
rect 5276 24274 5304 24511
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5448 24132 5500 24138
rect 5448 24074 5500 24080
rect 5170 23896 5226 23905
rect 5460 23866 5488 24074
rect 5170 23831 5226 23840
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5552 23730 5580 24550
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6288 23905 6316 24686
rect 6274 23896 6330 23905
rect 6274 23831 6276 23840
rect 6328 23831 6330 23840
rect 6276 23802 6328 23808
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22574 5488 22918
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5448 22568 5500 22574
rect 5552 22545 5580 22714
rect 5448 22510 5500 22516
rect 5538 22536 5594 22545
rect 5538 22471 5594 22480
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 22166 5304 22374
rect 6288 22166 6316 23054
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 5276 21690 5304 22102
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 6196 21622 6224 21830
rect 6184 21616 6236 21622
rect 6182 21584 6184 21593
rect 6236 21584 6238 21593
rect 6182 21519 6238 21528
rect 6196 21493 6224 21519
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5460 21146 5488 21422
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5460 20330 5488 20742
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5184 19990 5212 20198
rect 5552 19990 5580 20946
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20058 6040 21014
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 6104 20602 6132 20878
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6092 20324 6144 20330
rect 6092 20266 6144 20272
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5262 19816 5318 19825
rect 5262 19751 5318 19760
rect 5356 19780 5408 19786
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19242 5212 19654
rect 5172 19236 5224 19242
rect 5172 19178 5224 19184
rect 4816 18278 4936 18306
rect 5000 18686 5120 18714
rect 4618 18184 4674 18193
rect 4528 18148 4580 18154
rect 4618 18119 4674 18128
rect 4528 18090 4580 18096
rect 4540 17882 4568 18090
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4632 17082 4660 18119
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4724 17338 4752 17682
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4816 17134 4844 18278
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4804 17128 4856 17134
rect 4632 17054 4752 17082
rect 4804 17070 4856 17076
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14657 4568 14826
rect 4526 14648 4582 14657
rect 4526 14583 4582 14592
rect 4540 13938 4568 14583
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4528 12912 4580 12918
rect 4528 12854 4580 12860
rect 4540 12374 4568 12854
rect 4632 12617 4660 16934
rect 4724 15570 4752 17054
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16794 4844 16934
rect 4908 16794 4936 17614
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 16250 4844 16594
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 5000 14056 5028 18686
rect 5184 18630 5212 19178
rect 5172 18624 5224 18630
rect 5078 18592 5134 18601
rect 5172 18566 5224 18572
rect 5078 18527 5134 18536
rect 5092 18426 5120 18527
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5092 18222 5120 18362
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5184 18068 5212 18566
rect 5092 18040 5212 18068
rect 5092 17678 5120 18040
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 17338 5120 17614
rect 5276 17354 5304 19751
rect 5356 19722 5408 19728
rect 5368 19553 5396 19722
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5354 19544 5410 19553
rect 5622 19536 5918 19556
rect 5354 19479 5410 19488
rect 6104 19378 6132 20266
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5446 18864 5502 18873
rect 5644 18834 5672 19110
rect 5446 18799 5502 18808
rect 5632 18828 5684 18834
rect 5354 18456 5410 18465
rect 5460 18426 5488 18799
rect 5632 18770 5684 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5354 18391 5410 18400
rect 5448 18420 5500 18426
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5184 17326 5304 17354
rect 5184 16776 5212 17326
rect 5368 17270 5396 18391
rect 5448 18362 5500 18368
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5446 17232 5502 17241
rect 5264 17196 5316 17202
rect 5446 17167 5502 17176
rect 5264 17138 5316 17144
rect 5092 16748 5212 16776
rect 5092 15502 5120 16748
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5184 15910 5212 16594
rect 5276 16522 5304 17138
rect 5354 17096 5410 17105
rect 5354 17031 5410 17040
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5092 14521 5120 15302
rect 5078 14512 5134 14521
rect 5078 14447 5134 14456
rect 5184 14362 5212 15846
rect 5276 15638 5304 16458
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 15178 5304 15438
rect 5368 15337 5396 17031
rect 5460 16250 5488 17167
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5552 16114 5580 17002
rect 6104 16998 6132 17682
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6092 16992 6144 16998
rect 6090 16960 6092 16969
rect 6144 16960 6146 16969
rect 6090 16895 6146 16904
rect 5632 16720 5684 16726
rect 5630 16688 5632 16697
rect 5684 16688 5686 16697
rect 5630 16623 5686 16632
rect 5998 16552 6054 16561
rect 5998 16487 6054 16496
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 6012 16046 6040 16487
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15706 5580 15846
rect 6104 15706 6132 16050
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5354 15328 5410 15337
rect 5354 15263 5410 15272
rect 5276 15150 5396 15178
rect 5460 15162 5488 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 4908 14028 5028 14056
rect 5092 14334 5212 14362
rect 4908 13870 4936 14028
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 5000 13734 5028 13874
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4816 12986 4844 13330
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12986 4936 13262
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5000 12850 5028 13670
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4986 12744 5042 12753
rect 4804 12708 4856 12714
rect 4986 12679 5042 12688
rect 4804 12650 4856 12656
rect 4618 12608 4674 12617
rect 4618 12543 4674 12552
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11898 4752 12174
rect 4816 12102 4844 12650
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4816 11762 4844 12038
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3896 7857 3924 9959
rect 4080 9178 4108 10066
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 8650 4200 9590
rect 3988 8622 4200 8650
rect 3988 7993 4016 8622
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4080 8362 4108 8502
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3974 7984 4030 7993
rect 3974 7919 4030 7928
rect 3882 7848 3938 7857
rect 3882 7783 3938 7792
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3804 7177 3832 7346
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3790 7168 3846 7177
rect 3790 7103 3846 7112
rect 3698 7032 3754 7041
rect 3698 6967 3754 6976
rect 3606 5536 3662 5545
rect 3606 5471 3662 5480
rect 3712 5386 3740 6967
rect 3804 6934 3832 7103
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 3804 5846 3832 6870
rect 3896 6089 3924 7210
rect 3988 6458 4016 7919
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3882 6080 3938 6089
rect 3882 6015 3938 6024
rect 4080 5914 4108 8298
rect 4264 8294 4292 11154
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10606 4384 10950
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4356 9761 4384 10542
rect 4724 10470 4752 11222
rect 4816 11150 4844 11698
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4342 9752 4398 9761
rect 4342 9687 4398 9696
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7750 4292 8230
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3620 5358 3740 5386
rect 3514 3224 3570 3233
rect 3514 3159 3570 3168
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3332 2984 3384 2990
rect 3330 2952 3332 2961
rect 3384 2952 3386 2961
rect 3330 2887 3386 2896
rect 3528 2650 3556 2994
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3054 1456 3110 1465
rect 3054 1391 3110 1400
rect 2962 504 3018 513
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3160 480 3188 2042
rect 3620 2009 3648 5358
rect 4172 5352 4200 6054
rect 3988 5324 4200 5352
rect 3988 5098 4016 5324
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 2514 3740 4422
rect 3804 4321 3832 4966
rect 3790 4312 3846 4321
rect 3790 4247 3792 4256
rect 3844 4247 3846 4256
rect 3792 4218 3844 4224
rect 3804 4187 3832 4218
rect 3882 4176 3938 4185
rect 3882 4111 3938 4120
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3233 3832 3878
rect 3896 3738 3924 4111
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3790 3224 3846 3233
rect 3790 3159 3846 3168
rect 3804 3058 3832 3159
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3606 2000 3662 2009
rect 3606 1935 3662 1944
rect 3712 1465 3740 2450
rect 3698 1456 3754 1465
rect 3698 1391 3754 1400
rect 3804 1034 3832 2858
rect 3896 2582 3924 3674
rect 3988 2990 4016 5034
rect 4066 4720 4122 4729
rect 4066 4655 4068 4664
rect 4120 4655 4122 4664
rect 4068 4626 4120 4632
rect 4264 4457 4292 7686
rect 4356 6905 4384 9687
rect 4448 9382 4476 9998
rect 4540 9382 4568 10134
rect 4632 10062 4660 10406
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9586 4660 9998
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4436 9376 4488 9382
rect 4434 9344 4436 9353
rect 4528 9376 4580 9382
rect 4488 9344 4490 9353
rect 4528 9318 4580 9324
rect 4434 9279 4490 9288
rect 4434 8528 4490 8537
rect 4434 8463 4490 8472
rect 4448 8430 4476 8463
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4342 6896 4398 6905
rect 4342 6831 4398 6840
rect 4436 5840 4488 5846
rect 4342 5808 4398 5817
rect 4436 5782 4488 5788
rect 4342 5743 4398 5752
rect 4356 4758 4384 5743
rect 4448 5234 4476 5782
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4436 5024 4488 5030
rect 4434 4992 4436 5001
rect 4488 4992 4490 5001
rect 4434 4927 4490 4936
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4250 4448 4306 4457
rect 4250 4383 4306 4392
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4080 3194 4108 3606
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 4172 1737 4200 3878
rect 4250 3496 4306 3505
rect 4540 3482 4568 9318
rect 4632 9178 4660 9522
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4632 8974 4660 9114
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8498 4660 8910
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 8090 4660 8434
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4540 3454 4660 3482
rect 4250 3431 4306 3440
rect 4158 1728 4214 1737
rect 4158 1663 4214 1672
rect 3712 1006 3832 1034
rect 3712 480 3740 1006
rect 4264 480 4292 3431
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3058 4476 3334
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4632 1578 4660 3454
rect 4724 2689 4752 10406
rect 5000 10198 5028 12679
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 5092 9738 5120 14334
rect 5262 13696 5318 13705
rect 5262 13631 5318 13640
rect 5276 12782 5304 13631
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5170 11384 5226 11393
rect 5170 11319 5226 11328
rect 5184 10810 5212 11319
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5083 9710 5120 9738
rect 5083 9636 5111 9710
rect 5083 9608 5120 9636
rect 5092 9217 5120 9608
rect 5276 9382 5304 9862
rect 5264 9376 5316 9382
rect 5368 9353 5396 15150
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5540 15088 5592 15094
rect 5538 15056 5540 15065
rect 5592 15056 5594 15065
rect 5538 14991 5594 15000
rect 5538 14920 5594 14929
rect 5538 14855 5594 14864
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5460 14385 5488 14418
rect 5446 14376 5502 14385
rect 5446 14311 5502 14320
rect 5460 14074 5488 14311
rect 5552 14074 5580 14855
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6196 14074 6224 17614
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6288 17377 6316 17546
rect 6274 17368 6330 17377
rect 6274 17303 6330 17312
rect 6288 15570 6316 17303
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15162 6316 15506
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6380 15042 6408 24806
rect 6564 24585 6592 27520
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6550 24576 6606 24585
rect 6550 24511 6606 24520
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 6840 24070 6868 25298
rect 6920 24880 6972 24886
rect 6920 24822 6972 24828
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6656 22778 6684 23802
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6656 22386 6684 22714
rect 6840 22522 6868 24006
rect 6932 22642 6960 24822
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6840 22494 6960 22522
rect 6656 22358 6868 22386
rect 6840 21894 6868 22358
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6564 21350 6592 21830
rect 6932 21554 6960 22494
rect 7012 22160 7064 22166
rect 7012 22102 7064 22108
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6564 20806 6592 21286
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6564 19990 6592 20742
rect 6840 20398 6868 20742
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6564 19310 6592 19926
rect 6918 19680 6974 19689
rect 6918 19615 6974 19624
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6564 18630 6592 19246
rect 6932 19145 6960 19615
rect 6918 19136 6974 19145
rect 6918 19071 6974 19080
rect 7024 18970 7052 22102
rect 7116 22098 7144 27520
rect 7668 26466 7696 27520
rect 7668 26438 8156 26466
rect 7472 25968 7524 25974
rect 7472 25910 7524 25916
rect 7484 25430 7512 25910
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 7576 24954 7604 25298
rect 7852 25158 7880 25298
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24274 7236 24754
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7208 23594 7236 24210
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7300 23186 7328 24006
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7392 22778 7420 23122
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7116 20505 7144 20946
rect 7208 20602 7236 21014
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7102 20496 7158 20505
rect 7102 20431 7158 20440
rect 7116 20398 7144 20431
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19938 7144 20334
rect 7300 20330 7328 21898
rect 7378 20632 7434 20641
rect 7378 20567 7434 20576
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7392 20058 7420 20567
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7116 19910 7236 19938
rect 7208 19854 7236 19910
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7208 19514 7236 19790
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7392 19378 7420 19994
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7288 19304 7340 19310
rect 7102 19272 7158 19281
rect 7288 19246 7340 19252
rect 7102 19207 7158 19216
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6564 17882 6592 18566
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 16794 6592 17614
rect 6920 16992 6972 16998
rect 7116 16946 7144 19207
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18222 7236 18566
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7208 17542 7236 18022
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17241 7236 17478
rect 7194 17232 7250 17241
rect 7194 17167 7250 17176
rect 6920 16934 6972 16940
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6550 16552 6606 16561
rect 6550 16487 6606 16496
rect 6458 16008 6514 16017
rect 6458 15943 6514 15952
rect 6472 15638 6500 15943
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6288 15014 6408 15042
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 5460 12322 5488 14010
rect 6196 13870 6224 14010
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12442 5580 13330
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5460 12294 5580 12322
rect 5552 12170 5580 12294
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11354 6040 13262
rect 6288 12481 6316 15014
rect 6472 14822 6500 15438
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13326 6408 14214
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12646 6408 13262
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6274 12472 6330 12481
rect 6274 12407 6330 12416
rect 6184 12368 6236 12374
rect 6182 12336 6184 12345
rect 6236 12336 6238 12345
rect 6182 12271 6238 12280
rect 6196 11898 6224 12271
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5446 10840 5502 10849
rect 5446 10775 5502 10784
rect 5460 10742 5488 10775
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5552 10690 5580 11154
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10690 6040 10950
rect 6104 10849 6132 11494
rect 6090 10840 6146 10849
rect 6090 10775 6146 10784
rect 5552 10662 5672 10690
rect 6012 10674 6132 10690
rect 6012 10668 6144 10674
rect 6012 10662 6092 10668
rect 5540 10600 5592 10606
rect 5538 10568 5540 10577
rect 5592 10568 5594 10577
rect 5538 10503 5594 10512
rect 5644 10169 5672 10662
rect 6092 10610 6144 10616
rect 5630 10160 5686 10169
rect 5630 10095 5632 10104
rect 5684 10095 5686 10104
rect 6000 10124 6052 10130
rect 5632 10066 5684 10072
rect 6000 10066 6052 10072
rect 5644 10010 5672 10066
rect 5552 9982 5672 10010
rect 5448 9376 5500 9382
rect 5264 9318 5316 9324
rect 5354 9344 5410 9353
rect 5078 9208 5134 9217
rect 5078 9143 5134 9152
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4816 8362 4844 8978
rect 4908 8634 4936 9046
rect 5092 8673 5120 9143
rect 5078 8664 5134 8673
rect 4896 8628 4948 8634
rect 5078 8599 5134 8608
rect 4896 8570 4948 8576
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4710 2680 4766 2689
rect 4710 2615 4766 2624
rect 4710 1592 4766 1601
rect 4632 1550 4710 1578
rect 4710 1527 4766 1536
rect 4724 921 4752 1527
rect 4710 912 4766 921
rect 4710 847 4766 856
rect 4816 480 4844 8298
rect 5276 8265 5304 9318
rect 5448 9318 5500 9324
rect 5354 9279 5410 9288
rect 5460 8838 5488 9318
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8362 5488 8774
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5262 8256 5318 8265
rect 5552 8242 5580 9982
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5908 9036 5960 9042
rect 6012 9024 6040 10066
rect 5960 8996 6040 9024
rect 5908 8978 5960 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5262 8191 5318 8200
rect 5368 8214 5580 8242
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6866 4936 7142
rect 5000 6934 5028 7958
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7546 5212 7822
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5184 7002 5212 7482
rect 5368 7478 5396 8214
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 4988 6928 5040 6934
rect 5040 6888 5120 6916
rect 4988 6870 5040 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6458 4936 6802
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4908 5914 4936 6394
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3097 4936 3878
rect 4894 3088 4950 3097
rect 4894 3023 4950 3032
rect 4908 2922 4936 3023
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 5000 2446 5028 6054
rect 5092 5778 5120 6888
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5276 5370 5304 5782
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5368 4078 5396 5306
rect 5460 4808 5488 7686
rect 5552 6662 5580 8026
rect 6104 7936 6132 10610
rect 6196 8634 6224 11834
rect 6288 11150 6316 12174
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10810 6316 11086
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6276 10464 6328 10470
rect 6380 10452 6408 11154
rect 6472 11121 6500 14758
rect 6458 11112 6514 11121
rect 6458 11047 6514 11056
rect 6328 10424 6408 10452
rect 6276 10406 6328 10412
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6012 7908 6132 7936
rect 6184 7948 6236 7954
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7528 6040 7908
rect 6184 7890 6236 7896
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 5920 7500 6040 7528
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5644 7041 5672 7414
rect 5630 7032 5686 7041
rect 5630 6967 5686 6976
rect 5920 6730 5948 7500
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6012 6866 6040 7346
rect 6104 7002 6132 7754
rect 6196 7041 6224 7890
rect 6288 7274 6316 10406
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9450 6408 10066
rect 6564 9654 6592 16487
rect 6932 16114 6960 16934
rect 7024 16918 7144 16946
rect 7024 16794 7052 16918
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7024 15910 7052 16730
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6642 15736 6698 15745
rect 6642 15671 6644 15680
rect 6696 15671 6698 15680
rect 6644 15642 6696 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 13002 6684 13738
rect 6748 13530 6776 15506
rect 6840 13818 6868 15846
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14414 6960 14894
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 14074 6960 14350
rect 7024 14278 7052 14826
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6932 13920 6960 14010
rect 6932 13892 7052 13920
rect 6840 13790 6960 13818
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6656 12974 6776 13002
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6366 9344 6422 9353
rect 6366 9279 6422 9288
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6182 7032 6238 7041
rect 6092 6996 6144 7002
rect 6182 6967 6238 6976
rect 6092 6938 6144 6944
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6322 6040 6802
rect 6104 6458 6132 6938
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5953 5672 6054
rect 5630 5944 5686 5953
rect 5630 5879 5686 5888
rect 6104 5846 6132 6394
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6196 5302 6224 6967
rect 6276 6724 6328 6730
rect 6276 6666 6328 6672
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5540 4820 5592 4826
rect 5460 4780 5540 4808
rect 5540 4762 5592 4768
rect 5736 4593 5764 4966
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5722 4584 5778 4593
rect 5540 4548 5592 4554
rect 5722 4519 5778 4528
rect 5540 4490 5592 4496
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5184 2394 5212 3878
rect 5460 3641 5488 4422
rect 5552 4146 5580 4490
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5552 3670 5580 4082
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5736 3913 5764 3946
rect 5722 3904 5778 3913
rect 5722 3839 5778 3848
rect 6012 3738 6040 4762
rect 6104 4622 6132 5034
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 4214 6132 4558
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5540 3664 5592 3670
rect 5446 3632 5502 3641
rect 5540 3606 5592 3612
rect 5446 3567 5502 3576
rect 5552 3194 5580 3606
rect 6000 3392 6052 3398
rect 6104 3369 6132 3878
rect 6196 3738 6224 4694
rect 6288 3942 6316 6666
rect 6380 5545 6408 9279
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6472 7750 6500 8978
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6366 5536 6422 5545
rect 6366 5471 6422 5480
rect 6472 5273 6500 7686
rect 6564 7546 6592 7958
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6361 6592 7142
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6458 5264 6514 5273
rect 6458 5199 6514 5208
rect 6564 5098 6592 5510
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4010 6500 4422
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6000 3334 6052 3340
rect 6090 3360 6146 3369
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5354 2952 5410 2961
rect 5354 2887 5410 2896
rect 5184 2366 5304 2394
rect 5172 2304 5224 2310
rect 5170 2272 5172 2281
rect 5224 2272 5226 2281
rect 5170 2207 5226 2216
rect 5276 1057 5304 2366
rect 5262 1048 5318 1057
rect 5262 983 5318 992
rect 5368 480 5396 2887
rect 5552 2650 5580 3130
rect 6012 2961 6040 3334
rect 6090 3295 6146 3304
rect 6656 3210 6684 12854
rect 6748 9722 6776 12974
rect 6840 12306 6868 13670
rect 6932 13394 6960 13790
rect 7024 13530 7052 13892
rect 7208 13530 7236 15438
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 11898 6868 12242
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 10198 6868 11630
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6932 9518 6960 12718
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12442 7052 12582
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7102 10704 7158 10713
rect 7102 10639 7104 10648
rect 7156 10639 7158 10648
rect 7104 10610 7156 10616
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7208 9518 7236 9658
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6932 8974 6960 9454
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7024 9042 7052 9318
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7116 8820 7144 9386
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 9110 7236 9318
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7196 8832 7248 8838
rect 7116 8800 7196 8820
rect 7248 8800 7250 8809
rect 7116 8792 7194 8800
rect 7194 8735 7250 8744
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 7102 8256 7158 8265
rect 6840 8090 6868 8230
rect 7300 8242 7328 19246
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 17513 7420 17614
rect 7378 17504 7434 17513
rect 7378 17439 7434 17448
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7392 13802 7420 16458
rect 7484 13954 7512 22034
rect 7576 19310 7604 24550
rect 7746 23760 7802 23769
rect 7746 23695 7802 23704
rect 7760 23662 7788 23695
rect 7748 23656 7800 23662
rect 7748 23598 7800 23604
rect 7852 22778 7880 25094
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 21894 7788 22034
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 8024 21888 8076 21894
rect 8024 21830 8076 21836
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7668 19553 7696 19858
rect 7654 19544 7710 19553
rect 7654 19479 7656 19488
rect 7708 19479 7710 19488
rect 7656 19450 7708 19456
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7668 18306 7696 19450
rect 7760 19174 7788 21830
rect 8036 21486 8064 21830
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7932 21412 7984 21418
rect 7932 21354 7984 21360
rect 7944 20058 7972 21354
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7944 19378 7972 19994
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7852 18714 7880 19314
rect 7852 18686 7972 18714
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7576 18278 7696 18306
rect 7746 18320 7802 18329
rect 7852 18290 7880 18566
rect 7576 16697 7604 18278
rect 7746 18255 7748 18264
rect 7800 18255 7802 18264
rect 7840 18284 7892 18290
rect 7748 18226 7800 18232
rect 7840 18226 7892 18232
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 17746 7696 18158
rect 7852 17882 7880 18226
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7746 17776 7802 17785
rect 7656 17740 7708 17746
rect 7746 17711 7802 17720
rect 7656 17682 7708 17688
rect 7668 16998 7696 17682
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7760 16794 7788 17711
rect 7852 17338 7880 17818
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7562 16688 7618 16697
rect 7562 16623 7618 16632
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 16114 7604 16390
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7576 14385 7604 16050
rect 7852 15978 7880 16526
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 14822 7696 15438
rect 7746 15192 7802 15201
rect 7746 15127 7802 15136
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7668 14550 7696 14758
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7562 14376 7618 14385
rect 7562 14311 7618 14320
rect 7668 14074 7696 14486
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7484 13926 7696 13954
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7378 13424 7434 13433
rect 7378 13359 7434 13368
rect 7392 12986 7420 13359
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7392 11694 7420 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7378 11112 7434 11121
rect 7378 11047 7380 11056
rect 7432 11047 7434 11056
rect 7380 11018 7432 11024
rect 7392 10810 7420 11018
rect 7484 11014 7512 11562
rect 7472 11008 7524 11014
rect 7470 10976 7472 10985
rect 7524 10976 7526 10985
rect 7470 10911 7526 10920
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7484 10266 7512 10911
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8498 7512 8774
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7158 8214 7328 8242
rect 7378 8256 7434 8265
rect 7102 8191 7158 8200
rect 7378 8191 7434 8200
rect 7116 8090 7144 8191
rect 7392 8090 7420 8191
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 5370 6776 7686
rect 7116 7546 7144 8026
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6840 4826 6868 6054
rect 6932 5778 6960 7142
rect 7208 7002 7236 7822
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7410 7420 7754
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6932 4758 6960 5714
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 4826 7052 5646
rect 7102 5536 7158 5545
rect 7102 5471 7158 5480
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3777 7052 3878
rect 7010 3768 7066 3777
rect 7010 3703 7066 3712
rect 6196 3182 6684 3210
rect 5998 2952 6054 2961
rect 5998 2887 6000 2896
rect 6052 2887 6054 2896
rect 6000 2858 6052 2864
rect 6012 2827 6040 2858
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5552 2514 5580 2586
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6104 2310 6132 2450
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 2009 6132 2246
rect 6090 2000 6146 2009
rect 6090 1935 6146 1944
rect 6196 1442 6224 3182
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6564 2106 6592 2858
rect 6932 2530 6960 2994
rect 6840 2502 6960 2530
rect 6840 2446 6868 2502
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6012 1414 6224 1442
rect 6012 480 6040 1414
rect 6552 604 6604 610
rect 6552 546 6604 552
rect 6564 480 6592 546
rect 7116 480 7144 5471
rect 7208 2961 7236 6938
rect 7300 6662 7328 7278
rect 7392 6934 7420 7346
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 4282 7328 6598
rect 7392 6458 7420 6870
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5914 7420 6054
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7576 4826 7604 11834
rect 7668 9178 7696 13926
rect 7760 13530 7788 15127
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7760 12374 7788 13466
rect 7944 13002 7972 18686
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8036 15366 8064 16526
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7852 12974 7972 13002
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7852 11898 7880 12974
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10742 7788 11154
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7852 10577 7880 11018
rect 7838 10568 7894 10577
rect 7838 10503 7894 10512
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7668 6610 7696 9114
rect 7760 6769 7788 10066
rect 7944 9330 7972 12650
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8036 10441 8064 10542
rect 8022 10432 8078 10441
rect 8022 10367 8078 10376
rect 8036 10198 8064 10367
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7852 9302 7972 9330
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7852 8401 7880 9302
rect 8036 9178 8064 9318
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 8968 7984 8974
rect 8036 8945 8064 8978
rect 7932 8910 7984 8916
rect 8022 8936 8078 8945
rect 7838 8392 7894 8401
rect 7838 8327 7894 8336
rect 7944 8090 7972 8910
rect 8022 8871 8078 8880
rect 8036 8634 8064 8871
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7746 6760 7802 6769
rect 7746 6695 7802 6704
rect 8036 6662 8064 8434
rect 8024 6656 8076 6662
rect 7668 6582 7880 6610
rect 8024 6598 8076 6604
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 3942 7328 4218
rect 7576 4214 7604 4762
rect 7668 4622 7696 6394
rect 7746 5264 7802 5273
rect 7746 5199 7802 5208
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4214 7696 4558
rect 7564 4208 7616 4214
rect 7378 4176 7434 4185
rect 7564 4150 7616 4156
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7378 4111 7434 4120
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7194 2952 7250 2961
rect 7194 2887 7250 2896
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 1873 7236 2246
rect 7194 1864 7250 1873
rect 7194 1799 7250 1808
rect 7392 610 7420 4111
rect 7760 3738 7788 5199
rect 7852 4690 7880 6582
rect 8036 6186 8064 6598
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5710 8064 6122
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 4826 8064 5646
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 1465 7788 2246
rect 7746 1456 7802 1465
rect 7746 1391 7802 1400
rect 7852 1306 7880 3606
rect 7668 1278 7880 1306
rect 7380 604 7432 610
rect 7380 546 7432 552
rect 7668 480 7696 1278
rect 7944 921 7972 4218
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8036 3534 8064 4082
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8036 3126 8064 3470
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8128 2854 8156 26438
rect 8220 24177 8248 27520
rect 8298 27160 8354 27169
rect 8298 27095 8354 27104
rect 8312 25158 8340 27095
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8404 24614 8432 25230
rect 8576 24744 8628 24750
rect 8574 24712 8576 24721
rect 8628 24712 8630 24721
rect 8864 24682 8892 27520
rect 9416 24857 9444 27520
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9402 24848 9458 24857
rect 9402 24783 9458 24792
rect 8574 24647 8630 24656
rect 8852 24676 8904 24682
rect 8852 24618 8904 24624
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 8206 24168 8262 24177
rect 8206 24103 8262 24112
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8312 23905 8340 24006
rect 8298 23896 8354 23905
rect 8298 23831 8354 23840
rect 8404 23526 8432 24550
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8588 23594 8616 24006
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8208 23520 8260 23526
rect 8392 23520 8444 23526
rect 8260 23480 8340 23508
rect 8208 23462 8260 23468
rect 8312 23322 8340 23480
rect 8392 23462 8444 23468
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8404 23186 8432 23462
rect 8772 23225 8800 24550
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 8850 23760 8906 23769
rect 8850 23695 8906 23704
rect 8758 23216 8814 23225
rect 8392 23180 8444 23186
rect 8758 23151 8814 23160
rect 8392 23122 8444 23128
rect 8206 22808 8262 22817
rect 8864 22778 8892 23695
rect 9140 23322 9168 24006
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9324 22778 9352 22986
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 8206 22743 8262 22752
rect 8852 22772 8904 22778
rect 8220 22642 8248 22743
rect 8852 22714 8904 22720
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 9508 22574 9536 22918
rect 9692 22778 9720 25978
rect 9968 24834 9996 27520
rect 10520 25786 10548 27520
rect 9784 24806 9996 24834
rect 10060 25758 10548 25786
rect 11072 25786 11100 27520
rect 11244 25832 11296 25838
rect 11072 25758 11192 25786
rect 11244 25774 11296 25780
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8220 21962 8248 22374
rect 9508 22234 9536 22510
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 8576 22024 8628 22030
rect 8496 21984 8576 22012
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8404 21486 8432 21830
rect 8496 21690 8524 21984
rect 8576 21966 8628 21972
rect 8760 21956 8812 21962
rect 8760 21898 8812 21904
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8220 20874 8248 21422
rect 8404 21146 8432 21422
rect 8772 21146 8800 21898
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 9508 21078 9536 21626
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9496 21072 9548 21078
rect 9402 21040 9458 21049
rect 9496 21014 9548 21020
rect 9402 20975 9404 20984
rect 9456 20975 9458 20984
rect 9404 20946 9456 20952
rect 9218 20904 9274 20913
rect 8208 20868 8260 20874
rect 9218 20839 9274 20848
rect 8208 20810 8260 20816
rect 9232 20602 9260 20839
rect 9220 20596 9272 20602
rect 9220 20538 9272 20544
rect 9416 20534 9444 20946
rect 9494 20904 9550 20913
rect 9494 20839 9496 20848
rect 9548 20839 9550 20848
rect 9496 20810 9548 20816
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 8574 20088 8630 20097
rect 8574 20023 8630 20032
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8404 19292 8432 19858
rect 8298 19272 8354 19281
rect 8404 19264 8524 19292
rect 8298 19207 8354 19216
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8220 18970 8248 19110
rect 8312 18970 8340 19207
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8312 18714 8340 18906
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8220 18686 8340 18714
rect 8220 18358 8248 18686
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8312 17134 8340 18566
rect 8404 18358 8432 18770
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8404 17785 8432 18294
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 16794 8340 17070
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8220 16674 8248 16730
rect 8220 16646 8340 16674
rect 8312 16250 8340 16646
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8404 16046 8432 16390
rect 8392 16040 8444 16046
rect 8390 16008 8392 16017
rect 8444 16008 8446 16017
rect 8390 15943 8446 15952
rect 8496 15638 8524 19264
rect 8588 16250 8616 20023
rect 8666 19816 8722 19825
rect 8666 19751 8722 19760
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8220 14804 8248 15506
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8484 14816 8536 14822
rect 8220 14776 8484 14804
rect 8484 14758 8536 14764
rect 8496 14074 8524 14758
rect 8588 14278 8616 15302
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13258 8432 13670
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 11830 8248 12242
rect 8208 11824 8260 11830
rect 8206 11792 8208 11801
rect 8260 11792 8262 11801
rect 8206 11727 8262 11736
rect 8220 11354 8248 11727
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8484 11280 8536 11286
rect 8298 11248 8354 11257
rect 8484 11222 8536 11228
rect 8298 11183 8354 11192
rect 8392 11212 8444 11218
rect 8312 10033 8340 11183
rect 8392 11154 8444 11160
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8404 9568 8432 11154
rect 8496 10130 8524 11222
rect 8588 10606 8616 14214
rect 8680 12986 8708 19751
rect 8772 13530 8800 20470
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8956 19417 8984 20198
rect 9692 20058 9720 21082
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 8942 19408 8998 19417
rect 9416 19378 9444 19654
rect 8942 19343 8998 19352
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9232 18737 9260 19110
rect 9218 18728 9274 18737
rect 9218 18663 9274 18672
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18426 9076 18566
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 18290 9076 18362
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17202 9168 17478
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16726 8892 17070
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 9232 16522 9260 17206
rect 9324 17134 9352 19110
rect 9416 18766 9444 19314
rect 9692 19310 9720 19858
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9404 18624 9456 18630
rect 9508 18578 9536 19110
rect 9692 18970 9720 19246
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9456 18572 9536 18578
rect 9404 18566 9536 18572
rect 9416 18550 9536 18566
rect 9416 18193 9444 18550
rect 9402 18184 9458 18193
rect 9402 18119 9458 18128
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9416 17542 9444 18022
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9404 17536 9456 17542
rect 9600 17513 9628 17682
rect 9404 17478 9456 17484
rect 9586 17504 9642 17513
rect 9416 17338 9444 17478
rect 9586 17439 9642 17448
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9232 16250 9260 16458
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 9048 14618 9076 15574
rect 9036 14612 9088 14618
rect 8956 14572 9036 14600
rect 8956 14482 8984 14572
rect 9036 14554 9088 14560
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8956 13530 8984 14418
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 13530 9076 13670
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9416 13326 9444 17002
rect 9600 15638 9628 17439
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9496 15564 9548 15570
rect 9496 15506 9548 15512
rect 9508 15162 9536 15506
rect 9586 15464 9642 15473
rect 9586 15399 9588 15408
rect 9640 15399 9642 15408
rect 9588 15370 9640 15376
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9508 13870 9536 14418
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9692 13394 9720 16662
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8942 13016 8998 13025
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8852 12980 8904 12986
rect 8942 12951 8998 12960
rect 8852 12922 8904 12928
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8588 10266 8616 10542
rect 8680 10441 8708 12786
rect 8864 12753 8892 12922
rect 8956 12850 8984 12951
rect 9126 12880 9182 12889
rect 8944 12844 8996 12850
rect 9126 12815 9182 12824
rect 8944 12786 8996 12792
rect 8850 12744 8906 12753
rect 8850 12679 8906 12688
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8666 10432 8722 10441
rect 8666 10367 8722 10376
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8312 9540 8432 9568
rect 8312 5409 8340 9540
rect 8588 8974 8616 10202
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8392 8424 8444 8430
rect 8390 8392 8392 8401
rect 8444 8392 8446 8401
rect 8390 8327 8446 8336
rect 8588 8090 8616 8910
rect 8666 8528 8722 8537
rect 8666 8463 8722 8472
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8574 7984 8630 7993
rect 8574 7919 8576 7928
rect 8628 7919 8630 7928
rect 8576 7890 8628 7896
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 6866 8616 7346
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8588 6322 8616 6802
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8298 5400 8354 5409
rect 8298 5335 8354 5344
rect 8588 5166 8616 6258
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4214 8340 4626
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8392 4072 8444 4078
rect 8206 4040 8262 4049
rect 8392 4014 8444 4020
rect 8206 3975 8262 3984
rect 8300 4004 8352 4010
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8128 2553 8156 2586
rect 8114 2544 8170 2553
rect 8114 2479 8170 2488
rect 7930 912 7986 921
rect 7930 847 7986 856
rect 8220 480 8248 3975
rect 8300 3946 8352 3952
rect 8312 2650 8340 3946
rect 8404 3738 8432 4014
rect 8496 4010 8524 4422
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 3126 8432 3538
rect 8496 3194 8524 3946
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3120 8444 3126
rect 8588 3074 8616 5102
rect 8680 3602 8708 8463
rect 8772 8022 8800 11630
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8772 7002 8800 7958
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8772 3942 8800 3975
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8392 3062 8444 3068
rect 8496 3046 8616 3074
rect 8496 2990 8524 3046
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2281 8432 2790
rect 8390 2272 8446 2281
rect 8390 2207 8446 2216
rect 8864 480 8892 7783
rect 8956 7721 8984 12582
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9518 9076 9862
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 8634 9076 9454
rect 9140 9058 9168 12815
rect 9232 12782 9260 13126
rect 9312 12980 9364 12986
rect 9416 12968 9444 13262
rect 9588 13252 9640 13258
rect 9640 13212 9720 13240
rect 9588 13194 9640 13200
rect 9364 12940 9444 12968
rect 9312 12922 9364 12928
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9232 12102 9260 12718
rect 9310 12608 9366 12617
rect 9310 12543 9366 12552
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9140 9030 9260 9058
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8498 9168 8910
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9232 8378 9260 9030
rect 9324 8566 9352 12543
rect 9692 12442 9720 13212
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9416 11762 9444 12038
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9416 11393 9444 11562
rect 9402 11384 9458 11393
rect 9402 11319 9404 11328
rect 9456 11319 9458 11328
rect 9404 11290 9456 11296
rect 9416 11259 9444 11290
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 11121 9628 11154
rect 9586 11112 9642 11121
rect 9586 11047 9642 11056
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10266 9444 10950
rect 9692 10554 9720 12038
rect 9784 11626 9812 24806
rect 9864 24744 9916 24750
rect 9862 24712 9864 24721
rect 9916 24712 9918 24721
rect 9862 24647 9918 24656
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 24449 9904 24550
rect 9862 24440 9918 24449
rect 9862 24375 9918 24384
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9862 24032 9918 24041
rect 9862 23967 9918 23976
rect 9876 22098 9904 23967
rect 9968 23526 9996 24210
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9968 23050 9996 23462
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9876 21570 9904 22034
rect 9968 21690 9996 22714
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9876 21542 9996 21570
rect 9968 21350 9996 21542
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 20602 9904 21014
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9862 20224 9918 20233
rect 9862 20159 9918 20168
rect 9876 17134 9904 20159
rect 9968 17270 9996 21286
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9876 16250 9904 16934
rect 9968 16794 9996 17002
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 16726 10088 25758
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 11072 25498 11100 25638
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10612 24954 10640 25298
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10152 23662 10180 24006
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10784 23588 10836 23594
rect 10784 23530 10836 23536
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10796 23322 10824 23530
rect 10784 23316 10836 23322
rect 10784 23258 10836 23264
rect 10322 23216 10378 23225
rect 10322 23151 10324 23160
rect 10376 23151 10378 23160
rect 10324 23122 10376 23128
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10152 22778 10180 23054
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10336 22710 10364 23122
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10796 22574 10824 23258
rect 11072 22953 11100 24210
rect 11058 22944 11114 22953
rect 11058 22879 11114 22888
rect 10966 22808 11022 22817
rect 10966 22743 11022 22752
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10980 22522 11008 22743
rect 11072 22710 11100 22879
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11164 22522 11192 25758
rect 11256 24410 11284 25774
rect 11716 24562 11744 27520
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12072 24608 12124 24614
rect 11716 24534 12020 24562
rect 12072 24550 12124 24556
rect 11244 24404 11296 24410
rect 11244 24346 11296 24352
rect 11518 24168 11574 24177
rect 11518 24103 11574 24112
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 23769 11284 24006
rect 11242 23760 11298 23769
rect 11242 23695 11298 23704
rect 11242 22808 11298 22817
rect 11242 22743 11298 22752
rect 11256 22642 11284 22743
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 10980 22494 11192 22522
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22024 10192 22030
rect 10192 21984 10272 22012
rect 10140 21966 10192 21972
rect 10244 21729 10272 21984
rect 10888 21894 10916 22374
rect 11428 22092 11480 22098
rect 11428 22034 11480 22040
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10230 21720 10286 21729
rect 10230 21655 10286 21664
rect 10244 21622 10272 21655
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21146 10732 21286
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10244 20398 10272 20946
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10324 19984 10376 19990
rect 10324 19926 10376 19932
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 18970 10180 19790
rect 10336 19310 10364 19926
rect 10888 19786 10916 21830
rect 11256 21554 11284 21898
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11072 20330 11100 21082
rect 11150 20904 11206 20913
rect 11150 20839 11206 20848
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 20058 11100 20266
rect 11164 20074 11192 20839
rect 11256 20244 11284 21490
rect 11348 21486 11376 21830
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11348 21146 11376 21422
rect 11440 21350 11468 22034
rect 11428 21344 11480 21350
rect 11426 21312 11428 21321
rect 11480 21312 11482 21321
rect 11426 21247 11482 21256
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11426 20360 11482 20369
rect 11426 20295 11482 20304
rect 11336 20256 11388 20262
rect 11256 20216 11336 20244
rect 11336 20198 11388 20204
rect 11060 20052 11112 20058
rect 11164 20046 11284 20074
rect 11060 19994 11112 20000
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10324 19304 10376 19310
rect 10322 19272 10324 19281
rect 10376 19272 10378 19281
rect 10322 19207 10378 19216
rect 10336 19181 10364 19207
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 18426 10364 18770
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10336 18290 10364 18362
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9968 16114 9996 16458
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9968 15638 9996 16050
rect 10060 15706 10088 16526
rect 10244 16182 10272 16594
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9876 14822 9904 15438
rect 10152 15162 10180 15914
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15156 10192 15162
rect 10704 15144 10732 19722
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10782 19272 10838 19281
rect 10782 19207 10838 19216
rect 10796 18426 10824 19207
rect 10980 18952 11008 19314
rect 11164 19310 11192 19654
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10980 18924 11100 18952
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10796 16794 10824 17682
rect 10888 17678 10916 18566
rect 10980 17882 11008 18770
rect 11072 18426 11100 18924
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10980 17202 11008 17818
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10874 16688 10930 16697
rect 10874 16623 10930 16632
rect 10888 16250 10916 16623
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10888 16046 10916 16186
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10782 15736 10838 15745
rect 10782 15671 10838 15680
rect 10796 15473 10824 15671
rect 11072 15502 11100 18362
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11060 15496 11112 15502
rect 10782 15464 10838 15473
rect 10782 15399 10838 15408
rect 10980 15444 11060 15450
rect 10980 15438 11112 15444
rect 10980 15422 11100 15438
rect 10980 15162 11008 15422
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10968 15156 11020 15162
rect 10704 15116 10916 15144
rect 10140 15098 10192 15104
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9954 14784 10010 14793
rect 9876 12209 9904 14758
rect 9954 14719 10010 14728
rect 9862 12200 9918 12209
rect 9862 12135 9918 12144
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9876 11234 9904 12135
rect 9784 11206 9904 11234
rect 9784 10674 9812 11206
rect 9864 11144 9916 11150
rect 9968 11132 9996 14719
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14962
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10060 13530 10088 14350
rect 10796 14074 10824 14486
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 12986 10088 13466
rect 10152 13308 10180 13806
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10796 13530 10824 14010
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10888 13410 10916 15116
rect 10968 15098 11020 15104
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10980 14278 11008 14826
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10704 13382 10916 13410
rect 10324 13320 10376 13326
rect 10152 13280 10324 13308
rect 10324 13262 10376 13268
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10336 12918 10364 13262
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 11830 10088 12786
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12424 10732 13382
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12646 10824 13262
rect 10874 12744 10930 12753
rect 10874 12679 10930 12688
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10612 12396 10732 12424
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10152 11898 10180 12174
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10336 11830 10364 12174
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 12073 10548 12106
rect 10612 12102 10640 12396
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10600 12096 10652 12102
rect 10506 12064 10562 12073
rect 10600 12038 10652 12044
rect 10506 11999 10562 12008
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10520 11762 10548 11999
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11286 10088 11562
rect 10152 11558 10180 11630
rect 10704 11558 10732 12242
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9916 11104 9996 11132
rect 9864 11086 9916 11092
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9600 10526 9720 10554
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9402 9616 9458 9625
rect 9402 9551 9458 9560
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9140 8350 9260 8378
rect 9140 8294 9168 8350
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7750 9168 8230
rect 9128 7744 9180 7750
rect 8942 7712 8998 7721
rect 9128 7686 9180 7692
rect 8942 7647 8998 7656
rect 9140 7449 9168 7686
rect 9126 7440 9182 7449
rect 9126 7375 9182 7384
rect 8942 7304 8998 7313
rect 8942 7239 8944 7248
rect 8996 7239 8998 7248
rect 8944 7210 8996 7216
rect 8956 5370 8984 7210
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 5914 9076 6598
rect 9416 6304 9444 9551
rect 9496 8288 9548 8294
rect 9600 8265 9628 10526
rect 9876 10470 9904 11086
rect 10060 10810 10088 11222
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9956 10736 10008 10742
rect 10152 10690 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10322 11248 10378 11257
rect 10322 11183 10324 11192
rect 10376 11183 10378 11192
rect 10324 11154 10376 11160
rect 9956 10678 10008 10684
rect 9864 10464 9916 10470
rect 9678 10432 9734 10441
rect 9864 10406 9916 10412
rect 9678 10367 9734 10376
rect 9692 10062 9720 10367
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 8362 9720 9998
rect 9784 9178 9812 10066
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9784 8634 9812 9114
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9496 8230 9548 8236
rect 9586 8256 9642 8265
rect 9508 7342 9536 8230
rect 9586 8191 9642 8200
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 7041 9720 7278
rect 9678 7032 9734 7041
rect 9678 6967 9734 6976
rect 9784 6866 9812 7647
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6390 9812 6802
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9232 6276 9444 6304
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 2962 439 3018 448
rect 3146 0 3202 480
rect 3698 0 3754 480
rect 4250 0 4306 480
rect 4802 0 4858 480
rect 5354 0 5410 480
rect 5998 0 6054 480
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8850 0 8906 480
rect 8956 105 8984 3334
rect 9048 1329 9076 4150
rect 9034 1320 9090 1329
rect 9034 1255 9090 1264
rect 9232 610 9260 6276
rect 9310 6216 9366 6225
rect 9310 6151 9366 6160
rect 9324 5914 9352 6151
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5234 9352 5850
rect 9494 5808 9550 5817
rect 9494 5743 9550 5752
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9508 5166 9536 5743
rect 9772 5704 9824 5710
rect 9678 5672 9734 5681
rect 9772 5646 9824 5652
rect 9678 5607 9680 5616
rect 9732 5607 9734 5616
rect 9680 5578 9732 5584
rect 9784 5386 9812 5646
rect 9600 5370 9812 5386
rect 9588 5364 9812 5370
rect 9640 5358 9812 5364
rect 9588 5306 9640 5312
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9416 4554 9444 4966
rect 9600 4826 9628 5306
rect 9876 4826 9904 10406
rect 9968 10130 9996 10678
rect 10060 10662 10180 10690
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 9427 9996 10066
rect 9948 9382 9996 9427
rect 9936 9376 9996 9382
rect 9988 9324 9996 9376
rect 9936 9318 9996 9324
rect 9968 8838 9996 9318
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8090 9996 8774
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9968 7177 9996 7210
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9954 6760 10010 6769
rect 9954 6695 10010 6704
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9968 4758 9996 6695
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9416 3738 9444 4490
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9508 3210 9536 4558
rect 9680 4480 9732 4486
rect 9968 4457 9996 4558
rect 9680 4422 9732 4428
rect 9954 4448 10010 4457
rect 9692 4162 9720 4422
rect 9954 4383 10010 4392
rect 9600 4134 9720 4162
rect 9772 4140 9824 4146
rect 9600 4078 9628 4134
rect 9772 4082 9824 4088
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3505 9720 3878
rect 9678 3496 9734 3505
rect 9678 3431 9734 3440
rect 9508 3194 9720 3210
rect 9508 3188 9732 3194
rect 9508 3182 9680 3188
rect 9680 3130 9732 3136
rect 9494 3088 9550 3097
rect 9494 3023 9550 3032
rect 9508 2922 9536 3023
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9784 2854 9812 4082
rect 9968 3942 9996 4383
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9862 3632 9918 3641
rect 9862 3567 9864 3576
rect 9916 3567 9918 3576
rect 9864 3538 9916 3544
rect 9876 3126 9904 3538
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9772 2848 9824 2854
rect 10060 2802 10088 10662
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10152 9058 10180 9454
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10428 9110 10456 9141
rect 10416 9104 10468 9110
rect 10152 9052 10416 9058
rect 10152 9046 10468 9052
rect 10152 9030 10456 9046
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8838 10272 8910
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10336 8650 10364 8842
rect 10428 8786 10456 9030
rect 10704 8922 10732 11494
rect 10796 10962 10824 12582
rect 10888 11694 10916 12679
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10980 11082 11008 14214
rect 11072 13190 11100 15302
rect 11164 14822 11192 17206
rect 11256 16794 11284 20046
rect 11348 19922 11376 20198
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11348 19514 11376 19858
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11334 19408 11390 19417
rect 11334 19343 11390 19352
rect 11348 19242 11376 19343
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11440 18426 11468 20295
rect 11532 20097 11560 24103
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23662 11744 24006
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11888 23656 11940 23662
rect 11888 23598 11940 23604
rect 11716 23168 11744 23598
rect 11900 23254 11928 23598
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 11796 23180 11848 23186
rect 11716 23140 11796 23168
rect 11716 22642 11744 23140
rect 11796 23122 11848 23128
rect 11900 22778 11928 23190
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 21690 11744 22578
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11612 21480 11664 21486
rect 11612 21422 11664 21428
rect 11624 21049 11652 21422
rect 11610 21040 11666 21049
rect 11610 20975 11666 20984
rect 11716 20466 11744 21626
rect 11808 21350 11836 21966
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 21185 11836 21286
rect 11794 21176 11850 21185
rect 11794 21111 11850 21120
rect 11900 21078 11928 21966
rect 11888 21072 11940 21078
rect 11888 21014 11940 21020
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11518 20088 11574 20097
rect 11518 20023 11574 20032
rect 11716 19990 11744 20402
rect 11704 19984 11756 19990
rect 11704 19926 11756 19932
rect 11610 19408 11666 19417
rect 11610 19343 11666 19352
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11348 17542 11376 18022
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11348 17338 11376 17478
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11348 16114 11376 16594
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11164 14006 11192 14758
rect 11532 14550 11560 14758
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11242 13288 11298 13297
rect 11532 13258 11560 14486
rect 11242 13223 11298 13232
rect 11520 13252 11572 13258
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 13025 11100 13126
rect 11256 13025 11284 13223
rect 11520 13194 11572 13200
rect 11058 13016 11114 13025
rect 11058 12951 11114 12960
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 11060 12640 11112 12646
rect 11058 12608 11060 12617
rect 11112 12608 11114 12617
rect 11058 12543 11114 12552
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11532 12209 11560 12310
rect 11518 12200 11574 12209
rect 11518 12135 11574 12144
rect 11532 11558 11560 12135
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11164 11354 11192 11494
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11532 11150 11560 11494
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11152 11008 11204 11014
rect 10796 10934 11008 10962
rect 11152 10950 11204 10956
rect 10874 10840 10930 10849
rect 10874 10775 10930 10784
rect 10888 10577 10916 10775
rect 10874 10568 10930 10577
rect 10874 10503 10930 10512
rect 10784 10464 10836 10470
rect 10980 10452 11008 10934
rect 10784 10406 10836 10412
rect 10888 10424 11008 10452
rect 11164 10452 11192 10950
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11244 10464 11296 10470
rect 11164 10424 11244 10452
rect 10796 9761 10824 10406
rect 10782 9752 10838 9761
rect 10782 9687 10838 9696
rect 10888 9217 10916 10424
rect 11244 10406 11296 10412
rect 11256 10169 11284 10406
rect 11440 10266 11468 10610
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 10968 9512 11020 9518
rect 11072 9500 11100 9862
rect 11020 9472 11100 9500
rect 10968 9454 11020 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10874 9208 10930 9217
rect 10874 9143 10930 9152
rect 10782 9072 10838 9081
rect 10838 9016 11008 9024
rect 10782 9007 10784 9016
rect 10836 8996 11008 9016
rect 10784 8978 10836 8984
rect 10704 8894 10916 8922
rect 10428 8758 10732 8786
rect 10152 8622 10364 8650
rect 10152 8090 10180 8622
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10704 7954 10732 8758
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10704 7478 10732 7890
rect 10796 7546 10824 7890
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10782 7440 10838 7449
rect 10782 7375 10838 7384
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10690 7168 10746 7177
rect 10152 6186 10180 7142
rect 10289 7100 10585 7120
rect 10690 7103 10746 7112
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10152 5692 10180 6122
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5914 10732 7103
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10232 5704 10284 5710
rect 10152 5664 10232 5692
rect 10232 5646 10284 5652
rect 10244 5370 10272 5646
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10598 5400 10654 5409
rect 10232 5364 10284 5370
rect 10598 5335 10600 5344
rect 10232 5306 10284 5312
rect 10652 5335 10654 5344
rect 10600 5306 10652 5312
rect 10612 5166 10640 5306
rect 10704 5234 10732 5510
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 10152 4282 10180 4694
rect 10704 4622 10732 5170
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3632 10194 3641
rect 10138 3567 10140 3576
rect 10192 3567 10194 3576
rect 10140 3538 10192 3544
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10704 2854 10732 3062
rect 9772 2790 9824 2796
rect 9784 2446 9812 2790
rect 9948 2774 10088 2802
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 9948 2666 9976 2774
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9948 2638 9996 2666
rect 10704 2650 10732 2790
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9220 604 9272 610
rect 9220 546 9272 552
rect 9404 604 9456 610
rect 9404 546 9456 552
rect 9416 480 9444 546
rect 9968 480 9996 2638
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 8942 96 8998 105
rect 8942 31 8998 40
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10060 241 10088 2246
rect 10796 1442 10824 7375
rect 10888 4842 10916 8894
rect 10980 8362 11008 8996
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11072 8265 11100 9318
rect 11164 9110 11192 9862
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 8498 11284 8774
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11058 8256 11114 8265
rect 11058 8191 11114 8200
rect 10968 7948 11020 7954
rect 11072 7936 11100 8191
rect 11020 7908 11100 7936
rect 10968 7890 11020 7896
rect 11348 7410 11376 8298
rect 11624 7546 11652 19343
rect 11888 19168 11940 19174
rect 11886 19136 11888 19145
rect 11940 19136 11942 19145
rect 11886 19071 11942 19080
rect 11702 18728 11758 18737
rect 11702 18663 11758 18672
rect 11716 16522 11744 18663
rect 11794 17096 11850 17105
rect 11794 17031 11796 17040
rect 11848 17031 11850 17040
rect 11796 17002 11848 17008
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 16250 11744 16458
rect 11992 16454 12020 24534
rect 12084 23866 12112 24550
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12176 23633 12204 24686
rect 12162 23624 12218 23633
rect 12072 23588 12124 23594
rect 12162 23559 12218 23568
rect 12072 23530 12124 23536
rect 12084 22545 12112 23530
rect 12162 23080 12218 23089
rect 12162 23015 12218 23024
rect 12176 22778 12204 23015
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12176 22574 12204 22714
rect 12164 22568 12216 22574
rect 12070 22536 12126 22545
rect 12164 22510 12216 22516
rect 12070 22471 12126 22480
rect 12162 22128 12218 22137
rect 12162 22063 12218 22072
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 12084 21146 12112 21927
rect 12176 21690 12204 22063
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12176 19825 12204 21354
rect 12268 20641 12296 27520
rect 12820 27418 12848 27520
rect 12820 27390 13032 27418
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12452 25242 12480 25910
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12544 25362 12572 25842
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12452 25214 12572 25242
rect 12544 22098 12572 25214
rect 12636 24954 12664 26454
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12622 23760 12678 23769
rect 12728 23730 12756 24006
rect 12622 23695 12678 23704
rect 12716 23724 12768 23730
rect 12636 23202 12664 23695
rect 12716 23666 12768 23672
rect 12728 23322 12756 23666
rect 12900 23520 12952 23526
rect 12898 23488 12900 23497
rect 12952 23488 12954 23497
rect 12898 23423 12954 23432
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12636 23174 12756 23202
rect 12624 22704 12676 22710
rect 12622 22672 12624 22681
rect 12676 22672 12678 22681
rect 12622 22607 12678 22616
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12544 21486 12572 22034
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12254 20632 12310 20641
rect 12254 20567 12310 20576
rect 12452 19990 12480 20946
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 20602 12664 20878
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12162 19816 12218 19825
rect 12162 19751 12218 19760
rect 12452 19514 12480 19926
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12176 19174 12204 19246
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18290 12112 18566
rect 12176 18465 12204 19110
rect 12162 18456 12218 18465
rect 12162 18391 12218 18400
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12440 18352 12492 18358
rect 12438 18320 12440 18329
rect 12492 18320 12494 18329
rect 12072 18284 12124 18290
rect 12438 18255 12494 18264
rect 12072 18226 12124 18232
rect 12084 17746 12112 18226
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12084 16794 12112 17682
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 12176 16182 12204 17478
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12254 16824 12310 16833
rect 12254 16759 12256 16768
rect 12308 16759 12310 16768
rect 12348 16788 12400 16794
rect 12256 16730 12308 16736
rect 12348 16730 12400 16736
rect 12360 16250 12388 16730
rect 12452 16697 12480 16934
rect 12544 16794 12572 18362
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12438 16688 12494 16697
rect 12438 16623 12494 16632
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 16522 12572 16594
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12164 16176 12216 16182
rect 11794 16144 11850 16153
rect 11850 16102 11928 16130
rect 12164 16118 12216 16124
rect 11794 16079 11850 16088
rect 11900 15881 11928 16102
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12440 16040 12492 16046
rect 12636 16017 12664 16050
rect 12440 15982 12492 15988
rect 12622 16008 12678 16017
rect 11886 15872 11942 15881
rect 11886 15807 11942 15816
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12986 11744 13330
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11150 11836 11630
rect 11704 11144 11756 11150
rect 11702 11112 11704 11121
rect 11796 11144 11848 11150
rect 11756 11112 11758 11121
rect 11796 11086 11848 11092
rect 11702 11047 11758 11056
rect 11716 9654 11744 11047
rect 11808 10266 11836 11086
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11058 7304 11114 7313
rect 11058 7239 11114 7248
rect 11334 7304 11390 7313
rect 11334 7239 11336 7248
rect 11072 7041 11100 7239
rect 11388 7239 11390 7248
rect 11336 7210 11388 7216
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11058 7032 11114 7041
rect 11058 6967 11114 6976
rect 11072 6730 11100 6967
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5030 11008 6054
rect 11072 5846 11100 6287
rect 11152 6112 11204 6118
rect 11150 6080 11152 6089
rect 11204 6080 11206 6089
rect 11150 6015 11206 6024
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10968 5024 11020 5030
rect 11152 5024 11204 5030
rect 11020 4984 11100 5012
rect 10968 4966 11020 4972
rect 10888 4814 11008 4842
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 2689 10916 3878
rect 10980 2938 11008 4814
rect 11072 3058 11100 4984
rect 11152 4966 11204 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 4078 11284 7142
rect 11716 6905 11744 8434
rect 11702 6896 11758 6905
rect 11702 6831 11758 6840
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5953 11468 6054
rect 11426 5944 11482 5953
rect 11426 5879 11482 5888
rect 11334 5808 11390 5817
rect 11334 5743 11336 5752
rect 11388 5743 11390 5752
rect 11336 5714 11388 5720
rect 11348 4758 11376 5714
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4826 11468 5102
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11164 2990 11192 3470
rect 11152 2984 11204 2990
rect 10980 2910 11100 2938
rect 11152 2926 11204 2932
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10874 2680 10930 2689
rect 10980 2650 11008 2790
rect 10874 2615 10930 2624
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10520 1414 10824 1442
rect 10520 480 10548 1414
rect 11072 480 11100 2910
rect 11256 2802 11284 4014
rect 11348 3738 11376 4082
rect 11532 3942 11560 6598
rect 11624 4060 11652 6598
rect 11716 6458 11744 6831
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11716 4758 11744 6394
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5370 11836 5782
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 4214 11744 4694
rect 11794 4584 11850 4593
rect 11794 4519 11796 4528
rect 11848 4519 11850 4528
rect 11796 4490 11848 4496
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11624 4049 11744 4060
rect 11624 4040 11758 4049
rect 11624 4032 11702 4040
rect 11702 3975 11758 3984
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11348 3398 11376 3674
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 2922 11376 3334
rect 11716 3108 11744 3975
rect 11808 3942 11836 4490
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3505 11836 3878
rect 11794 3496 11850 3505
rect 11794 3431 11850 3440
rect 11900 3380 11928 15807
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11992 13530 12020 13670
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11992 10130 12020 12922
rect 12084 10810 12112 15506
rect 12452 15162 12480 15982
rect 12622 15943 12678 15952
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12544 15094 12572 15438
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14618 12572 14758
rect 12728 14634 12756 23174
rect 12900 22976 12952 22982
rect 12898 22944 12900 22953
rect 12952 22944 12954 22953
rect 12898 22879 12954 22888
rect 13004 21729 13032 27390
rect 13372 25514 13400 27520
rect 13728 26308 13780 26314
rect 13728 26250 13780 26256
rect 13280 25486 13400 25514
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 12990 21720 13046 21729
rect 12990 21655 13046 21664
rect 12808 19168 12860 19174
rect 12806 19136 12808 19145
rect 12860 19136 12862 19145
rect 12806 19071 12862 19080
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 18086 12848 18702
rect 13004 18578 13032 21655
rect 13096 21554 13124 22918
rect 13280 22817 13308 25486
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13372 24954 13400 25298
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13556 24750 13584 25094
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 13556 24313 13584 24686
rect 13648 24614 13676 25298
rect 13740 24954 13768 26250
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13924 24834 13952 27520
rect 14568 27418 14596 27520
rect 14476 27390 14596 27418
rect 13924 24806 14320 24834
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13542 24304 13598 24313
rect 13452 24268 13504 24274
rect 13542 24239 13598 24248
rect 13452 24210 13504 24216
rect 13464 23594 13492 24210
rect 14004 24064 14056 24070
rect 14108 24041 14136 24550
rect 14004 24006 14056 24012
rect 14094 24032 14150 24041
rect 14016 23730 14044 24006
rect 14094 23967 14150 23976
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13740 23610 13768 23666
rect 14016 23610 14044 23666
rect 13452 23588 13504 23594
rect 13740 23582 13860 23610
rect 14016 23582 14136 23610
rect 13452 23530 13504 23536
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13266 22808 13322 22817
rect 13556 22778 13584 23054
rect 13266 22743 13322 22752
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13740 22506 13768 23258
rect 13832 22778 13860 23582
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13740 22234 13768 22442
rect 13924 22438 13952 23190
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13372 21554 13400 22170
rect 13726 22128 13782 22137
rect 13726 22063 13728 22072
rect 13780 22063 13782 22072
rect 13728 22034 13780 22040
rect 13452 22024 13504 22030
rect 13740 22003 13768 22034
rect 13452 21966 13504 21972
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13464 21146 13492 21966
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 21457 13676 21830
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13634 21448 13690 21457
rect 13634 21383 13690 21392
rect 13740 21146 13768 21490
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20942 13860 21286
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 13096 19786 13124 20266
rect 13188 20058 13216 20742
rect 13832 20602 13860 20878
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 20058 13860 20198
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13924 19938 13952 22374
rect 14016 21962 14044 23462
rect 14108 23322 14136 23582
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14108 22574 14136 23054
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 14108 22137 14136 22510
rect 14094 22128 14150 22137
rect 14094 22063 14150 22072
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14004 21956 14056 21962
rect 14004 21898 14056 21904
rect 14016 21690 14044 21898
rect 14108 21690 14136 21966
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14108 21078 14136 21626
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20602 14136 20878
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14108 20210 14136 20538
rect 14200 20262 14228 24686
rect 14292 21185 14320 24806
rect 14278 21176 14334 21185
rect 14278 21111 14334 21120
rect 14476 20890 14504 27390
rect 15120 25242 15148 27520
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 14752 25214 15148 25242
rect 14646 23488 14702 23497
rect 14646 23423 14702 23432
rect 14384 20862 14504 20890
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 13832 19910 13952 19938
rect 14016 20182 14136 20210
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 13096 19378 13124 19722
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 18970 13124 19314
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13648 18970 13676 19178
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13450 18864 13506 18873
rect 13450 18799 13506 18808
rect 13004 18550 13308 18578
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17377 12848 18022
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12806 17368 12862 17377
rect 12806 17303 12862 17312
rect 12912 17270 12940 17478
rect 12900 17264 12952 17270
rect 12820 17212 12900 17218
rect 12820 17206 12952 17212
rect 12820 17190 12940 17206
rect 13004 17202 13032 18158
rect 13174 17912 13230 17921
rect 13174 17847 13230 17856
rect 12820 16590 12848 17190
rect 12912 17141 12940 17190
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13188 17134 13216 17847
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 15706 12848 16526
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12532 14612 12584 14618
rect 12728 14606 12848 14634
rect 12532 14554 12584 14560
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12268 13938 12296 14214
rect 12544 14074 12572 14554
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 14346 12756 14418
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12728 14074 12756 14282
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12176 10985 12204 13738
rect 12268 13462 12296 13874
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12360 13394 12388 13670
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12256 12096 12308 12102
rect 12308 12044 12388 12050
rect 12256 12038 12388 12044
rect 12268 12022 12388 12038
rect 12360 11694 12388 12022
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12254 11384 12310 11393
rect 12254 11319 12310 11328
rect 12162 10976 12218 10985
rect 12162 10911 12218 10920
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12084 10538 12112 10746
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11980 8900 12032 8906
rect 12176 8888 12204 10066
rect 12268 9654 12296 11319
rect 12360 10130 12388 11630
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10606 12572 10950
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12032 8860 12204 8888
rect 11980 8842 12032 8848
rect 11992 8276 12020 8842
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12072 8288 12124 8294
rect 11992 8248 12072 8276
rect 11992 7818 12020 8248
rect 12072 8230 12124 8236
rect 12176 8090 12204 8298
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7342 12020 7754
rect 12072 7744 12124 7750
rect 12070 7712 12072 7721
rect 12124 7712 12126 7721
rect 12070 7647 12126 7656
rect 12084 7449 12112 7647
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12084 6798 12112 7210
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 5914 12020 6598
rect 12084 6254 12112 6734
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12084 3670 12112 5306
rect 12162 4856 12218 4865
rect 12162 4791 12164 4800
rect 12216 4791 12218 4800
rect 12164 4762 12216 4768
rect 12176 3942 12204 4762
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11532 3080 11744 3108
rect 11808 3352 11928 3380
rect 11532 2972 11560 3080
rect 11440 2944 11560 2972
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11164 2774 11284 2802
rect 11164 2553 11192 2774
rect 11440 2650 11468 2944
rect 11808 2666 11836 3352
rect 11992 3194 12020 3538
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12176 3097 12204 3878
rect 12162 3088 12218 3097
rect 11980 3052 12032 3058
rect 12162 3023 12218 3032
rect 11980 2994 12032 3000
rect 11992 2922 12020 2994
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11716 2638 11836 2666
rect 11992 2650 12020 2858
rect 11980 2644 12032 2650
rect 11150 2544 11206 2553
rect 11150 2479 11206 2488
rect 11716 480 11744 2638
rect 11980 2586 12032 2592
rect 11992 2446 12020 2586
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12268 480 12296 7482
rect 12360 5710 12388 9279
rect 12452 9178 12480 10406
rect 12544 9586 12572 10542
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12452 9042 12480 9114
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12452 5658 12480 7890
rect 12532 6928 12584 6934
rect 12530 6896 12532 6905
rect 12584 6896 12586 6905
rect 12530 6831 12586 6840
rect 12360 5370 12388 5646
rect 12452 5630 12572 5658
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5234 12480 5510
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12544 5114 12572 5630
rect 12452 5086 12572 5114
rect 12452 3738 12480 5086
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 3738 12572 4966
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12452 3466 12480 3674
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12636 1850 12664 13942
rect 12728 13258 12756 14010
rect 12820 13530 12848 14606
rect 12912 14278 12940 15506
rect 13004 15366 13032 16050
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 14550 13032 15302
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14414 13032 14486
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 13004 13938 13032 14350
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12986 12756 13194
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12820 12889 12848 13466
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12806 12880 12862 12889
rect 12806 12815 12808 12824
rect 12860 12815 12862 12824
rect 12808 12786 12860 12792
rect 12820 12755 12848 12786
rect 13004 12646 13032 13330
rect 13188 13297 13216 13806
rect 13174 13288 13230 13297
rect 13174 13223 13230 13232
rect 13280 13172 13308 18550
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15026 13400 15846
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13188 13144 13308 13172
rect 12992 12640 13044 12646
rect 12990 12608 12992 12617
rect 13044 12608 13046 12617
rect 12990 12543 13046 12552
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13004 11694 13032 12310
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 12714 10976 12770 10985
rect 12714 10911 12770 10920
rect 12728 5030 12756 10911
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12820 9625 12848 10678
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12898 10296 12954 10305
rect 12898 10231 12954 10240
rect 12912 9897 12940 10231
rect 13004 10130 13032 10610
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12898 9888 12954 9897
rect 12898 9823 12954 9832
rect 12898 9752 12954 9761
rect 12898 9687 12954 9696
rect 12806 9616 12862 9625
rect 12806 9551 12862 9560
rect 12912 9178 12940 9687
rect 13004 9382 13032 10066
rect 12992 9376 13044 9382
rect 12990 9344 12992 9353
rect 13044 9344 13046 9353
rect 12990 9279 13046 9288
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12912 8634 12940 9114
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 8090 12940 8230
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13004 7585 13032 8978
rect 12990 7576 13046 7585
rect 12990 7511 13046 7520
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12990 6080 13046 6089
rect 12820 5914 12848 6054
rect 12990 6015 13046 6024
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12898 5672 12954 5681
rect 12820 5370 12848 5646
rect 12898 5607 12900 5616
rect 12952 5607 12954 5616
rect 12900 5578 12952 5584
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 4146 12940 4422
rect 12900 4140 12952 4146
rect 12820 4100 12900 4128
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12728 2009 12756 3946
rect 12820 3602 12848 4100
rect 12900 4082 12952 4088
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12912 3398 12940 3878
rect 13004 3777 13032 6015
rect 12990 3768 13046 3777
rect 12990 3703 13046 3712
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3097 12940 3334
rect 12898 3088 12954 3097
rect 12898 3023 12954 3032
rect 13188 2582 13216 13144
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11286 13308 12038
rect 13464 11354 13492 18799
rect 13740 17882 13768 18906
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13556 13530 13584 13806
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 12850 13584 13126
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13556 12442 13584 12786
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13556 12170 13584 12378
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13358 11248 13414 11257
rect 13358 11183 13414 11192
rect 13372 11150 13400 11183
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 10810 13584 11086
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13648 10010 13676 17070
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 16114 13768 16390
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13832 15162 13860 19910
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13924 19446 13952 19790
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 14016 19258 14044 20182
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13924 19230 14044 19258
rect 13924 15552 13952 19230
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18834 14044 19110
rect 14108 18873 14136 19858
rect 14292 19378 14320 19926
rect 14384 19446 14412 20862
rect 14568 20602 14596 20878
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14660 20466 14688 23423
rect 14752 20806 14780 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15488 24954 15516 25298
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 15198 24848 15254 24857
rect 15198 24783 15254 24792
rect 15212 24177 15240 24783
rect 15672 24698 15700 27520
rect 16118 24848 16174 24857
rect 16118 24783 16174 24792
rect 15304 24670 15700 24698
rect 15936 24676 15988 24682
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23338 15332 24670
rect 15936 24618 15988 24624
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 24313 15700 24550
rect 15658 24304 15714 24313
rect 15568 24268 15620 24274
rect 15658 24239 15714 24248
rect 15568 24210 15620 24216
rect 15580 23866 15608 24210
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15120 23310 15332 23338
rect 15120 23186 15148 23310
rect 15290 23216 15346 23225
rect 15108 23180 15160 23186
rect 15290 23151 15292 23160
rect 15108 23122 15160 23128
rect 15344 23151 15346 23160
rect 15292 23122 15344 23128
rect 15396 23118 15424 23462
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22778 15424 23054
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15752 22568 15804 22574
rect 15752 22510 15804 22516
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14830 21176 14886 21185
rect 14830 21111 14886 21120
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 14094 18864 14150 18873
rect 14004 18828 14056 18834
rect 14094 18799 14150 18808
rect 14004 18770 14056 18776
rect 14016 17882 14044 18770
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14108 18426 14136 18702
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14200 17882 14228 19178
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14108 16454 14136 17070
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14200 15706 14228 15914
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 13924 15524 14044 15552
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13924 15201 13952 15370
rect 13910 15192 13966 15201
rect 13820 15156 13872 15162
rect 13910 15127 13966 15136
rect 13820 15098 13872 15104
rect 13832 10690 13860 15098
rect 14016 13841 14044 15524
rect 14186 14784 14242 14793
rect 14186 14719 14242 14728
rect 14002 13832 14058 13841
rect 14002 13767 14058 13776
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12102 13952 13126
rect 13912 12096 13964 12102
rect 13910 12064 13912 12073
rect 13964 12064 13966 12073
rect 13910 11999 13966 12008
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13740 10662 13860 10690
rect 13740 10305 13768 10662
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 13726 10296 13782 10305
rect 13726 10231 13782 10240
rect 13740 10198 13768 10231
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13372 9982 13676 10010
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13280 6254 13308 8502
rect 13372 7954 13400 9982
rect 13832 9926 13860 10474
rect 13452 9920 13504 9926
rect 13820 9920 13872 9926
rect 13452 9862 13504 9868
rect 13648 9868 13820 9874
rect 13648 9862 13872 9868
rect 13464 9722 13492 9862
rect 13648 9846 13860 9862
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13464 8974 13492 9658
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 9110 13584 9454
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13464 7886 13492 8910
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 7880 13504 7886
rect 13372 7828 13452 7834
rect 13372 7822 13504 7828
rect 13372 7806 13492 7822
rect 13372 7546 13400 7806
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7274 13492 7686
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5914 13308 6190
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13372 5370 13400 5714
rect 13464 5710 13492 7210
rect 13556 7002 13584 8298
rect 13648 8090 13676 9846
rect 13818 8936 13874 8945
rect 13818 8871 13874 8880
rect 13726 8120 13782 8129
rect 13636 8084 13688 8090
rect 13726 8055 13728 8064
rect 13636 8026 13688 8032
rect 13780 8055 13782 8064
rect 13728 8026 13780 8032
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13556 6118 13584 6938
rect 13648 6662 13676 7890
rect 13740 7002 13768 8026
rect 13832 7954 13860 8871
rect 13924 8090 13952 11766
rect 14016 11218 14044 13767
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14108 11898 14136 12650
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14108 11150 14136 11834
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13556 5234 13584 6054
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13188 2310 13216 2518
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13004 2009 13032 2246
rect 12714 2000 12770 2009
rect 12714 1935 12770 1944
rect 12990 2000 13046 2009
rect 12990 1935 13046 1944
rect 12636 1822 12848 1850
rect 12820 480 12848 1822
rect 13372 480 13400 4966
rect 13556 4826 13584 5170
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13648 4078 13676 5578
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5250 13860 5510
rect 13740 5222 13860 5250
rect 13740 5166 13768 5222
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13726 4992 13782 5001
rect 13726 4927 13782 4936
rect 13740 4826 13768 4927
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13818 4720 13874 4729
rect 13818 4655 13874 4664
rect 13832 4622 13860 4655
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13726 4312 13782 4321
rect 13726 4247 13782 4256
rect 13636 4072 13688 4078
rect 13740 4049 13768 4247
rect 13636 4014 13688 4020
rect 13726 4040 13782 4049
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3233 13584 3878
rect 13648 3738 13676 4014
rect 13832 4010 13860 4558
rect 13726 3975 13782 3984
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13542 3224 13598 3233
rect 13542 3159 13598 3168
rect 13450 2680 13506 2689
rect 13450 2615 13452 2624
rect 13504 2615 13506 2624
rect 13452 2586 13504 2592
rect 13648 2553 13676 3470
rect 13740 3194 13768 3606
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13634 2544 13690 2553
rect 13634 2479 13690 2488
rect 13740 2446 13768 2790
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13924 480 13952 7686
rect 14016 5234 14044 10950
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10305 14136 10406
rect 14094 10296 14150 10305
rect 14094 10231 14150 10240
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14108 9489 14136 10134
rect 14094 9480 14150 9489
rect 14094 9415 14150 9424
rect 14200 9194 14228 14719
rect 14292 12594 14320 19314
rect 14384 12730 14412 19382
rect 14476 19378 14504 19654
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14568 18154 14596 19994
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14660 18698 14688 19314
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14660 18222 14688 18634
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14568 17882 14596 18090
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14476 14958 14504 15098
rect 14568 15026 14596 15506
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14464 14952 14516 14958
rect 14660 14906 14688 18022
rect 14464 14894 14516 14900
rect 14568 14878 14688 14906
rect 14568 12782 14596 14878
rect 14646 14512 14702 14521
rect 14646 14447 14702 14456
rect 14556 12776 14608 12782
rect 14384 12702 14504 12730
rect 14556 12718 14608 12724
rect 14292 12566 14412 12594
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11286 14320 12038
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14384 11121 14412 12566
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10470 14320 10950
rect 14370 10704 14426 10713
rect 14370 10639 14426 10648
rect 14384 10606 14412 10639
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14108 9166 14228 9194
rect 14108 7750 14136 9166
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14200 8498 14228 9046
rect 14292 8906 14320 10406
rect 14476 10112 14504 12702
rect 14660 12442 14688 14447
rect 14752 12866 14780 20742
rect 14844 20482 14872 21111
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14844 20454 14964 20482
rect 14830 20088 14886 20097
rect 14830 20023 14886 20032
rect 14844 18086 14872 20023
rect 14936 19802 14964 20454
rect 15200 19916 15252 19922
rect 15304 19904 15332 22442
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15580 21554 15608 22034
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15384 21140 15436 21146
rect 15384 21082 15436 21088
rect 15396 20534 15424 21082
rect 15580 20874 15608 21490
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20602 15608 20810
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15396 20074 15424 20470
rect 15396 20058 15516 20074
rect 15384 20052 15516 20058
rect 15436 20046 15516 20052
rect 15384 19994 15436 20000
rect 15252 19876 15332 19904
rect 15384 19916 15436 19922
rect 15200 19858 15252 19864
rect 15384 19858 15436 19864
rect 14936 19774 15332 19802
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14844 16794 14872 17682
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16017 15332 19774
rect 15396 19174 15424 19858
rect 15488 19514 15516 20046
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15568 19304 15620 19310
rect 15566 19272 15568 19281
rect 15620 19272 15622 19281
rect 15566 19207 15622 19216
rect 15384 19168 15436 19174
rect 15672 19156 15700 21286
rect 15764 19825 15792 22510
rect 15948 21350 15976 24618
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 16040 22642 16068 23462
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15750 19816 15806 19825
rect 15750 19751 15806 19760
rect 15856 19378 15884 20334
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15384 19110 15436 19116
rect 15580 19128 15700 19156
rect 15396 18426 15424 19110
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15382 16688 15438 16697
rect 15488 16658 15516 16934
rect 15382 16623 15438 16632
rect 15476 16652 15528 16658
rect 15290 16008 15346 16017
rect 15290 15943 15346 15952
rect 15396 15706 15424 16623
rect 15476 16594 15528 16600
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15396 14958 15424 15302
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15396 14414 15424 14894
rect 15384 14408 15436 14414
rect 15014 14376 15070 14385
rect 14844 14334 15014 14362
rect 14844 12986 14872 14334
rect 15384 14350 15436 14356
rect 15014 14311 15070 14320
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 13870 15424 14350
rect 15488 14074 15516 16594
rect 15580 15570 15608 19128
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15672 18154 15700 18770
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15764 18222 15792 18702
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 14618 15608 15370
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15580 13002 15608 14554
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15488 12974 15608 13002
rect 14752 12838 14872 12866
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14556 12232 14608 12238
rect 14752 12186 14780 12718
rect 14556 12174 14608 12180
rect 14568 11898 14596 12174
rect 14660 12158 14780 12186
rect 14660 11898 14688 12158
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14646 11792 14702 11801
rect 14646 11727 14702 11736
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14384 10084 14504 10112
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14384 8537 14412 10084
rect 14462 10024 14518 10033
rect 14462 9959 14518 9968
rect 14370 8528 14426 8537
rect 14188 8492 14240 8498
rect 14370 8463 14426 8472
rect 14188 8434 14240 8440
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 6186 14228 7686
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 5710 14136 6054
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14200 5574 14228 6122
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14096 5160 14148 5166
rect 14002 5128 14058 5137
rect 14096 5102 14148 5108
rect 14002 5063 14058 5072
rect 14016 4826 14044 5063
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14016 4457 14044 4762
rect 14002 4448 14058 4457
rect 14002 4383 14058 4392
rect 14016 4282 14044 4383
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14016 2650 14044 3538
rect 14108 2689 14136 5102
rect 14200 4554 14228 5510
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14200 4078 14228 4490
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14200 2922 14228 4014
rect 14292 3534 14320 4558
rect 14384 4486 14412 8026
rect 14476 7392 14504 9959
rect 14568 9722 14596 10610
rect 14660 10198 14688 11727
rect 14752 11354 14780 12038
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14738 11112 14794 11121
rect 14738 11047 14794 11056
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14568 8634 14596 9658
rect 14648 8832 14700 8838
rect 14646 8800 14648 8809
rect 14700 8800 14702 8809
rect 14646 8735 14702 8744
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14568 8362 14596 8570
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14476 7364 14596 7392
rect 14462 7304 14518 7313
rect 14462 7239 14518 7248
rect 14476 7206 14504 7239
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14384 3398 14412 3946
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14384 2854 14412 3334
rect 14476 3074 14504 6734
rect 14568 5658 14596 7364
rect 14660 5778 14688 7754
rect 14752 6798 14780 11047
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 5914 14780 6598
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14738 5808 14794 5817
rect 14648 5772 14700 5778
rect 14738 5743 14794 5752
rect 14648 5714 14700 5720
rect 14568 5630 14688 5658
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14568 3369 14596 3538
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14476 3046 14596 3074
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14094 2680 14150 2689
rect 14004 2644 14056 2650
rect 14094 2615 14150 2624
rect 14004 2586 14056 2592
rect 14568 480 14596 3046
rect 14660 2666 14688 5630
rect 14752 4826 14780 5743
rect 14844 5166 14872 12838
rect 15488 12617 15516 12974
rect 15566 12880 15622 12889
rect 15566 12815 15568 12824
rect 15620 12815 15622 12824
rect 15568 12786 15620 12792
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15198 11656 15254 11665
rect 15198 11591 15200 11600
rect 15252 11591 15254 11600
rect 15200 11562 15252 11568
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11098 15148 11494
rect 15304 11257 15332 12038
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15120 11070 15332 11098
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15200 10600 15252 10606
rect 15014 10568 15070 10577
rect 15014 10503 15016 10512
rect 15068 10503 15070 10512
rect 15198 10568 15200 10577
rect 15252 10568 15254 10577
rect 15198 10503 15254 10512
rect 15016 10474 15068 10480
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9382 15332 11070
rect 15396 10810 15424 11154
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15396 10606 15424 10746
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9042 15332 9318
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15396 8974 15424 9998
rect 15488 9654 15516 11562
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10470 15608 11154
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8480 15332 8774
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15212 8452 15332 8480
rect 15212 8129 15240 8452
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15198 8120 15254 8129
rect 15304 8090 15332 8298
rect 15198 8055 15254 8064
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6730 15240 7142
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6186 15332 6734
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5234 15424 8502
rect 15580 7857 15608 10066
rect 15566 7848 15622 7857
rect 15566 7783 15622 7792
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15488 6458 15516 7414
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14936 4690 14964 5170
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14752 3194 14780 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4078 15332 4762
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14752 2922 14780 3130
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14660 2638 14872 2666
rect 15120 2650 15148 3062
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 14660 2281 14688 2518
rect 14646 2272 14702 2281
rect 14646 2207 14702 2216
rect 14844 1442 14872 2638
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15396 2417 15424 4966
rect 15488 3369 15516 6054
rect 15580 5914 15608 6598
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15568 5092 15620 5098
rect 15568 5034 15620 5040
rect 15580 3738 15608 5034
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15474 3360 15530 3369
rect 15474 3295 15530 3304
rect 15488 3194 15516 3295
rect 15476 3188 15528 3194
rect 15528 3148 15608 3176
rect 15476 3130 15528 3136
rect 15474 3088 15530 3097
rect 15474 3023 15530 3032
rect 15488 2650 15516 3023
rect 15580 2990 15608 3148
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15382 2408 15438 2417
rect 15382 2343 15438 2352
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1414 15148 1442
rect 15120 480 15148 1414
rect 15672 480 15700 18090
rect 15764 16794 15792 18158
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15856 16998 15884 17682
rect 15934 17368 15990 17377
rect 15934 17303 15990 17312
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15856 16590 15884 16934
rect 15948 16726 15976 17303
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15764 15978 15792 16526
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15948 16182 15976 16662
rect 16040 16250 16068 22374
rect 16132 20602 16160 24783
rect 16224 24410 16252 27520
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16210 24168 16266 24177
rect 16210 24103 16266 24112
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16224 17218 16252 24103
rect 16684 23526 16712 24210
rect 16776 23866 16804 27520
rect 17420 24857 17448 27520
rect 17406 24848 17462 24857
rect 17406 24783 17462 24792
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17052 24177 17080 24550
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17038 24168 17094 24177
rect 17038 24103 17094 24112
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 17512 23526 17540 24210
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 16486 23216 16542 23225
rect 16304 23180 16356 23186
rect 16486 23151 16542 23160
rect 16304 23122 16356 23128
rect 16316 22438 16344 23122
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16316 19145 16344 20878
rect 16408 20806 16436 21286
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16302 19136 16358 19145
rect 16302 19071 16358 19080
rect 16500 18850 16528 23151
rect 16684 21486 16712 23462
rect 17512 23254 17540 23462
rect 17500 23248 17552 23254
rect 17500 23190 17552 23196
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16762 21448 16818 21457
rect 16762 21383 16818 21392
rect 16670 20496 16726 20505
rect 16670 20431 16726 20440
rect 16684 20058 16712 20431
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16408 18822 16528 18850
rect 16302 17640 16358 17649
rect 16302 17575 16358 17584
rect 16132 17190 16252 17218
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15948 15881 15976 16118
rect 15934 15872 15990 15881
rect 15934 15807 15990 15816
rect 15750 15736 15806 15745
rect 15750 15671 15806 15680
rect 15764 14226 15792 15671
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14385 15884 15438
rect 15948 14822 15976 15506
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15842 14376 15898 14385
rect 15842 14311 15844 14320
rect 15896 14311 15898 14320
rect 15844 14282 15896 14288
rect 15764 14198 15884 14226
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 12986 15792 13330
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15856 11937 15884 14198
rect 15842 11928 15898 11937
rect 15842 11863 15898 11872
rect 15842 11792 15898 11801
rect 15842 11727 15898 11736
rect 15856 11150 15884 11727
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15844 10056 15896 10062
rect 15948 10033 15976 14758
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12986 16068 13262
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 11898 16068 12922
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16132 11098 16160 17190
rect 16316 17082 16344 17575
rect 16040 11070 16160 11098
rect 16224 17054 16344 17082
rect 16224 11082 16252 17054
rect 16408 16810 16436 18822
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18086 16528 18702
rect 16488 18080 16540 18086
rect 16540 18028 16620 18034
rect 16488 18022 16620 18028
rect 16500 18006 16620 18022
rect 16592 17882 16620 18006
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16316 16782 16436 16810
rect 16316 16561 16344 16782
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16408 15910 16436 16662
rect 16592 16232 16620 16934
rect 16684 16833 16712 17070
rect 16776 16998 16804 21383
rect 17788 21321 17816 24550
rect 17972 24154 18000 27520
rect 18524 24410 18552 27520
rect 18786 24712 18842 24721
rect 18786 24647 18842 24656
rect 18800 24410 18828 24647
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 17880 24138 18000 24154
rect 17868 24132 18000 24138
rect 17920 24126 18000 24132
rect 17868 24074 17920 24080
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17880 22506 17908 23122
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 17774 21312 17830 21321
rect 17696 21270 17774 21298
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16670 16824 16726 16833
rect 16670 16759 16672 16768
rect 16724 16759 16726 16768
rect 16672 16730 16724 16736
rect 16868 16658 16896 17138
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17052 16250 17080 16526
rect 17040 16244 17092 16250
rect 16592 16204 16712 16232
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16316 14278 16344 14826
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 13326 16344 14214
rect 16408 13530 16436 15846
rect 16500 15706 16528 15846
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16488 15360 16540 15366
rect 16592 15314 16620 16050
rect 16684 15638 16712 16204
rect 17040 16186 17092 16192
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 16540 15308 16620 15314
rect 16488 15302 16620 15308
rect 16500 15286 16620 15302
rect 16592 14550 16620 15286
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 13954 16528 14350
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 14074 16896 14214
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16500 13926 16620 13954
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12442 16344 13262
rect 16500 12918 16528 13806
rect 16592 13462 16620 13926
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16212 11076 16264 11082
rect 16040 10198 16068 11070
rect 16212 11018 16264 11024
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16210 10976 16266 10985
rect 16132 10713 16160 10950
rect 16210 10911 16266 10920
rect 16118 10704 16174 10713
rect 16118 10639 16120 10648
rect 16172 10639 16174 10648
rect 16120 10610 16172 10616
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15844 9998 15896 10004
rect 15934 10024 15990 10033
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 7410 15792 9318
rect 15856 8945 15884 9998
rect 15934 9959 15990 9968
rect 15934 9344 15990 9353
rect 15934 9279 15990 9288
rect 15948 8974 15976 9279
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15936 8968 15988 8974
rect 15842 8936 15898 8945
rect 15936 8910 15988 8916
rect 15842 8871 15898 8880
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 7886 15884 8774
rect 15948 8090 15976 8910
rect 16040 8566 16068 8978
rect 16028 8560 16080 8566
rect 16026 8528 16028 8537
rect 16080 8528 16082 8537
rect 16026 8463 16082 8472
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15844 7880 15896 7886
rect 15842 7848 15844 7857
rect 15896 7848 15898 7857
rect 15842 7783 15898 7792
rect 16132 7732 16160 10474
rect 15856 7704 16160 7732
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15856 7290 15884 7704
rect 16224 7562 16252 10911
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9586 16344 9862
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9178 16344 9522
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 15764 7262 15884 7290
rect 15948 7534 16252 7562
rect 15764 5250 15792 7262
rect 15948 6118 15976 7534
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6934 16160 7346
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16316 6746 16344 9114
rect 16408 8634 16436 12854
rect 16500 11898 16528 12854
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16684 11558 16712 12310
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16592 10962 16620 11222
rect 16684 11121 16712 11494
rect 16776 11286 16804 13194
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16592 10934 16712 10962
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9636 16528 10066
rect 16580 9648 16632 9654
rect 16500 9608 16580 9636
rect 16580 9590 16632 9596
rect 16684 9382 16712 10934
rect 16776 10266 16804 11222
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16960 9722 16988 15914
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17512 15570 17540 15846
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 14890 17448 15438
rect 17696 15162 17724 21270
rect 17774 21247 17830 21256
rect 18064 19961 18092 23598
rect 18156 23594 18184 24210
rect 19076 23866 19104 27520
rect 19628 25684 19656 27520
rect 19536 25656 19656 25684
rect 19536 23866 19564 25656
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19982 24848 20038 24857
rect 19982 24783 20038 24792
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19996 24410 20024 24783
rect 20272 24721 20300 27520
rect 20258 24712 20314 24721
rect 20258 24647 20314 24656
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 18050 19952 18106 19961
rect 18050 19887 18106 19896
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15706 17816 15846
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15450 17908 15506
rect 17880 15422 18000 15450
rect 17972 15162 18000 15422
rect 18156 15366 18184 23530
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17696 14890 17724 15098
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17132 14816 17184 14822
rect 17696 14793 17724 14826
rect 17132 14758 17184 14764
rect 17682 14784 17738 14793
rect 17144 14550 17172 14758
rect 17682 14719 17738 14728
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17144 14074 17172 14486
rect 17972 14278 18000 14894
rect 18524 14822 18552 15302
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17592 13456 17644 13462
rect 17406 13424 17462 13433
rect 17406 13359 17462 13368
rect 17590 13424 17592 13433
rect 17644 13424 17646 13433
rect 17590 13359 17646 13368
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12782 17172 13262
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 11898 17356 12378
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17328 11354 17356 11834
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17328 10810 17356 11290
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16408 8430 16436 8570
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16500 8362 16528 8774
rect 16960 8498 16988 9114
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 7546 16436 8230
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16408 7342 16436 7482
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16684 7206 16712 7958
rect 17420 7546 17448 13359
rect 17880 12238 17908 14214
rect 17972 13802 18000 14214
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17500 12232 17552 12238
rect 17498 12200 17500 12209
rect 17868 12232 17920 12238
rect 17552 12200 17554 12209
rect 17868 12174 17920 12180
rect 17498 12135 17554 12144
rect 17512 11898 17540 12135
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17512 10674 17540 11086
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17604 10470 17632 11154
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 18326 10432 18382 10441
rect 17604 9994 17632 10406
rect 18326 10367 18382 10376
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17880 9382 17908 10202
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17512 8838 17540 9318
rect 17880 8838 17908 9318
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17512 8430 17540 8774
rect 17500 8424 17552 8430
rect 17498 8392 17500 8401
rect 17552 8392 17554 8401
rect 17880 8362 17908 8774
rect 17498 8327 17554 8336
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17590 8256 17646 8265
rect 17590 8191 17646 8200
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16224 6718 16344 6746
rect 16224 6254 16252 6718
rect 16684 6662 16712 7142
rect 16304 6656 16356 6662
rect 16672 6656 16724 6662
rect 16356 6604 16436 6610
rect 16304 6598 16436 6604
rect 16672 6598 16724 6604
rect 16316 6582 16436 6598
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15856 5370 15884 5646
rect 15948 5370 15976 5850
rect 16040 5794 16068 6122
rect 16118 5944 16174 5953
rect 16302 5944 16358 5953
rect 16174 5902 16252 5930
rect 16118 5879 16174 5888
rect 16040 5766 16160 5794
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15764 5222 15884 5250
rect 15856 2281 15884 5222
rect 16040 3738 16068 5578
rect 16132 4826 16160 5766
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16132 3942 16160 4626
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15948 3126 15976 3606
rect 16040 3194 16068 3674
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16132 3058 16160 3878
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16026 2544 16082 2553
rect 16026 2479 16082 2488
rect 16040 2446 16068 2479
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15842 2272 15898 2281
rect 15842 2207 15898 2216
rect 15856 785 15884 2207
rect 15842 776 15898 785
rect 15842 711 15898 720
rect 16224 480 16252 5902
rect 16302 5879 16358 5888
rect 16316 5574 16344 5879
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16408 5030 16436 6582
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16500 5234 16528 5850
rect 16684 5710 16712 6598
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16776 5914 16804 6394
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16592 5098 16620 5578
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 17328 5030 17356 5646
rect 17604 5642 17632 8191
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 7342 17816 7822
rect 17776 7336 17828 7342
rect 17774 7304 17776 7313
rect 17828 7304 17830 7313
rect 17774 7239 17830 7248
rect 17788 6458 17816 7239
rect 17880 6905 17908 8298
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7410 18000 7686
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17972 7041 18000 7346
rect 18064 7342 18092 9590
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 7449 18276 9522
rect 18234 7440 18290 7449
rect 18234 7375 18290 7384
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18052 7200 18104 7206
rect 18050 7168 18052 7177
rect 18104 7168 18106 7177
rect 18050 7103 18106 7112
rect 17958 7032 18014 7041
rect 17958 6967 18014 6976
rect 17866 6896 17922 6905
rect 17866 6831 17922 6840
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 18050 6216 18106 6225
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17604 5234 17632 5578
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 16396 5024 16448 5030
rect 16394 4992 16396 5001
rect 17316 5024 17368 5030
rect 16448 4992 16450 5001
rect 17316 4966 17368 4972
rect 16394 4927 16450 4936
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16408 3534 16436 4762
rect 17328 4729 17356 4966
rect 17604 4826 17632 5170
rect 17696 5030 17724 5714
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17696 4865 17724 4966
rect 17682 4856 17738 4865
rect 17592 4820 17644 4826
rect 17880 4826 17908 6190
rect 17960 6180 18012 6186
rect 18050 6151 18106 6160
rect 17960 6122 18012 6128
rect 17972 5370 18000 6122
rect 18064 6118 18092 6151
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18248 5846 18276 7278
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18248 5166 18276 5782
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 17682 4791 17738 4800
rect 17868 4820 17920 4826
rect 17592 4762 17644 4768
rect 17868 4762 17920 4768
rect 18248 4729 18276 5102
rect 17314 4720 17370 4729
rect 18234 4720 18290 4729
rect 17314 4655 17370 4664
rect 17960 4684 18012 4690
rect 18234 4655 18290 4664
rect 17960 4626 18012 4632
rect 17774 4584 17830 4593
rect 17972 4570 18000 4626
rect 17830 4542 18000 4570
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 17774 4519 17830 4528
rect 16854 4312 16910 4321
rect 16854 4247 16910 4256
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3670 16620 4014
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3777 16804 3946
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 2825 16620 3334
rect 16578 2816 16634 2825
rect 16578 2751 16634 2760
rect 16302 2544 16358 2553
rect 16302 2479 16304 2488
rect 16356 2479 16358 2488
rect 16304 2450 16356 2456
rect 16868 1170 16896 4247
rect 17498 4176 17554 4185
rect 17788 4146 17816 4519
rect 18248 4214 18276 4558
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 17498 4111 17554 4120
rect 17776 4140 17828 4146
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 17144 3738 17172 3975
rect 17512 3738 17540 4111
rect 17776 4082 17828 4088
rect 18052 4072 18104 4078
rect 18248 4049 18276 4150
rect 18052 4014 18104 4020
rect 18234 4040 18290 4049
rect 17958 3768 18014 3777
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17500 3732 17552 3738
rect 17958 3703 17960 3712
rect 17500 3674 17552 3680
rect 18012 3703 18014 3712
rect 17960 3674 18012 3680
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17420 3058 17448 3538
rect 17512 3194 17540 3674
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17604 3233 17632 3538
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17590 3224 17646 3233
rect 17500 3188 17552 3194
rect 17590 3159 17646 3168
rect 17500 3130 17552 3136
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17604 2922 17632 3159
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17696 2825 17724 3470
rect 17682 2816 17738 2825
rect 17682 2751 17738 2760
rect 17038 2680 17094 2689
rect 17038 2615 17094 2624
rect 17052 2514 17080 2615
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17696 2446 17724 2751
rect 17958 2680 18014 2689
rect 17958 2615 17960 2624
rect 18012 2615 18014 2624
rect 17960 2586 18012 2592
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17236 2009 17264 2246
rect 17222 2000 17278 2009
rect 17222 1935 17278 1944
rect 18064 1873 18092 4014
rect 18144 4004 18196 4010
rect 18234 3975 18290 3984
rect 18144 3946 18196 3952
rect 17406 1864 17462 1873
rect 17406 1799 17462 1808
rect 18050 1864 18106 1873
rect 18050 1799 18106 1808
rect 16776 1142 16896 1170
rect 16776 480 16804 1142
rect 17420 480 17448 1799
rect 17958 1728 18014 1737
rect 17958 1663 18014 1672
rect 17972 480 18000 1663
rect 18156 649 18184 3946
rect 18340 3942 18368 10367
rect 18418 9752 18474 9761
rect 18524 9722 18552 14758
rect 18616 12442 18644 18119
rect 19076 18057 19104 23598
rect 20088 23526 20116 24210
rect 20442 23896 20498 23905
rect 20442 23831 20444 23840
rect 20496 23831 20498 23840
rect 20444 23802 20496 23808
rect 20260 23656 20312 23662
rect 20824 23610 20852 27520
rect 21376 24857 21404 27520
rect 21362 24848 21418 24857
rect 21362 24783 21418 24792
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20916 23769 20944 24210
rect 21546 24032 21602 24041
rect 21546 23967 21602 23976
rect 21560 23866 21588 23967
rect 21928 23905 21956 27520
rect 22480 24562 22508 27520
rect 22020 24534 22508 24562
rect 22020 24410 22048 24534
rect 22190 24440 22246 24449
rect 22008 24404 22060 24410
rect 22190 24375 22192 24384
rect 22008 24346 22060 24352
rect 22244 24375 22246 24384
rect 22192 24346 22244 24352
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 21914 23896 21970 23905
rect 21548 23860 21600 23866
rect 21914 23831 21970 23840
rect 21548 23802 21600 23808
rect 20902 23760 20958 23769
rect 20902 23695 20904 23704
rect 20956 23695 20958 23704
rect 20904 23666 20956 23672
rect 20260 23598 20312 23604
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19168 22778 19196 23122
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20088 18193 20116 23462
rect 20272 22982 20300 23598
rect 20640 23582 20852 23610
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20640 23322 20668 23582
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 21100 22982 21128 23598
rect 22020 23526 22048 24210
rect 23124 24041 23152 27520
rect 23676 24698 23704 27520
rect 23400 24670 23704 24698
rect 23110 24032 23166 24041
rect 23110 23967 23166 23976
rect 23400 23866 23428 24670
rect 24228 24449 24256 27520
rect 24780 25226 24808 27520
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24440 24270 24449
rect 24214 24375 24270 24384
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 25332 23866 25360 27520
rect 25976 24177 26004 27520
rect 26528 25158 26556 27520
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 27080 24313 27108 27520
rect 27066 24304 27122 24313
rect 27066 24239 27122 24248
rect 25962 24168 26018 24177
rect 25962 24103 26018 24112
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 20074 18184 20130 18193
rect 20074 18119 20130 18128
rect 19062 18048 19118 18057
rect 19062 17983 19118 17992
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20272 16697 20300 22918
rect 20258 16688 20314 16697
rect 20258 16623 20314 16632
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 21100 15638 21128 22918
rect 22020 19417 22048 23462
rect 22374 23216 22430 23225
rect 22374 23151 22376 23160
rect 22428 23151 22430 23160
rect 22376 23122 22428 23128
rect 22388 22778 22416 23122
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22006 19408 22062 19417
rect 22006 19343 22062 19352
rect 22480 17377 22508 23598
rect 23492 23338 23520 23598
rect 23400 23310 23520 23338
rect 23570 23352 23626 23361
rect 23400 23254 23428 23310
rect 23570 23287 23626 23296
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23584 21593 23612 23287
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 23570 21584 23626 21593
rect 23570 21519 23626 21528
rect 27632 21457 27660 27520
rect 27618 21448 27674 21457
rect 27618 21383 27674 21392
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 22466 17368 22522 17377
rect 24289 17360 24585 17380
rect 22466 17303 22522 17312
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 21088 15632 21140 15638
rect 20902 15600 20958 15609
rect 21088 15574 21140 15580
rect 20902 15535 20904 15544
rect 20956 15535 20958 15544
rect 20904 15506 20956 15512
rect 20916 15162 20944 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19352 14074 19380 14855
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 24674 13968 24730 13977
rect 24674 13903 24730 13912
rect 24688 13870 24716 13903
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24412 13462 24440 13806
rect 24400 13456 24452 13462
rect 24398 13424 24400 13433
rect 24452 13424 24454 13433
rect 24398 13359 24454 13368
rect 24122 13288 24178 13297
rect 24122 13223 24178 13232
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18694 12336 18750 12345
rect 18694 12271 18750 12280
rect 18418 9687 18474 9696
rect 18512 9716 18564 9722
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18432 3194 18460 9687
rect 18512 9658 18564 9664
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 7342 18552 7686
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18616 7206 18644 7482
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 18142 640 18198 649
rect 18142 575 18198 584
rect 18248 513 18276 2858
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 1193 18368 2246
rect 18326 1184 18382 1193
rect 18326 1119 18382 1128
rect 18234 504 18290 513
rect 10046 232 10102 241
rect 10046 167 10102 176
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17406 0 17462 480
rect 17958 0 18014 480
rect 18524 480 18552 6598
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18616 5710 18644 6258
rect 18708 5846 18736 12271
rect 20350 11928 20406 11937
rect 20350 11863 20406 11872
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18786 10568 18842 10577
rect 18786 10503 18842 10512
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18708 5166 18736 5782
rect 18800 5522 18828 10503
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19062 9480 19118 9489
rect 19062 9415 19118 9424
rect 18972 8016 19024 8022
rect 18878 7984 18934 7993
rect 18972 7958 19024 7964
rect 18878 7919 18880 7928
rect 18932 7919 18934 7928
rect 18880 7890 18932 7896
rect 18892 7002 18920 7890
rect 18984 7546 19012 7958
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18878 5808 18934 5817
rect 18878 5743 18934 5752
rect 18892 5642 18920 5743
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18800 5494 18920 5522
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 4593 18736 5102
rect 18694 4584 18750 4593
rect 18694 4519 18750 4528
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18800 4078 18828 4422
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18892 3466 18920 5494
rect 18972 3664 19024 3670
rect 19076 3652 19104 9415
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19522 8392 19578 8401
rect 19522 8327 19578 8336
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6186 19196 6734
rect 19444 6458 19472 6802
rect 19536 6730 19564 8327
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20258 6896 20314 6905
rect 20258 6831 20314 6840
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 20272 6662 20300 6831
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19156 6180 19208 6186
rect 19156 6122 19208 6128
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19168 4826 19196 5646
rect 19260 5370 19288 5714
rect 19352 5370 19380 5850
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19260 5137 19288 5306
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19246 5128 19302 5137
rect 19246 5063 19302 5072
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19352 4282 19380 5170
rect 19444 4758 19472 6394
rect 20272 6118 20300 6598
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19522 5808 19578 5817
rect 19522 5743 19578 5752
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19536 4690 19564 5743
rect 20258 5672 20314 5681
rect 20258 5607 20314 5616
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19536 4282 19564 4626
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19024 3624 19104 3652
rect 18972 3606 19024 3612
rect 19260 3534 19288 4082
rect 19996 4078 20024 5510
rect 20074 5264 20130 5273
rect 20074 5199 20130 5208
rect 20088 4826 20116 5199
rect 20272 5166 20300 5607
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20076 4820 20128 4826
rect 20128 4780 20208 4808
rect 20076 4762 20128 4768
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19248 3528 19300 3534
rect 19062 3496 19118 3505
rect 18880 3460 18932 3466
rect 19248 3470 19300 3476
rect 19062 3431 19118 3440
rect 18880 3402 18932 3408
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18708 2514 18736 2790
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18708 1601 18736 2450
rect 18694 1592 18750 1601
rect 18694 1527 18750 1536
rect 19076 480 19104 3431
rect 19352 1057 19380 4014
rect 20088 3942 20116 4558
rect 20180 4214 20208 4780
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20364 4010 20392 11863
rect 21454 10160 21510 10169
rect 21454 10095 21510 10104
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20456 5574 20484 6666
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20640 5522 20668 6122
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5710 20760 6054
rect 20720 5704 20772 5710
rect 20718 5672 20720 5681
rect 20772 5672 20774 5681
rect 20718 5607 20774 5616
rect 20456 4865 20484 5510
rect 20640 5494 20760 5522
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20442 4856 20498 4865
rect 20442 4791 20498 4800
rect 20548 4690 20576 5034
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20732 4554 20760 5494
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 21008 4282 21036 4626
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 21180 4072 21232 4078
rect 21178 4040 21180 4049
rect 21232 4040 21234 4049
rect 20352 4004 20404 4010
rect 21178 3975 21234 3984
rect 20352 3946 20404 3952
rect 20076 3936 20128 3942
rect 20074 3904 20076 3913
rect 20128 3904 20130 3913
rect 19622 3836 19918 3856
rect 20074 3839 20130 3848
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 21468 3738 21496 10095
rect 24030 7848 24086 7857
rect 24030 7783 24086 7792
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22480 5166 22508 5714
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23662 5672 23718 5681
rect 23492 5166 23520 5646
rect 23662 5607 23718 5616
rect 22468 5160 22520 5166
rect 22466 5128 22468 5137
rect 23480 5160 23532 5166
rect 22520 5128 22522 5137
rect 23480 5102 23532 5108
rect 22466 5063 22522 5072
rect 22098 4856 22154 4865
rect 22098 4791 22100 4800
rect 22152 4791 22154 4800
rect 22560 4820 22612 4826
rect 22100 4762 22152 4768
rect 22560 4762 22612 4768
rect 22190 4720 22246 4729
rect 22100 4684 22152 4690
rect 22190 4655 22246 4664
rect 22100 4626 22152 4632
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21456 3732 21508 3738
rect 21376 3692 21456 3720
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3194 19472 3334
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20088 2990 20116 3130
rect 20180 3058 20208 3470
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20076 2984 20128 2990
rect 19522 2952 19578 2961
rect 20076 2926 20128 2932
rect 20456 2922 20484 3334
rect 20628 3120 20680 3126
rect 20680 3080 20760 3108
rect 20628 3062 20680 3068
rect 19522 2887 19578 2896
rect 20444 2916 20496 2922
rect 19536 1170 19564 2887
rect 20444 2858 20496 2864
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 20258 2816 20314 2825
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19904 2417 19932 2450
rect 19890 2408 19946 2417
rect 19890 2343 19946 2352
rect 19996 2310 20024 2790
rect 20258 2751 20314 2760
rect 19984 2304 20036 2310
rect 19982 2272 19984 2281
rect 20036 2272 20038 2281
rect 19982 2207 20038 2216
rect 19996 2181 20024 2207
rect 19536 1142 19656 1170
rect 19338 1048 19394 1057
rect 19338 983 19394 992
rect 19628 480 19656 1142
rect 20272 480 20300 2751
rect 20732 2650 20760 3080
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20732 1465 20760 2382
rect 20718 1456 20774 1465
rect 20718 1391 20774 1400
rect 20824 480 20852 3402
rect 20916 3369 20944 3538
rect 21088 3392 21140 3398
rect 20902 3360 20958 3369
rect 21088 3334 21140 3340
rect 20902 3295 20958 3304
rect 20916 3194 20944 3295
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21100 3097 21128 3334
rect 21086 3088 21142 3097
rect 21086 3023 21142 3032
rect 21376 2990 21404 3692
rect 21456 3674 21508 3680
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 2145 21220 2450
rect 21178 2136 21234 2145
rect 21178 2071 21234 2080
rect 21362 1456 21418 1465
rect 21362 1391 21418 1400
rect 21376 480 21404 1391
rect 21652 610 21680 4422
rect 21836 3738 21864 4422
rect 22112 3942 22140 4626
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 22112 3641 22140 3878
rect 22098 3632 22154 3641
rect 22008 3596 22060 3602
rect 22098 3567 22154 3576
rect 22008 3538 22060 3544
rect 22020 3194 22048 3538
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22204 2990 22232 4655
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 4321 22508 4422
rect 22466 4312 22522 4321
rect 22466 4247 22522 4256
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 22204 2650 22232 2790
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22204 2394 22232 2450
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 22020 2366 22232 2394
rect 21836 1170 21864 2314
rect 21836 1142 21956 1170
rect 21640 604 21692 610
rect 21640 546 21692 552
rect 21928 480 21956 1142
rect 22020 921 22048 2366
rect 22296 1329 22324 4014
rect 22376 4004 22428 4010
rect 22376 3946 22428 3952
rect 22388 1986 22416 3946
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3505 22508 3878
rect 22572 3738 22600 4762
rect 23676 3738 23704 5607
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 22466 3496 22522 3505
rect 22466 3431 22522 3440
rect 22572 2854 22600 3674
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23124 3194 23152 3538
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23308 2961 23336 3334
rect 23570 3224 23626 3233
rect 23388 3188 23440 3194
rect 23570 3159 23626 3168
rect 23388 3130 23440 3136
rect 23294 2952 23350 2961
rect 23294 2887 23350 2896
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 23400 2553 23428 3130
rect 23584 2990 23612 3159
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23386 2544 23442 2553
rect 23386 2479 23442 2488
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 22388 1958 22508 1986
rect 22282 1320 22338 1329
rect 22282 1255 22338 1264
rect 22006 912 22062 921
rect 22006 847 22062 856
rect 22480 480 22508 1958
rect 23492 1465 23520 2246
rect 23478 1456 23534 1465
rect 23478 1391 23534 1400
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23124 480 23152 546
rect 23676 480 23704 3062
rect 23848 2848 23900 2854
rect 23846 2816 23848 2825
rect 23900 2816 23902 2825
rect 23846 2751 23902 2760
rect 24044 2514 24072 7783
rect 24136 4729 24164 13223
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 24122 4720 24178 4729
rect 24122 4655 24178 4664
rect 25134 4584 25190 4593
rect 25134 4519 25190 4528
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 25148 2514 25176 4519
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 24124 2372 24176 2378
rect 24176 2332 24256 2360
rect 24124 2314 24176 2320
rect 24228 480 24256 2332
rect 24860 2304 24912 2310
rect 24860 2246 24912 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24872 1737 24900 2246
rect 24858 1728 24914 1737
rect 24858 1663 24914 1672
rect 24688 598 24808 626
rect 18234 439 18290 448
rect 18510 0 18566 480
rect 19062 0 19118 480
rect 19614 0 19670 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
rect 23110 0 23166 480
rect 23662 0 23718 480
rect 24214 0 24270 480
rect 24688 241 24716 598
rect 24780 480 24808 598
rect 25332 480 25360 4966
rect 27618 3904 27674 3913
rect 27618 3839 27674 3848
rect 25962 3088 26018 3097
rect 25962 3023 26018 3032
rect 25976 480 26004 3023
rect 27066 2000 27122 2009
rect 27066 1935 27122 1944
rect 26436 598 26556 626
rect 24674 232 24730 241
rect 24674 167 24730 176
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25962 0 26018 480
rect 26436 105 26464 598
rect 26528 480 26556 598
rect 27080 480 27108 1935
rect 27632 480 27660 3839
rect 26422 96 26478 105
rect 26422 31 26478 40
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3974 27648 4030 27704
rect 294 20304 350 20360
rect 1950 24268 2006 24304
rect 1950 24248 1952 24268
rect 1952 24248 2004 24268
rect 2004 24248 2006 24268
rect 2502 24112 2558 24168
rect 2410 23860 2466 23896
rect 2410 23840 2412 23860
rect 2412 23840 2464 23860
rect 2464 23840 2466 23860
rect 1858 23588 1914 23624
rect 1858 23568 1860 23588
rect 1860 23568 1912 23588
rect 1912 23568 1914 23588
rect 1306 13096 1362 13152
rect 1674 18536 1730 18592
rect 1674 17720 1730 17776
rect 1582 17584 1638 17640
rect 1950 20324 2006 20360
rect 1950 20304 1952 20324
rect 1952 20304 2004 20324
rect 2004 20304 2006 20324
rect 1766 14184 1822 14240
rect 294 6296 350 6352
rect 2042 17040 2098 17096
rect 2686 21392 2742 21448
rect 2410 17040 2466 17096
rect 2410 16904 2466 16960
rect 2318 12960 2374 13016
rect 1858 9016 1914 9072
rect 2134 8472 2190 8528
rect 2962 21800 3018 21856
rect 2778 21256 2834 21312
rect 2686 18944 2742 19000
rect 3514 24676 3570 24712
rect 3514 24656 3516 24676
rect 3516 24656 3568 24676
rect 3568 24656 3570 24676
rect 4066 25880 4122 25936
rect 3974 25336 4030 25392
rect 4066 24792 4122 24848
rect 3238 18672 3294 18728
rect 3146 18128 3202 18184
rect 2594 16496 2650 16552
rect 3330 16108 3386 16144
rect 3330 16088 3332 16108
rect 3332 16088 3384 16108
rect 3384 16088 3386 16108
rect 2594 15272 2650 15328
rect 3514 15408 3570 15464
rect 3238 14320 3294 14376
rect 2410 11212 2466 11248
rect 2410 11192 2412 11212
rect 2412 11192 2464 11212
rect 2464 11192 2466 11212
rect 2502 11092 2504 11112
rect 2504 11092 2556 11112
rect 2556 11092 2558 11112
rect 2502 11056 2558 11092
rect 2134 5752 2190 5808
rect 1858 5072 1914 5128
rect 1582 4972 1584 4992
rect 1584 4972 1636 4992
rect 1636 4972 1638 4992
rect 1582 4936 1638 4972
rect 1674 4528 1730 4584
rect 1490 4256 1546 4312
rect 1398 3848 1454 3904
rect 846 3576 902 3632
rect 1858 4392 1914 4448
rect 3238 12280 3294 12336
rect 2410 4664 2466 4720
rect 2686 9596 2688 9616
rect 2688 9596 2740 9616
rect 2740 9596 2742 9616
rect 2686 9560 2742 9596
rect 3974 23432 4030 23488
rect 3974 22616 4030 22672
rect 4894 26560 4950 26616
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4434 23024 4490 23080
rect 4526 21936 4582 21992
rect 4894 21392 4950 21448
rect 3790 19216 3846 19272
rect 4250 19760 4306 19816
rect 3698 18264 3754 18320
rect 4250 19080 4306 19136
rect 3974 17176 4030 17232
rect 3698 15000 3754 15056
rect 3606 13640 3662 13696
rect 3514 13232 3570 13288
rect 3422 11328 3478 11384
rect 3514 11056 3570 11112
rect 2686 7948 2742 7984
rect 2686 7928 2688 7948
rect 2688 7928 2740 7948
rect 2740 7928 2742 7948
rect 3054 9560 3110 9616
rect 3422 9460 3424 9480
rect 3424 9460 3476 9480
rect 3476 9460 3478 9480
rect 3422 9424 3478 9460
rect 3698 13096 3754 13152
rect 3606 8336 3662 8392
rect 3146 6840 3202 6896
rect 2962 3712 3018 3768
rect 2134 3052 2190 3088
rect 2134 3032 2136 3052
rect 2136 3032 2188 3052
rect 2188 3032 2190 3052
rect 1950 2216 2006 2272
rect 2410 1672 2466 1728
rect 2870 584 2926 640
rect 3514 8200 3570 8256
rect 4342 17720 4398 17776
rect 4066 16632 4122 16688
rect 4066 14864 4122 14920
rect 4066 14184 4122 14240
rect 4158 12960 4214 13016
rect 4342 12416 4398 12472
rect 4710 18964 4766 19000
rect 4710 18944 4712 18964
rect 4712 18944 4764 18964
rect 4764 18944 4766 18964
rect 4986 18944 5042 19000
rect 5262 24520 5318 24576
rect 5170 23840 5226 23896
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6274 23860 6330 23896
rect 6274 23840 6276 23860
rect 6276 23840 6328 23860
rect 6328 23840 6330 23860
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 22480 5594 22536
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6182 21564 6184 21584
rect 6184 21564 6236 21584
rect 6236 21564 6238 21584
rect 6182 21528 6238 21564
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5262 19760 5318 19816
rect 4618 18128 4674 18184
rect 4526 14592 4582 14648
rect 5078 18536 5134 18592
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5354 19488 5410 19544
rect 5446 18808 5502 18864
rect 5354 18400 5410 18456
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5446 17176 5502 17232
rect 5354 17040 5410 17096
rect 5078 14456 5134 14512
rect 6090 16940 6092 16960
rect 6092 16940 6144 16960
rect 6144 16940 6146 16960
rect 6090 16904 6146 16940
rect 5630 16668 5632 16688
rect 5632 16668 5684 16688
rect 5684 16668 5686 16688
rect 5630 16632 5686 16668
rect 5998 16496 6054 16552
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5354 15272 5410 15328
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4986 12688 5042 12744
rect 4618 12552 4674 12608
rect 3882 9968 3938 10024
rect 3974 7928 4030 7984
rect 3882 7792 3938 7848
rect 3790 7112 3846 7168
rect 3698 6976 3754 7032
rect 3606 5480 3662 5536
rect 3882 6024 3938 6080
rect 4342 9696 4398 9752
rect 3514 3168 3570 3224
rect 3330 2932 3332 2952
rect 3332 2932 3384 2952
rect 3384 2932 3386 2952
rect 3330 2896 3386 2932
rect 3054 1400 3110 1456
rect 2962 448 3018 504
rect 3790 4276 3846 4312
rect 3790 4256 3792 4276
rect 3792 4256 3844 4276
rect 3844 4256 3846 4276
rect 3882 4120 3938 4176
rect 3790 3168 3846 3224
rect 3606 1944 3662 2000
rect 3698 1400 3754 1456
rect 4066 4684 4122 4720
rect 4066 4664 4068 4684
rect 4068 4664 4120 4684
rect 4120 4664 4122 4684
rect 4434 9324 4436 9344
rect 4436 9324 4488 9344
rect 4488 9324 4490 9344
rect 4434 9288 4490 9324
rect 4434 8472 4490 8528
rect 4342 6840 4398 6896
rect 4342 5752 4398 5808
rect 4434 4972 4436 4992
rect 4436 4972 4488 4992
rect 4488 4972 4490 4992
rect 4434 4936 4490 4972
rect 4250 4392 4306 4448
rect 4250 3440 4306 3496
rect 4158 1672 4214 1728
rect 5262 13640 5318 13696
rect 5170 11328 5226 11384
rect 5538 15036 5540 15056
rect 5540 15036 5592 15056
rect 5592 15036 5594 15056
rect 5538 15000 5594 15036
rect 5538 14864 5594 14920
rect 5446 14320 5502 14376
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6274 17312 6330 17368
rect 6550 24520 6606 24576
rect 6918 19624 6974 19680
rect 6918 19080 6974 19136
rect 7102 20440 7158 20496
rect 7378 20576 7434 20632
rect 7102 19216 7158 19272
rect 7194 17176 7250 17232
rect 6550 16496 6606 16552
rect 6458 15952 6514 16008
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6274 12416 6330 12472
rect 6182 12316 6184 12336
rect 6184 12316 6236 12336
rect 6236 12316 6238 12336
rect 6182 12280 6238 12316
rect 5446 10784 5502 10840
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6090 10784 6146 10840
rect 5538 10548 5540 10568
rect 5540 10548 5592 10568
rect 5592 10548 5594 10568
rect 5538 10512 5594 10548
rect 5630 10124 5686 10160
rect 5630 10104 5632 10124
rect 5632 10104 5684 10124
rect 5684 10104 5686 10124
rect 5078 9152 5134 9208
rect 5078 8608 5134 8664
rect 4710 2624 4766 2680
rect 4710 1536 4766 1592
rect 4710 856 4766 912
rect 5354 9288 5410 9344
rect 5262 8200 5318 8256
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4894 3032 4950 3088
rect 6458 11056 6514 11112
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5630 6976 5686 7032
rect 6642 15700 6698 15736
rect 6642 15680 6644 15700
rect 6644 15680 6696 15700
rect 6696 15680 6698 15700
rect 6366 9288 6422 9344
rect 6182 6976 6238 7032
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5630 5888 5686 5944
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5722 4528 5778 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5722 3848 5778 3904
rect 5446 3576 5502 3632
rect 6366 5480 6422 5536
rect 6550 6296 6606 6352
rect 6458 5208 6514 5264
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5354 2896 5410 2952
rect 5170 2252 5172 2272
rect 5172 2252 5224 2272
rect 5224 2252 5226 2272
rect 5170 2216 5226 2252
rect 5262 992 5318 1048
rect 6090 3304 6146 3360
rect 7102 10668 7158 10704
rect 7102 10648 7104 10668
rect 7104 10648 7156 10668
rect 7156 10648 7158 10668
rect 7194 8780 7196 8800
rect 7196 8780 7248 8800
rect 7248 8780 7250 8800
rect 7194 8744 7250 8780
rect 7102 8200 7158 8256
rect 7378 17448 7434 17504
rect 7746 23704 7802 23760
rect 7654 19508 7710 19544
rect 7654 19488 7656 19508
rect 7656 19488 7708 19508
rect 7708 19488 7710 19508
rect 7746 18284 7802 18320
rect 7746 18264 7748 18284
rect 7748 18264 7800 18284
rect 7800 18264 7802 18284
rect 7746 17720 7802 17776
rect 7562 16632 7618 16688
rect 7746 15136 7802 15192
rect 7562 14320 7618 14376
rect 7378 13368 7434 13424
rect 7378 11076 7434 11112
rect 7378 11056 7380 11076
rect 7380 11056 7432 11076
rect 7432 11056 7434 11076
rect 7470 10956 7472 10976
rect 7472 10956 7524 10976
rect 7524 10956 7526 10976
rect 7470 10920 7526 10956
rect 7378 8200 7434 8256
rect 7102 5480 7158 5536
rect 7010 3712 7066 3768
rect 5998 2916 6054 2952
rect 5998 2896 6000 2916
rect 6000 2896 6052 2916
rect 6052 2896 6054 2916
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6090 1944 6146 2000
rect 7838 10512 7894 10568
rect 8022 10376 8078 10432
rect 7838 8336 7894 8392
rect 8022 8880 8078 8936
rect 7746 6704 7802 6760
rect 7746 5208 7802 5264
rect 7378 4120 7434 4176
rect 7194 2896 7250 2952
rect 7194 1808 7250 1864
rect 7746 1400 7802 1456
rect 8298 27104 8354 27160
rect 8574 24692 8576 24712
rect 8576 24692 8628 24712
rect 8628 24692 8630 24712
rect 8574 24656 8630 24692
rect 9402 24792 9458 24848
rect 8206 24112 8262 24168
rect 8298 23840 8354 23896
rect 8850 23704 8906 23760
rect 8758 23160 8814 23216
rect 8206 22752 8262 22808
rect 9402 21004 9458 21040
rect 9402 20984 9404 21004
rect 9404 20984 9456 21004
rect 9456 20984 9458 21004
rect 9218 20848 9274 20904
rect 9494 20868 9550 20904
rect 9494 20848 9496 20868
rect 9496 20848 9548 20868
rect 9548 20848 9550 20868
rect 8574 20032 8630 20088
rect 8298 19216 8354 19272
rect 8390 17720 8446 17776
rect 8390 15988 8392 16008
rect 8392 15988 8444 16008
rect 8444 15988 8446 16008
rect 8390 15952 8446 15988
rect 8666 19760 8722 19816
rect 8206 11772 8208 11792
rect 8208 11772 8260 11792
rect 8260 11772 8262 11792
rect 8206 11736 8262 11772
rect 8298 11192 8354 11248
rect 8298 9968 8354 10024
rect 8942 19352 8998 19408
rect 9218 18672 9274 18728
rect 9402 18128 9458 18184
rect 9586 17448 9642 17504
rect 9586 15428 9642 15464
rect 9586 15408 9588 15428
rect 9588 15408 9640 15428
rect 9640 15408 9642 15428
rect 8942 12960 8998 13016
rect 9126 12824 9182 12880
rect 8850 12688 8906 12744
rect 8666 10376 8722 10432
rect 8390 8372 8392 8392
rect 8392 8372 8444 8392
rect 8444 8372 8446 8392
rect 8390 8336 8446 8372
rect 8666 8472 8722 8528
rect 8574 7948 8630 7984
rect 8574 7928 8576 7948
rect 8576 7928 8628 7948
rect 8628 7928 8630 7948
rect 8298 5344 8354 5400
rect 8206 3984 8262 4040
rect 8114 2488 8170 2544
rect 7930 856 7986 912
rect 8850 7792 8906 7848
rect 8758 3984 8814 4040
rect 8390 2216 8446 2272
rect 9310 12552 9366 12608
rect 9402 11348 9458 11384
rect 9402 11328 9404 11348
rect 9404 11328 9456 11348
rect 9456 11328 9458 11348
rect 9586 11056 9642 11112
rect 9862 24692 9864 24712
rect 9864 24692 9916 24712
rect 9916 24692 9918 24712
rect 9862 24656 9918 24692
rect 9862 24384 9918 24440
rect 9862 23976 9918 24032
rect 9862 20168 9918 20224
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10322 23180 10378 23216
rect 10322 23160 10324 23180
rect 10324 23160 10376 23180
rect 10376 23160 10378 23180
rect 11058 22888 11114 22944
rect 10966 22752 11022 22808
rect 11518 24112 11574 24168
rect 11242 23704 11298 23760
rect 11242 22752 11298 22808
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10230 21664 10286 21720
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 11150 20848 11206 20904
rect 11426 21292 11428 21312
rect 11428 21292 11480 21312
rect 11480 21292 11482 21312
rect 11426 21256 11482 21292
rect 11426 20304 11482 20360
rect 10322 19252 10324 19272
rect 10324 19252 10376 19272
rect 10376 19252 10378 19272
rect 10322 19216 10378 19252
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10782 19216 10838 19272
rect 10874 16632 10930 16688
rect 10782 15680 10838 15736
rect 10782 15408 10838 15464
rect 9954 14728 10010 14784
rect 9862 12144 9918 12200
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10874 12688 10930 12744
rect 10506 12008 10562 12064
rect 9402 9560 9458 9616
rect 8942 7656 8998 7712
rect 9126 7384 9182 7440
rect 8942 7268 8998 7304
rect 8942 7248 8944 7268
rect 8944 7248 8996 7268
rect 8996 7248 8998 7268
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10322 11212 10378 11248
rect 10322 11192 10324 11212
rect 10324 11192 10376 11212
rect 10376 11192 10378 11212
rect 9678 10376 9734 10432
rect 9586 8200 9642 8256
rect 9770 7656 9826 7712
rect 9678 6976 9734 7032
rect 9034 1264 9090 1320
rect 9310 6160 9366 6216
rect 9494 5752 9550 5808
rect 9678 5636 9734 5672
rect 9678 5616 9680 5636
rect 9680 5616 9732 5636
rect 9732 5616 9734 5636
rect 9954 7112 10010 7168
rect 9954 6704 10010 6760
rect 9954 4392 10010 4448
rect 9678 3440 9734 3496
rect 9494 3032 9550 3088
rect 9862 3596 9918 3632
rect 9862 3576 9864 3596
rect 9864 3576 9916 3596
rect 9916 3576 9918 3596
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11334 19352 11390 19408
rect 11610 20984 11666 21040
rect 11794 21120 11850 21176
rect 11518 20032 11574 20088
rect 11610 19352 11666 19408
rect 11242 13232 11298 13288
rect 11058 12960 11114 13016
rect 11242 12960 11298 13016
rect 11058 12588 11060 12608
rect 11060 12588 11112 12608
rect 11112 12588 11114 12608
rect 11058 12552 11114 12588
rect 11518 12144 11574 12200
rect 10874 10784 10930 10840
rect 10874 10512 10930 10568
rect 10782 9696 10838 9752
rect 11242 10104 11298 10160
rect 10874 9152 10930 9208
rect 10782 9036 10838 9072
rect 10782 9016 10784 9036
rect 10784 9016 10836 9036
rect 10836 9016 10838 9036
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10782 7384 10838 7440
rect 10690 7112 10746 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10598 5364 10654 5400
rect 10598 5344 10600 5364
rect 10600 5344 10652 5364
rect 10652 5344 10654 5364
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3596 10194 3632
rect 10138 3576 10140 3596
rect 10140 3576 10192 3596
rect 10192 3576 10194 3596
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 8942 40 8998 96
rect 11058 8200 11114 8256
rect 11886 19116 11888 19136
rect 11888 19116 11940 19136
rect 11940 19116 11942 19136
rect 11886 19080 11942 19116
rect 11702 18672 11758 18728
rect 11794 17060 11850 17096
rect 11794 17040 11796 17060
rect 11796 17040 11848 17060
rect 11848 17040 11850 17060
rect 12162 23568 12218 23624
rect 12162 23024 12218 23080
rect 12070 22480 12126 22536
rect 12162 22072 12218 22128
rect 12070 21936 12126 21992
rect 12622 23704 12678 23760
rect 12898 23468 12900 23488
rect 12900 23468 12952 23488
rect 12952 23468 12954 23488
rect 12898 23432 12954 23468
rect 12622 22652 12624 22672
rect 12624 22652 12676 22672
rect 12676 22652 12678 22672
rect 12622 22616 12678 22652
rect 12254 20576 12310 20632
rect 12162 19760 12218 19816
rect 12162 18400 12218 18456
rect 12438 18300 12440 18320
rect 12440 18300 12492 18320
rect 12492 18300 12494 18320
rect 12438 18264 12494 18300
rect 12254 16788 12310 16824
rect 12254 16768 12256 16788
rect 12256 16768 12308 16788
rect 12308 16768 12310 16788
rect 12438 16632 12494 16688
rect 11794 16088 11850 16144
rect 11886 15816 11942 15872
rect 11702 11092 11704 11112
rect 11704 11092 11756 11112
rect 11756 11092 11758 11112
rect 11702 11056 11758 11092
rect 11058 7248 11114 7304
rect 11334 7268 11390 7304
rect 11334 7248 11336 7268
rect 11336 7248 11388 7268
rect 11388 7248 11390 7268
rect 11058 6976 11114 7032
rect 11058 6296 11114 6352
rect 11150 6060 11152 6080
rect 11152 6060 11204 6080
rect 11204 6060 11206 6080
rect 11150 6024 11206 6060
rect 11702 6840 11758 6896
rect 11426 5888 11482 5944
rect 11334 5772 11390 5808
rect 11334 5752 11336 5772
rect 11336 5752 11388 5772
rect 11388 5752 11390 5772
rect 10874 2624 10930 2680
rect 11794 4548 11850 4584
rect 11794 4528 11796 4548
rect 11796 4528 11848 4548
rect 11848 4528 11850 4548
rect 11702 3984 11758 4040
rect 11794 3440 11850 3496
rect 12622 15952 12678 16008
rect 12898 22924 12900 22944
rect 12900 22924 12952 22944
rect 12952 22924 12954 22944
rect 12898 22888 12954 22924
rect 12990 21664 13046 21720
rect 12806 19116 12808 19136
rect 12808 19116 12860 19136
rect 12860 19116 12862 19136
rect 12806 19080 12862 19116
rect 13542 24248 13598 24304
rect 14094 23976 14150 24032
rect 13266 22752 13322 22808
rect 13726 22092 13782 22128
rect 13726 22072 13728 22092
rect 13728 22072 13780 22092
rect 13780 22072 13782 22092
rect 13634 21392 13690 21448
rect 14094 22072 14150 22128
rect 14278 21120 14334 21176
rect 14646 23432 14702 23488
rect 13450 18808 13506 18864
rect 12806 17312 12862 17368
rect 13174 17856 13230 17912
rect 12254 11328 12310 11384
rect 12162 10920 12218 10976
rect 12346 9288 12402 9344
rect 12070 7692 12072 7712
rect 12072 7692 12124 7712
rect 12124 7692 12126 7712
rect 12070 7656 12126 7692
rect 12070 7384 12126 7440
rect 12162 4820 12218 4856
rect 12162 4800 12164 4820
rect 12164 4800 12216 4820
rect 12216 4800 12218 4820
rect 12162 3032 12218 3088
rect 11150 2488 11206 2544
rect 12530 6876 12532 6896
rect 12532 6876 12584 6896
rect 12584 6876 12586 6896
rect 12530 6840 12586 6876
rect 12806 12844 12862 12880
rect 12806 12824 12808 12844
rect 12808 12824 12860 12844
rect 12860 12824 12862 12844
rect 13174 13232 13230 13288
rect 12990 12588 12992 12608
rect 12992 12588 13044 12608
rect 13044 12588 13046 12608
rect 12990 12552 13046 12588
rect 12714 10920 12770 10976
rect 12898 10240 12954 10296
rect 12898 9832 12954 9888
rect 12898 9696 12954 9752
rect 12806 9560 12862 9616
rect 12990 9324 12992 9344
rect 12992 9324 13044 9344
rect 13044 9324 13046 9344
rect 12990 9288 13046 9324
rect 12990 7520 13046 7576
rect 12990 6024 13046 6080
rect 12898 5636 12954 5672
rect 12898 5616 12900 5636
rect 12900 5616 12952 5636
rect 12952 5616 12954 5636
rect 12990 3712 13046 3768
rect 12898 3032 12954 3088
rect 13358 11192 13414 11248
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15198 24792 15254 24848
rect 16118 24792 16174 24848
rect 15198 24112 15254 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15658 24248 15714 24304
rect 15290 23180 15346 23216
rect 15290 23160 15292 23180
rect 15292 23160 15344 23180
rect 15344 23160 15346 23180
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14830 21120 14886 21176
rect 14094 18808 14150 18864
rect 13910 15136 13966 15192
rect 14186 14728 14242 14784
rect 14002 13776 14058 13832
rect 13910 12044 13912 12064
rect 13912 12044 13964 12064
rect 13964 12044 13966 12064
rect 13910 12008 13966 12044
rect 13726 10240 13782 10296
rect 13818 8880 13874 8936
rect 13726 8084 13782 8120
rect 13726 8064 13728 8084
rect 13728 8064 13780 8084
rect 13780 8064 13782 8084
rect 12714 1944 12770 2000
rect 12990 1944 13046 2000
rect 13726 4936 13782 4992
rect 13818 4664 13874 4720
rect 13726 4256 13782 4312
rect 13726 3984 13782 4040
rect 13542 3168 13598 3224
rect 13450 2644 13506 2680
rect 13450 2624 13452 2644
rect 13452 2624 13504 2644
rect 13504 2624 13506 2644
rect 13634 2488 13690 2544
rect 14094 10240 14150 10296
rect 14094 9424 14150 9480
rect 14646 14456 14702 14512
rect 14370 11056 14426 11112
rect 14370 10648 14426 10704
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14830 20032 14886 20088
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15566 19252 15568 19272
rect 15568 19252 15620 19272
rect 15620 19252 15622 19272
rect 15566 19216 15622 19252
rect 15750 19760 15806 19816
rect 15382 16632 15438 16688
rect 15290 15952 15346 16008
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15014 14320 15070 14376
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14646 11736 14702 11792
rect 14462 9968 14518 10024
rect 14370 8472 14426 8528
rect 14002 5072 14058 5128
rect 14002 4392 14058 4448
rect 14738 11056 14794 11112
rect 14646 8780 14648 8800
rect 14648 8780 14700 8800
rect 14700 8780 14702 8800
rect 14646 8744 14702 8780
rect 14462 7248 14518 7304
rect 14738 5752 14794 5808
rect 14554 3304 14610 3360
rect 14094 2624 14150 2680
rect 15566 12844 15622 12880
rect 15566 12824 15568 12844
rect 15568 12824 15620 12844
rect 15620 12824 15622 12844
rect 15474 12552 15530 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15198 11620 15254 11656
rect 15198 11600 15200 11620
rect 15200 11600 15252 11620
rect 15252 11600 15254 11620
rect 15290 11192 15346 11248
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15014 10532 15070 10568
rect 15014 10512 15016 10532
rect 15016 10512 15068 10532
rect 15068 10512 15070 10532
rect 15198 10548 15200 10568
rect 15200 10548 15252 10568
rect 15252 10548 15254 10568
rect 15198 10512 15254 10548
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15198 8064 15254 8120
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15566 7792 15622 7848
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14646 2216 14702 2272
rect 15474 3304 15530 3360
rect 15474 3032 15530 3088
rect 15382 2352 15438 2408
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15934 17312 15990 17368
rect 16210 24112 16266 24168
rect 17406 24792 17462 24848
rect 17038 24112 17094 24168
rect 16486 23160 16542 23216
rect 16302 19080 16358 19136
rect 16762 21392 16818 21448
rect 16670 20440 16726 20496
rect 16302 17584 16358 17640
rect 15934 15816 15990 15872
rect 15750 15680 15806 15736
rect 15842 14340 15898 14376
rect 15842 14320 15844 14340
rect 15844 14320 15896 14340
rect 15896 14320 15898 14340
rect 15842 11872 15898 11928
rect 15842 11736 15898 11792
rect 16302 16496 16358 16552
rect 18786 24656 18842 24712
rect 16670 16788 16726 16824
rect 16670 16768 16672 16788
rect 16672 16768 16724 16788
rect 16724 16768 16726 16788
rect 16210 10920 16266 10976
rect 16118 10668 16174 10704
rect 16118 10648 16120 10668
rect 16120 10648 16172 10668
rect 16172 10648 16174 10668
rect 15934 9968 15990 10024
rect 15934 9288 15990 9344
rect 15842 8880 15898 8936
rect 16026 8508 16028 8528
rect 16028 8508 16080 8528
rect 16080 8508 16082 8528
rect 16026 8472 16082 8508
rect 15842 7828 15844 7848
rect 15844 7828 15896 7848
rect 15896 7828 15898 7848
rect 15842 7792 15898 7828
rect 16670 11056 16726 11112
rect 17774 21256 17830 21312
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19982 24792 20038 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20258 24656 20314 24712
rect 18050 19896 18106 19952
rect 18602 18128 18658 18184
rect 17682 14728 17738 14784
rect 17406 13368 17462 13424
rect 17590 13404 17592 13424
rect 17592 13404 17644 13424
rect 17644 13404 17646 13424
rect 17590 13368 17646 13404
rect 17498 12180 17500 12200
rect 17500 12180 17552 12200
rect 17552 12180 17554 12200
rect 17498 12144 17554 12180
rect 18326 10376 18382 10432
rect 17498 8372 17500 8392
rect 17500 8372 17552 8392
rect 17552 8372 17554 8392
rect 17498 8336 17554 8372
rect 17590 8200 17646 8256
rect 16118 5888 16174 5944
rect 16026 2488 16082 2544
rect 15842 2216 15898 2272
rect 15842 720 15898 776
rect 16302 5888 16358 5944
rect 17774 7284 17776 7304
rect 17776 7284 17828 7304
rect 17828 7284 17830 7304
rect 17774 7248 17830 7284
rect 18234 7384 18290 7440
rect 18050 7148 18052 7168
rect 18052 7148 18104 7168
rect 18104 7148 18106 7168
rect 18050 7112 18106 7148
rect 17958 6976 18014 7032
rect 17866 6840 17922 6896
rect 16394 4972 16396 4992
rect 16396 4972 16448 4992
rect 16448 4972 16450 4992
rect 16394 4936 16450 4972
rect 17682 4800 17738 4856
rect 18050 6160 18106 6216
rect 17314 4664 17370 4720
rect 18234 4664 18290 4720
rect 17774 4528 17830 4584
rect 16854 4256 16910 4312
rect 16762 3712 16818 3768
rect 16578 2760 16634 2816
rect 16302 2508 16358 2544
rect 16302 2488 16304 2508
rect 16304 2488 16356 2508
rect 16356 2488 16358 2508
rect 17498 4120 17554 4176
rect 17130 3984 17186 4040
rect 17958 3732 18014 3768
rect 17958 3712 17960 3732
rect 17960 3712 18012 3732
rect 18012 3712 18014 3732
rect 17590 3168 17646 3224
rect 17682 2760 17738 2816
rect 17038 2624 17094 2680
rect 17958 2644 18014 2680
rect 17958 2624 17960 2644
rect 17960 2624 18012 2644
rect 18012 2624 18014 2644
rect 17222 1944 17278 2000
rect 18234 3984 18290 4040
rect 17406 1808 17462 1864
rect 18050 1808 18106 1864
rect 17958 1672 18014 1728
rect 18418 9696 18474 9752
rect 20442 23860 20498 23896
rect 20442 23840 20444 23860
rect 20444 23840 20496 23860
rect 20496 23840 20498 23860
rect 21362 24792 21418 24848
rect 21546 23976 21602 24032
rect 22190 24404 22246 24440
rect 22190 24384 22192 24404
rect 22192 24384 22244 24404
rect 22244 24384 22246 24404
rect 21914 23840 21970 23896
rect 20902 23724 20958 23760
rect 20902 23704 20904 23724
rect 20904 23704 20956 23724
rect 20956 23704 20958 23724
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 23110 23976 23166 24032
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24384 24270 24440
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27066 24248 27122 24304
rect 25962 24112 26018 24168
rect 20074 18128 20130 18184
rect 19062 17992 19118 18048
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20258 16632 20314 16688
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 22374 23180 22430 23216
rect 22374 23160 22376 23180
rect 22376 23160 22428 23180
rect 22428 23160 22430 23180
rect 22006 19352 22062 19408
rect 23570 23296 23626 23352
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23570 21528 23626 21584
rect 27618 21392 27674 21448
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 22466 17312 22522 17368
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 20902 15564 20958 15600
rect 20902 15544 20904 15564
rect 20904 15544 20956 15564
rect 20956 15544 20958 15564
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19338 14864 19394 14920
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24674 13912 24730 13968
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24398 13404 24400 13424
rect 24400 13404 24452 13424
rect 24452 13404 24454 13424
rect 24398 13368 24454 13404
rect 24122 13232 24178 13288
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18694 12280 18750 12336
rect 18142 584 18198 640
rect 18326 1128 18382 1184
rect 10046 176 10102 232
rect 18234 448 18290 504
rect 20350 11872 20406 11928
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18786 10512 18842 10568
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19062 9424 19118 9480
rect 18878 7948 18934 7984
rect 18878 7928 18880 7948
rect 18880 7928 18932 7948
rect 18932 7928 18934 7948
rect 18878 5752 18934 5808
rect 18694 4528 18750 4584
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19522 8336 19578 8392
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20258 6840 20314 6896
rect 19246 5072 19302 5128
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19522 5752 19578 5808
rect 20258 5616 20314 5672
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20074 5208 20130 5264
rect 19062 3440 19118 3496
rect 18694 1536 18750 1592
rect 21454 10104 21510 10160
rect 20718 5652 20720 5672
rect 20720 5652 20772 5672
rect 20772 5652 20774 5672
rect 20718 5616 20774 5652
rect 20442 4800 20498 4856
rect 21178 4020 21180 4040
rect 21180 4020 21232 4040
rect 21232 4020 21234 4040
rect 21178 3984 21234 4020
rect 20074 3884 20076 3904
rect 20076 3884 20128 3904
rect 20128 3884 20130 3904
rect 20074 3848 20130 3884
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 24030 7792 24086 7848
rect 23662 5616 23718 5672
rect 22466 5108 22468 5128
rect 22468 5108 22520 5128
rect 22520 5108 22522 5128
rect 22466 5072 22522 5108
rect 22098 4820 22154 4856
rect 22098 4800 22100 4820
rect 22100 4800 22152 4820
rect 22152 4800 22154 4820
rect 22190 4664 22246 4720
rect 19522 2896 19578 2952
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19890 2352 19946 2408
rect 20258 2760 20314 2816
rect 19982 2252 19984 2272
rect 19984 2252 20036 2272
rect 20036 2252 20038 2272
rect 19982 2216 20038 2252
rect 19338 992 19394 1048
rect 20718 1400 20774 1456
rect 20902 3304 20958 3360
rect 21086 3032 21142 3088
rect 21178 2080 21234 2136
rect 21362 1400 21418 1456
rect 22098 3576 22154 3632
rect 22466 4256 22522 4312
rect 22466 3440 22522 3496
rect 23570 3168 23626 3224
rect 23294 2896 23350 2952
rect 23386 2488 23442 2544
rect 22282 1264 22338 1320
rect 22006 856 22062 912
rect 23478 1400 23534 1456
rect 23846 2796 23848 2816
rect 23848 2796 23900 2816
rect 23900 2796 23902 2816
rect 23846 2760 23902 2796
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24122 4664 24178 4720
rect 25134 4528 25190 4584
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24858 1672 24914 1728
rect 27618 3848 27674 3904
rect 25962 3032 26018 3088
rect 27066 1944 27122 2000
rect 24674 176 24730 232
rect 26422 40 26478 96
<< metal3 >>
rect 0 27706 480 27736
rect 3969 27706 4035 27709
rect 0 27704 4035 27706
rect 0 27648 3974 27704
rect 4030 27648 4035 27704
rect 0 27646 4035 27648
rect 0 27616 480 27646
rect 3969 27643 4035 27646
rect 0 27162 480 27192
rect 8293 27162 8359 27165
rect 0 27160 8359 27162
rect 0 27104 8298 27160
rect 8354 27104 8359 27160
rect 0 27102 8359 27104
rect 0 27072 480 27102
rect 8293 27099 8359 27102
rect 0 26618 480 26648
rect 4889 26618 4955 26621
rect 0 26616 4955 26618
rect 0 26560 4894 26616
rect 4950 26560 4955 26616
rect 0 26558 4955 26560
rect 0 26528 480 26558
rect 4889 26555 4955 26558
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3969 25394 4035 25397
rect 0 25392 4035 25394
rect 0 25336 3974 25392
rect 4030 25336 4035 25392
rect 0 25334 4035 25336
rect 0 25304 480 25334
rect 3969 25331 4035 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 4061 24850 4127 24853
rect 0 24848 4127 24850
rect 0 24792 4066 24848
rect 4122 24792 4127 24848
rect 0 24790 4127 24792
rect 0 24760 480 24790
rect 4061 24787 4127 24790
rect 9397 24850 9463 24853
rect 15193 24850 15259 24853
rect 9397 24848 15259 24850
rect 9397 24792 9402 24848
rect 9458 24792 15198 24848
rect 15254 24792 15259 24848
rect 9397 24790 15259 24792
rect 9397 24787 9463 24790
rect 15193 24787 15259 24790
rect 16113 24850 16179 24853
rect 17401 24850 17467 24853
rect 16113 24848 17467 24850
rect 16113 24792 16118 24848
rect 16174 24792 17406 24848
rect 17462 24792 17467 24848
rect 16113 24790 17467 24792
rect 16113 24787 16179 24790
rect 17401 24787 17467 24790
rect 19977 24850 20043 24853
rect 21357 24850 21423 24853
rect 19977 24848 21423 24850
rect 19977 24792 19982 24848
rect 20038 24792 21362 24848
rect 21418 24792 21423 24848
rect 19977 24790 21423 24792
rect 19977 24787 20043 24790
rect 21357 24787 21423 24790
rect 3509 24714 3575 24717
rect 8569 24714 8635 24717
rect 9857 24716 9923 24717
rect 3509 24712 8635 24714
rect 3509 24656 3514 24712
rect 3570 24656 8574 24712
rect 8630 24656 8635 24712
rect 3509 24654 8635 24656
rect 3509 24651 3575 24654
rect 8569 24651 8635 24654
rect 9806 24652 9812 24716
rect 9876 24714 9923 24716
rect 18781 24714 18847 24717
rect 20253 24714 20319 24717
rect 9876 24712 9968 24714
rect 9918 24656 9968 24712
rect 9876 24654 9968 24656
rect 18781 24712 20319 24714
rect 18781 24656 18786 24712
rect 18842 24656 20258 24712
rect 20314 24656 20319 24712
rect 18781 24654 20319 24656
rect 9876 24652 9923 24654
rect 9857 24651 9923 24652
rect 18781 24651 18847 24654
rect 20253 24651 20319 24654
rect 5257 24578 5323 24581
rect 6545 24578 6611 24581
rect 5257 24576 6611 24578
rect 5257 24520 5262 24576
rect 5318 24520 6550 24576
rect 6606 24520 6611 24576
rect 5257 24518 6611 24520
rect 5257 24515 5323 24518
rect 6545 24515 6611 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 9857 24442 9923 24445
rect 1350 24440 9923 24442
rect 1350 24384 9862 24440
rect 9918 24384 9923 24440
rect 1350 24382 9923 24384
rect 0 24170 480 24200
rect 1350 24170 1410 24382
rect 9857 24379 9923 24382
rect 22185 24442 22251 24445
rect 24209 24442 24275 24445
rect 22185 24440 24275 24442
rect 22185 24384 22190 24440
rect 22246 24384 24214 24440
rect 24270 24384 24275 24440
rect 22185 24382 24275 24384
rect 22185 24379 22251 24382
rect 24209 24379 24275 24382
rect 1945 24306 2011 24309
rect 13537 24306 13603 24309
rect 1945 24304 13603 24306
rect 1945 24248 1950 24304
rect 2006 24248 13542 24304
rect 13598 24248 13603 24304
rect 1945 24246 13603 24248
rect 1945 24243 2011 24246
rect 13537 24243 13603 24246
rect 15653 24306 15719 24309
rect 27061 24306 27127 24309
rect 15653 24304 27127 24306
rect 15653 24248 15658 24304
rect 15714 24248 27066 24304
rect 27122 24248 27127 24304
rect 15653 24246 27127 24248
rect 15653 24243 15719 24246
rect 27061 24243 27127 24246
rect 0 24110 1410 24170
rect 2497 24170 2563 24173
rect 2630 24170 2636 24172
rect 2497 24168 2636 24170
rect 2497 24112 2502 24168
rect 2558 24112 2636 24168
rect 2497 24110 2636 24112
rect 0 24080 480 24110
rect 2497 24107 2563 24110
rect 2630 24108 2636 24110
rect 2700 24108 2706 24172
rect 8201 24170 8267 24173
rect 11513 24170 11579 24173
rect 8201 24168 11579 24170
rect 8201 24112 8206 24168
rect 8262 24112 11518 24168
rect 11574 24112 11579 24168
rect 8201 24110 11579 24112
rect 8201 24107 8267 24110
rect 11513 24107 11579 24110
rect 15193 24170 15259 24173
rect 16205 24170 16271 24173
rect 15193 24168 16271 24170
rect 15193 24112 15198 24168
rect 15254 24112 16210 24168
rect 16266 24112 16271 24168
rect 15193 24110 16271 24112
rect 15193 24107 15259 24110
rect 16205 24107 16271 24110
rect 17033 24170 17099 24173
rect 25957 24170 26023 24173
rect 17033 24168 26023 24170
rect 17033 24112 17038 24168
rect 17094 24112 25962 24168
rect 26018 24112 26023 24168
rect 17033 24110 26023 24112
rect 17033 24107 17099 24110
rect 25957 24107 26023 24110
rect 9857 24034 9923 24037
rect 14089 24034 14155 24037
rect 9857 24032 14155 24034
rect 9857 23976 9862 24032
rect 9918 23976 14094 24032
rect 14150 23976 14155 24032
rect 9857 23974 14155 23976
rect 9857 23971 9923 23974
rect 14089 23971 14155 23974
rect 21541 24034 21607 24037
rect 23105 24034 23171 24037
rect 21541 24032 23171 24034
rect 21541 23976 21546 24032
rect 21602 23976 23110 24032
rect 23166 23976 23171 24032
rect 21541 23974 23171 23976
rect 21541 23971 21607 23974
rect 23105 23971 23171 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2405 23898 2471 23901
rect 5165 23898 5231 23901
rect 2405 23896 5231 23898
rect 2405 23840 2410 23896
rect 2466 23840 5170 23896
rect 5226 23840 5231 23896
rect 2405 23838 5231 23840
rect 2405 23835 2471 23838
rect 5165 23835 5231 23838
rect 6269 23898 6335 23901
rect 8293 23898 8359 23901
rect 6269 23896 8359 23898
rect 6269 23840 6274 23896
rect 6330 23840 8298 23896
rect 8354 23840 8359 23896
rect 6269 23838 8359 23840
rect 6269 23835 6335 23838
rect 8293 23835 8359 23838
rect 20437 23898 20503 23901
rect 21909 23898 21975 23901
rect 20437 23896 21975 23898
rect 20437 23840 20442 23896
rect 20498 23840 21914 23896
rect 21970 23840 21975 23896
rect 20437 23838 21975 23840
rect 20437 23835 20503 23838
rect 21909 23835 21975 23838
rect 7741 23762 7807 23765
rect 8845 23762 8911 23765
rect 11237 23762 11303 23765
rect 7741 23760 11303 23762
rect 7741 23704 7746 23760
rect 7802 23704 8850 23760
rect 8906 23704 11242 23760
rect 11298 23704 11303 23760
rect 7741 23702 11303 23704
rect 7741 23699 7807 23702
rect 8845 23699 8911 23702
rect 11237 23699 11303 23702
rect 12617 23762 12683 23765
rect 20897 23762 20963 23765
rect 12617 23760 20963 23762
rect 12617 23704 12622 23760
rect 12678 23704 20902 23760
rect 20958 23704 20963 23760
rect 12617 23702 20963 23704
rect 12617 23699 12683 23702
rect 20897 23699 20963 23702
rect 0 23626 480 23656
rect 1853 23626 1919 23629
rect 12157 23626 12223 23629
rect 0 23566 1410 23626
rect 0 23536 480 23566
rect 1350 23490 1410 23566
rect 1853 23624 12223 23626
rect 1853 23568 1858 23624
rect 1914 23568 12162 23624
rect 12218 23568 12223 23624
rect 1853 23566 12223 23568
rect 1853 23563 1919 23566
rect 12157 23563 12223 23566
rect 3969 23490 4035 23493
rect 1350 23488 4035 23490
rect 1350 23432 3974 23488
rect 4030 23432 4035 23488
rect 1350 23430 4035 23432
rect 3969 23427 4035 23430
rect 12893 23490 12959 23493
rect 14641 23490 14707 23493
rect 12893 23488 14707 23490
rect 12893 23432 12898 23488
rect 12954 23432 14646 23488
rect 14702 23432 14707 23488
rect 12893 23430 14707 23432
rect 12893 23427 12959 23430
rect 14641 23427 14707 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 23565 23354 23631 23357
rect 27520 23354 28000 23384
rect 23565 23352 28000 23354
rect 23565 23296 23570 23352
rect 23626 23296 28000 23352
rect 23565 23294 28000 23296
rect 23565 23291 23631 23294
rect 27520 23264 28000 23294
rect 8753 23218 8819 23221
rect 4294 23216 8819 23218
rect 4294 23160 8758 23216
rect 8814 23160 8819 23216
rect 4294 23158 8819 23160
rect 0 23082 480 23112
rect 4294 23082 4354 23158
rect 8753 23155 8819 23158
rect 10317 23218 10383 23221
rect 15285 23218 15351 23221
rect 10317 23216 15351 23218
rect 10317 23160 10322 23216
rect 10378 23160 15290 23216
rect 15346 23160 15351 23216
rect 10317 23158 15351 23160
rect 10317 23155 10383 23158
rect 15285 23155 15351 23158
rect 16481 23218 16547 23221
rect 22369 23218 22435 23221
rect 16481 23216 22435 23218
rect 16481 23160 16486 23216
rect 16542 23160 22374 23216
rect 22430 23160 22435 23216
rect 16481 23158 22435 23160
rect 16481 23155 16547 23158
rect 22369 23155 22435 23158
rect 0 23022 4354 23082
rect 4429 23082 4495 23085
rect 12157 23082 12223 23085
rect 4429 23080 12223 23082
rect 4429 23024 4434 23080
rect 4490 23024 12162 23080
rect 12218 23024 12223 23080
rect 4429 23022 12223 23024
rect 0 22992 480 23022
rect 4429 23019 4495 23022
rect 12157 23019 12223 23022
rect 11053 22946 11119 22949
rect 12893 22946 12959 22949
rect 11053 22944 12959 22946
rect 11053 22888 11058 22944
rect 11114 22888 12898 22944
rect 12954 22888 12959 22944
rect 11053 22886 12959 22888
rect 11053 22883 11119 22886
rect 12893 22883 12959 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 8201 22810 8267 22813
rect 10961 22810 11027 22813
rect 8201 22808 11027 22810
rect 8201 22752 8206 22808
rect 8262 22752 10966 22808
rect 11022 22752 11027 22808
rect 8201 22750 11027 22752
rect 8201 22747 8267 22750
rect 10961 22747 11027 22750
rect 11237 22810 11303 22813
rect 13261 22810 13327 22813
rect 11237 22808 13327 22810
rect 11237 22752 11242 22808
rect 11298 22752 13266 22808
rect 13322 22752 13327 22808
rect 11237 22750 13327 22752
rect 11237 22747 11303 22750
rect 13261 22747 13327 22750
rect 3969 22674 4035 22677
rect 12617 22674 12683 22677
rect 3969 22672 12683 22674
rect 3969 22616 3974 22672
rect 4030 22616 12622 22672
rect 12678 22616 12683 22672
rect 3969 22614 12683 22616
rect 3969 22611 4035 22614
rect 12617 22611 12683 22614
rect 0 22538 480 22568
rect 5533 22538 5599 22541
rect 12065 22538 12131 22541
rect 0 22478 4952 22538
rect 0 22448 480 22478
rect 4892 22130 4952 22478
rect 5533 22536 12131 22538
rect 5533 22480 5538 22536
rect 5594 22480 12070 22536
rect 12126 22480 12131 22536
rect 5533 22478 12131 22480
rect 5533 22475 5599 22478
rect 12065 22475 12131 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 12157 22130 12223 22133
rect 4892 22128 12223 22130
rect 4892 22072 12162 22128
rect 12218 22072 12223 22128
rect 4892 22070 12223 22072
rect 12157 22067 12223 22070
rect 13721 22130 13787 22133
rect 14089 22130 14155 22133
rect 13721 22128 14155 22130
rect 13721 22072 13726 22128
rect 13782 22072 14094 22128
rect 14150 22072 14155 22128
rect 13721 22070 14155 22072
rect 13721 22067 13787 22070
rect 14089 22067 14155 22070
rect 4521 21994 4587 21997
rect 12065 21994 12131 21997
rect 4521 21992 12131 21994
rect 4521 21936 4526 21992
rect 4582 21936 12070 21992
rect 12126 21936 12131 21992
rect 4521 21934 12131 21936
rect 4521 21931 4587 21934
rect 12065 21931 12131 21934
rect 0 21858 480 21888
rect 2957 21858 3023 21861
rect 0 21856 3023 21858
rect 0 21800 2962 21856
rect 3018 21800 3023 21856
rect 0 21798 3023 21800
rect 0 21768 480 21798
rect 2957 21795 3023 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10225 21722 10291 21725
rect 12985 21722 13051 21725
rect 10225 21720 13051 21722
rect 10225 21664 10230 21720
rect 10286 21664 12990 21720
rect 13046 21664 13051 21720
rect 10225 21662 13051 21664
rect 10225 21659 10291 21662
rect 12985 21659 13051 21662
rect 6177 21586 6243 21589
rect 23565 21586 23631 21589
rect 6177 21584 23631 21586
rect 6177 21528 6182 21584
rect 6238 21528 23570 21584
rect 23626 21528 23631 21584
rect 6177 21526 23631 21528
rect 6177 21523 6243 21526
rect 23565 21523 23631 21526
rect 2681 21452 2747 21453
rect 2630 21388 2636 21452
rect 2700 21450 2747 21452
rect 4889 21450 4955 21453
rect 13629 21450 13695 21453
rect 2700 21448 2792 21450
rect 2742 21392 2792 21448
rect 2700 21390 2792 21392
rect 4889 21448 13695 21450
rect 4889 21392 4894 21448
rect 4950 21392 13634 21448
rect 13690 21392 13695 21448
rect 4889 21390 13695 21392
rect 2700 21388 2747 21390
rect 2681 21387 2747 21388
rect 4889 21387 4955 21390
rect 13629 21387 13695 21390
rect 16757 21450 16823 21453
rect 27613 21450 27679 21453
rect 16757 21448 27679 21450
rect 16757 21392 16762 21448
rect 16818 21392 27618 21448
rect 27674 21392 27679 21448
rect 16757 21390 27679 21392
rect 16757 21387 16823 21390
rect 27613 21387 27679 21390
rect 0 21314 480 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 480 21254
rect 2773 21251 2839 21254
rect 11421 21314 11487 21317
rect 17769 21314 17835 21317
rect 11421 21312 17835 21314
rect 11421 21256 11426 21312
rect 11482 21256 17774 21312
rect 17830 21256 17835 21312
rect 11421 21254 17835 21256
rect 11421 21251 11487 21254
rect 17769 21251 17835 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 11789 21178 11855 21181
rect 14273 21178 14339 21181
rect 14825 21178 14891 21181
rect 11789 21176 14891 21178
rect 11789 21120 11794 21176
rect 11850 21120 14278 21176
rect 14334 21120 14830 21176
rect 14886 21120 14891 21176
rect 11789 21118 14891 21120
rect 11789 21115 11855 21118
rect 14273 21115 14339 21118
rect 14825 21115 14891 21118
rect 9397 21042 9463 21045
rect 11605 21042 11671 21045
rect 9397 21040 11671 21042
rect 9397 20984 9402 21040
rect 9458 20984 11610 21040
rect 11666 20984 11671 21040
rect 9397 20982 11671 20984
rect 9397 20979 9463 20982
rect 11605 20979 11671 20982
rect 9213 20906 9279 20909
rect 1350 20904 9279 20906
rect 1350 20848 9218 20904
rect 9274 20848 9279 20904
rect 1350 20846 9279 20848
rect 0 20770 480 20800
rect 1350 20770 1410 20846
rect 9213 20843 9279 20846
rect 9489 20906 9555 20909
rect 11145 20906 11211 20909
rect 9489 20904 11211 20906
rect 9489 20848 9494 20904
rect 9550 20848 11150 20904
rect 11206 20848 11211 20904
rect 9489 20846 11211 20848
rect 9489 20843 9555 20846
rect 11145 20843 11211 20846
rect 0 20710 1410 20770
rect 0 20680 480 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 7373 20634 7439 20637
rect 12249 20634 12315 20637
rect 7373 20632 12315 20634
rect 7373 20576 7378 20632
rect 7434 20576 12254 20632
rect 12310 20576 12315 20632
rect 7373 20574 12315 20576
rect 7373 20571 7439 20574
rect 12249 20571 12315 20574
rect 7097 20498 7163 20501
rect 16665 20498 16731 20501
rect 7097 20496 16731 20498
rect 7097 20440 7102 20496
rect 7158 20440 16670 20496
rect 16726 20440 16731 20496
rect 7097 20438 16731 20440
rect 7097 20435 7163 20438
rect 16665 20435 16731 20438
rect 289 20362 355 20365
rect 1945 20362 2011 20365
rect 11421 20362 11487 20365
rect 289 20360 11487 20362
rect 289 20304 294 20360
rect 350 20304 1950 20360
rect 2006 20304 11426 20360
rect 11482 20304 11487 20360
rect 289 20302 11487 20304
rect 289 20299 355 20302
rect 1945 20299 2011 20302
rect 11421 20299 11487 20302
rect 9857 20228 9923 20229
rect 9806 20226 9812 20228
rect 9766 20166 9812 20226
rect 9876 20224 9923 20228
rect 9918 20168 9923 20224
rect 9806 20164 9812 20166
rect 9876 20164 9923 20168
rect 9857 20163 9923 20164
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 8569 20090 8635 20093
rect 0 20088 8635 20090
rect 0 20032 8574 20088
rect 8630 20032 8635 20088
rect 0 20030 8635 20032
rect 0 20000 480 20030
rect 8569 20027 8635 20030
rect 11513 20090 11579 20093
rect 14825 20090 14891 20093
rect 11513 20088 14891 20090
rect 11513 20032 11518 20088
rect 11574 20032 14830 20088
rect 14886 20032 14891 20088
rect 11513 20030 14891 20032
rect 11513 20027 11579 20030
rect 14825 20027 14891 20030
rect 18045 19954 18111 19957
rect 5398 19952 18111 19954
rect 5398 19896 18050 19952
rect 18106 19896 18111 19952
rect 5398 19894 18111 19896
rect 4245 19818 4311 19821
rect 5257 19818 5323 19821
rect 5398 19818 5458 19894
rect 12344 19860 12450 19894
rect 18045 19891 18111 19894
rect 4245 19816 5458 19818
rect 4245 19760 4250 19816
rect 4306 19760 5262 19816
rect 5318 19760 5458 19816
rect 4245 19758 5458 19760
rect 8661 19818 8727 19821
rect 12157 19818 12223 19821
rect 15745 19818 15811 19821
rect 8661 19816 12223 19818
rect 8661 19760 8666 19816
rect 8722 19760 12162 19816
rect 12218 19760 12223 19816
rect 8661 19758 12223 19760
rect 4245 19755 4311 19758
rect 5257 19755 5323 19758
rect 8661 19755 8727 19758
rect 12157 19755 12223 19758
rect 14046 19816 15811 19818
rect 14046 19760 15750 19816
rect 15806 19760 15811 19816
rect 14046 19758 15811 19760
rect 6913 19682 6979 19685
rect 14046 19682 14106 19758
rect 15745 19755 15811 19758
rect 6913 19680 14106 19682
rect 6913 19624 6918 19680
rect 6974 19624 14106 19680
rect 6913 19622 14106 19624
rect 6913 19619 6979 19622
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 5349 19546 5415 19549
rect 0 19544 5415 19546
rect 0 19488 5354 19544
rect 5410 19488 5415 19544
rect 0 19486 5415 19488
rect 0 19456 480 19486
rect 5349 19483 5415 19486
rect 7649 19546 7715 19549
rect 7649 19544 11530 19546
rect 7649 19488 7654 19544
rect 7710 19488 11530 19544
rect 7649 19486 11530 19488
rect 7649 19483 7715 19486
rect 8937 19410 9003 19413
rect 11329 19410 11395 19413
rect 8937 19408 11395 19410
rect 8937 19352 8942 19408
rect 8998 19352 11334 19408
rect 11390 19352 11395 19408
rect 8937 19350 11395 19352
rect 11470 19410 11530 19486
rect 11605 19410 11671 19413
rect 22001 19410 22067 19413
rect 11470 19408 22067 19410
rect 11470 19352 11610 19408
rect 11666 19352 22006 19408
rect 22062 19352 22067 19408
rect 11470 19350 22067 19352
rect 8937 19347 9003 19350
rect 11329 19347 11395 19350
rect 11605 19347 11671 19350
rect 22001 19347 22067 19350
rect 3785 19274 3851 19277
rect 7097 19274 7163 19277
rect 8293 19274 8359 19277
rect 10317 19274 10383 19277
rect 3785 19272 8359 19274
rect 3785 19216 3790 19272
rect 3846 19216 7102 19272
rect 7158 19216 8298 19272
rect 8354 19216 8359 19272
rect 3785 19214 8359 19216
rect 3785 19211 3851 19214
rect 7097 19211 7163 19214
rect 8293 19211 8359 19214
rect 9998 19272 10383 19274
rect 9998 19216 10322 19272
rect 10378 19216 10383 19272
rect 9998 19214 10383 19216
rect 4245 19138 4311 19141
rect 6913 19138 6979 19141
rect 4245 19136 6979 19138
rect 4245 19080 4250 19136
rect 4306 19080 6918 19136
rect 6974 19080 6979 19136
rect 4245 19078 6979 19080
rect 4245 19075 4311 19078
rect 6913 19075 6979 19078
rect 0 19002 480 19032
rect 2681 19002 2747 19005
rect 4705 19002 4771 19005
rect 0 18942 1410 19002
rect 0 18912 480 18942
rect 1350 18866 1410 18942
rect 2681 19000 4771 19002
rect 2681 18944 2686 19000
rect 2742 18944 4710 19000
rect 4766 18944 4771 19000
rect 2681 18942 4771 18944
rect 2681 18939 2747 18942
rect 4705 18939 4771 18942
rect 4981 19002 5047 19005
rect 9998 19002 10058 19214
rect 10317 19211 10383 19214
rect 10777 19274 10843 19277
rect 15561 19274 15627 19277
rect 10777 19272 15627 19274
rect 10777 19216 10782 19272
rect 10838 19216 15566 19272
rect 15622 19216 15627 19272
rect 10777 19214 15627 19216
rect 10777 19211 10843 19214
rect 15561 19211 15627 19214
rect 11881 19138 11947 19141
rect 12801 19138 12867 19141
rect 16297 19138 16363 19141
rect 11881 19136 16363 19138
rect 11881 19080 11886 19136
rect 11942 19080 12806 19136
rect 12862 19080 16302 19136
rect 16358 19080 16363 19136
rect 11881 19078 16363 19080
rect 11881 19075 11947 19078
rect 12801 19075 12867 19078
rect 16297 19075 16363 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 4981 19000 10058 19002
rect 4981 18944 4986 19000
rect 5042 18944 10058 19000
rect 4981 18942 10058 18944
rect 4981 18939 5047 18942
rect 5441 18866 5507 18869
rect 1350 18864 5507 18866
rect 1350 18808 5446 18864
rect 5502 18808 5507 18864
rect 1350 18806 5507 18808
rect 5441 18803 5507 18806
rect 13445 18866 13511 18869
rect 14089 18866 14155 18869
rect 13445 18864 14155 18866
rect 13445 18808 13450 18864
rect 13506 18808 14094 18864
rect 14150 18808 14155 18864
rect 13445 18806 14155 18808
rect 13445 18803 13511 18806
rect 14089 18803 14155 18806
rect 3233 18730 3299 18733
rect 9213 18730 9279 18733
rect 11697 18730 11763 18733
rect 3233 18728 11763 18730
rect 3233 18672 3238 18728
rect 3294 18672 9218 18728
rect 9274 18672 11702 18728
rect 11758 18672 11763 18728
rect 3233 18670 11763 18672
rect 3233 18667 3299 18670
rect 9213 18667 9279 18670
rect 11697 18667 11763 18670
rect 1669 18594 1735 18597
rect 5073 18594 5139 18597
rect 1669 18592 5139 18594
rect 1669 18536 1674 18592
rect 1730 18536 5078 18592
rect 5134 18536 5139 18592
rect 1669 18534 5139 18536
rect 1669 18531 1735 18534
rect 5073 18531 5139 18534
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 5349 18458 5415 18461
rect 12157 18458 12223 18461
rect 0 18456 5415 18458
rect 0 18400 5354 18456
rect 5410 18400 5415 18456
rect 0 18398 5415 18400
rect 0 18368 480 18398
rect 5349 18395 5415 18398
rect 5996 18456 12223 18458
rect 5996 18400 12162 18456
rect 12218 18400 12223 18456
rect 5996 18398 12223 18400
rect 3693 18322 3759 18325
rect 5996 18322 6056 18398
rect 12157 18395 12223 18398
rect 3693 18320 6056 18322
rect 3693 18264 3698 18320
rect 3754 18264 6056 18320
rect 3693 18262 6056 18264
rect 7741 18322 7807 18325
rect 12433 18322 12499 18325
rect 7741 18320 12499 18322
rect 7741 18264 7746 18320
rect 7802 18264 12438 18320
rect 12494 18264 12499 18320
rect 7741 18262 12499 18264
rect 3693 18259 3759 18262
rect 7741 18259 7807 18262
rect 12433 18259 12499 18262
rect 3141 18186 3207 18189
rect 4613 18186 4679 18189
rect 9397 18186 9463 18189
rect 3141 18184 9463 18186
rect 3141 18128 3146 18184
rect 3202 18128 4618 18184
rect 4674 18128 9402 18184
rect 9458 18128 9463 18184
rect 3141 18126 9463 18128
rect 3141 18123 3207 18126
rect 4613 18123 4679 18126
rect 9397 18123 9463 18126
rect 18597 18186 18663 18189
rect 20069 18186 20135 18189
rect 18597 18184 20135 18186
rect 18597 18128 18602 18184
rect 18658 18128 20074 18184
rect 20130 18128 20135 18184
rect 18597 18126 20135 18128
rect 18597 18123 18663 18126
rect 20069 18123 20135 18126
rect 19057 18050 19123 18053
rect 15150 18048 19123 18050
rect 15150 17992 19062 18048
rect 19118 17992 19123 18048
rect 15150 17990 19123 17992
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 13169 17914 13235 17917
rect 15150 17914 15210 17990
rect 19057 17987 19123 17990
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 13169 17912 15210 17914
rect 13169 17856 13174 17912
rect 13230 17856 15210 17912
rect 13169 17854 15210 17856
rect 13169 17851 13235 17854
rect 0 17778 480 17808
rect 1669 17778 1735 17781
rect 0 17776 1735 17778
rect 0 17720 1674 17776
rect 1730 17720 1735 17776
rect 0 17718 1735 17720
rect 0 17688 480 17718
rect 1669 17715 1735 17718
rect 4337 17778 4403 17781
rect 7741 17778 7807 17781
rect 8385 17778 8451 17781
rect 4337 17776 8451 17778
rect 4337 17720 4342 17776
rect 4398 17720 7746 17776
rect 7802 17720 8390 17776
rect 8446 17720 8451 17776
rect 4337 17718 8451 17720
rect 4337 17715 4403 17718
rect 7741 17715 7807 17718
rect 8385 17715 8451 17718
rect 1577 17642 1643 17645
rect 16297 17642 16363 17645
rect 1577 17640 16363 17642
rect 1577 17584 1582 17640
rect 1638 17584 16302 17640
rect 16358 17584 16363 17640
rect 1577 17582 16363 17584
rect 1577 17579 1643 17582
rect 16297 17579 16363 17582
rect 7373 17506 7439 17509
rect 9581 17506 9647 17509
rect 7373 17504 9647 17506
rect 7373 17448 7378 17504
rect 7434 17448 9586 17504
rect 9642 17448 9647 17504
rect 7373 17446 9647 17448
rect 7373 17443 7439 17446
rect 9581 17443 9647 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 6269 17370 6335 17373
rect 12801 17370 12867 17373
rect 6269 17368 12867 17370
rect 6269 17312 6274 17368
rect 6330 17312 12806 17368
rect 12862 17312 12867 17368
rect 6269 17310 12867 17312
rect 6269 17307 6335 17310
rect 12801 17307 12867 17310
rect 15929 17370 15995 17373
rect 22461 17370 22527 17373
rect 15929 17368 22527 17370
rect 15929 17312 15934 17368
rect 15990 17312 22466 17368
rect 22522 17312 22527 17368
rect 15929 17310 22527 17312
rect 15929 17307 15995 17310
rect 22461 17307 22527 17310
rect 0 17234 480 17264
rect 3969 17234 4035 17237
rect 0 17232 4035 17234
rect 0 17176 3974 17232
rect 4030 17176 4035 17232
rect 0 17174 4035 17176
rect 0 17144 480 17174
rect 3969 17171 4035 17174
rect 5441 17234 5507 17237
rect 7189 17234 7255 17237
rect 5441 17232 7255 17234
rect 5441 17176 5446 17232
rect 5502 17176 7194 17232
rect 7250 17176 7255 17232
rect 5441 17174 7255 17176
rect 5441 17171 5507 17174
rect 7189 17171 7255 17174
rect 2037 17098 2103 17101
rect 2405 17098 2471 17101
rect 2037 17096 2471 17098
rect 2037 17040 2042 17096
rect 2098 17040 2410 17096
rect 2466 17040 2471 17096
rect 2037 17038 2471 17040
rect 2037 17035 2103 17038
rect 2405 17035 2471 17038
rect 5349 17098 5415 17101
rect 11789 17098 11855 17101
rect 5349 17096 11855 17098
rect 5349 17040 5354 17096
rect 5410 17040 11794 17096
rect 11850 17040 11855 17096
rect 5349 17038 11855 17040
rect 5349 17035 5415 17038
rect 11789 17035 11855 17038
rect 2405 16962 2471 16965
rect 6085 16962 6151 16965
rect 2405 16960 6151 16962
rect 2405 16904 2410 16960
rect 2466 16904 6090 16960
rect 6146 16904 6151 16960
rect 2405 16902 6151 16904
rect 2405 16899 2471 16902
rect 6085 16899 6151 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 12249 16826 12315 16829
rect 16665 16826 16731 16829
rect 12249 16824 16731 16826
rect 12249 16768 12254 16824
rect 12310 16768 16670 16824
rect 16726 16768 16731 16824
rect 12249 16766 16731 16768
rect 12249 16763 12315 16766
rect 16665 16763 16731 16766
rect 0 16690 480 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 480 16630
rect 4061 16627 4127 16630
rect 5625 16690 5691 16693
rect 7557 16690 7623 16693
rect 5625 16688 7623 16690
rect 5625 16632 5630 16688
rect 5686 16632 7562 16688
rect 7618 16632 7623 16688
rect 5625 16630 7623 16632
rect 5625 16627 5691 16630
rect 7557 16627 7623 16630
rect 10869 16690 10935 16693
rect 12433 16690 12499 16693
rect 10869 16688 12499 16690
rect 10869 16632 10874 16688
rect 10930 16632 12438 16688
rect 12494 16632 12499 16688
rect 10869 16630 12499 16632
rect 10869 16627 10935 16630
rect 12433 16627 12499 16630
rect 15377 16690 15443 16693
rect 20253 16690 20319 16693
rect 15377 16688 20319 16690
rect 15377 16632 15382 16688
rect 15438 16632 20258 16688
rect 20314 16632 20319 16688
rect 15377 16630 20319 16632
rect 15377 16627 15443 16630
rect 20253 16627 20319 16630
rect 2589 16554 2655 16557
rect 5993 16554 6059 16557
rect 2589 16552 6059 16554
rect 2589 16496 2594 16552
rect 2650 16496 5998 16552
rect 6054 16496 6059 16552
rect 2589 16494 6059 16496
rect 2589 16491 2655 16494
rect 5993 16491 6059 16494
rect 6545 16554 6611 16557
rect 16297 16554 16363 16557
rect 6545 16552 16363 16554
rect 6545 16496 6550 16552
rect 6606 16496 16302 16552
rect 16358 16496 16363 16552
rect 6545 16494 16363 16496
rect 6545 16491 6611 16494
rect 16297 16491 16363 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 3325 16146 3391 16149
rect 11789 16146 11855 16149
rect 3325 16144 11855 16146
rect 3325 16088 3330 16144
rect 3386 16088 11794 16144
rect 11850 16088 11855 16144
rect 3325 16086 11855 16088
rect 3325 16083 3391 16086
rect 11789 16083 11855 16086
rect 0 16010 480 16040
rect 6453 16010 6519 16013
rect 0 16008 6519 16010
rect 0 15952 6458 16008
rect 6514 15952 6519 16008
rect 0 15950 6519 15952
rect 0 15920 480 15950
rect 6453 15947 6519 15950
rect 8385 16010 8451 16013
rect 12617 16010 12683 16013
rect 15285 16012 15351 16013
rect 15285 16010 15332 16012
rect 8385 16008 12683 16010
rect 8385 15952 8390 16008
rect 8446 15952 12622 16008
rect 12678 15952 12683 16008
rect 8385 15950 12683 15952
rect 15240 16008 15332 16010
rect 15240 15952 15290 16008
rect 15240 15950 15332 15952
rect 8385 15947 8451 15950
rect 12617 15947 12683 15950
rect 15285 15948 15332 15950
rect 15396 15948 15402 16012
rect 15285 15947 15351 15948
rect 11881 15874 11947 15877
rect 15929 15874 15995 15877
rect 11881 15872 15995 15874
rect 11881 15816 11886 15872
rect 11942 15816 15934 15872
rect 15990 15816 15995 15872
rect 11881 15814 15995 15816
rect 11881 15811 11947 15814
rect 15929 15811 15995 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 6637 15738 6703 15741
rect 10777 15738 10843 15741
rect 15745 15738 15811 15741
rect 6637 15736 9552 15738
rect 6637 15680 6642 15736
rect 6698 15704 9552 15736
rect 10777 15736 15811 15738
rect 6698 15680 9644 15704
rect 6637 15678 9644 15680
rect 6637 15675 6703 15678
rect 9492 15644 9644 15678
rect 10777 15680 10782 15736
rect 10838 15680 15750 15736
rect 15806 15680 15811 15736
rect 10777 15678 15811 15680
rect 10777 15675 10843 15678
rect 15745 15675 15811 15678
rect 9584 15602 9644 15644
rect 20897 15602 20963 15605
rect 9584 15600 20963 15602
rect 9584 15544 20902 15600
rect 20958 15544 20963 15600
rect 9584 15542 20963 15544
rect 20897 15539 20963 15542
rect 0 15466 480 15496
rect 3509 15466 3575 15469
rect 0 15464 3575 15466
rect 0 15408 3514 15464
rect 3570 15408 3575 15464
rect 0 15406 3575 15408
rect 0 15376 480 15406
rect 3509 15403 3575 15406
rect 9581 15466 9647 15469
rect 10777 15466 10843 15469
rect 9581 15464 10843 15466
rect 9581 15408 9586 15464
rect 9642 15408 10782 15464
rect 10838 15408 10843 15464
rect 9581 15406 10843 15408
rect 9581 15403 9647 15406
rect 10777 15403 10843 15406
rect 2589 15330 2655 15333
rect 5349 15330 5415 15333
rect 2589 15328 5415 15330
rect 2589 15272 2594 15328
rect 2650 15272 5354 15328
rect 5410 15272 5415 15328
rect 2589 15270 5415 15272
rect 2589 15267 2655 15270
rect 5349 15267 5415 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 7741 15194 7807 15197
rect 13905 15194 13971 15197
rect 7741 15192 13971 15194
rect 7741 15136 7746 15192
rect 7802 15136 13910 15192
rect 13966 15136 13971 15192
rect 7741 15134 13971 15136
rect 7741 15131 7807 15134
rect 13905 15131 13971 15134
rect 3693 15058 3759 15061
rect 5533 15058 5599 15061
rect 3693 15056 5599 15058
rect 3693 15000 3698 15056
rect 3754 15000 5538 15056
rect 5594 15000 5599 15056
rect 3693 14998 5599 15000
rect 3693 14995 3759 14998
rect 5533 14995 5599 14998
rect 0 14922 480 14952
rect 4061 14922 4127 14925
rect 5533 14922 5599 14925
rect 19333 14922 19399 14925
rect 0 14862 3986 14922
rect 0 14832 480 14862
rect 3926 14786 3986 14862
rect 4061 14920 5599 14922
rect 4061 14864 4066 14920
rect 4122 14864 5538 14920
rect 5594 14864 5599 14920
rect 4061 14862 5599 14864
rect 4061 14859 4127 14862
rect 5533 14859 5599 14862
rect 10136 14920 19399 14922
rect 10136 14864 19338 14920
rect 19394 14864 19399 14920
rect 10136 14862 19399 14864
rect 9949 14786 10015 14789
rect 3926 14784 10015 14786
rect 3926 14728 9954 14784
rect 10010 14728 10015 14784
rect 3926 14726 10015 14728
rect 9949 14723 10015 14726
rect 4521 14650 4587 14653
rect 10136 14650 10196 14862
rect 19333 14859 19399 14862
rect 14181 14786 14247 14789
rect 17677 14786 17743 14789
rect 14181 14784 17743 14786
rect 14181 14728 14186 14784
rect 14242 14728 17682 14784
rect 17738 14728 17743 14784
rect 14181 14726 17743 14728
rect 14181 14723 14247 14726
rect 17677 14723 17743 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 4521 14648 10196 14650
rect 4521 14592 4526 14648
rect 4582 14592 10196 14648
rect 4521 14590 10196 14592
rect 4521 14587 4587 14590
rect 5073 14514 5139 14517
rect 14641 14514 14707 14517
rect 5073 14512 14707 14514
rect 5073 14456 5078 14512
rect 5134 14456 14646 14512
rect 14702 14456 14707 14512
rect 5073 14454 14707 14456
rect 5073 14451 5139 14454
rect 14641 14451 14707 14454
rect 0 14378 480 14408
rect 3233 14378 3299 14381
rect 0 14376 3299 14378
rect 0 14320 3238 14376
rect 3294 14320 3299 14376
rect 0 14318 3299 14320
rect 0 14288 480 14318
rect 3233 14315 3299 14318
rect 5441 14378 5507 14381
rect 7557 14378 7623 14381
rect 15009 14378 15075 14381
rect 15837 14378 15903 14381
rect 5441 14376 15903 14378
rect 5441 14320 5446 14376
rect 5502 14320 7562 14376
rect 7618 14320 15014 14376
rect 15070 14320 15842 14376
rect 15898 14320 15903 14376
rect 5441 14318 15903 14320
rect 5441 14315 5507 14318
rect 7557 14315 7623 14318
rect 15009 14315 15075 14318
rect 15837 14315 15903 14318
rect 1761 14242 1827 14245
rect 4061 14242 4127 14245
rect 1761 14240 4127 14242
rect 1761 14184 1766 14240
rect 1822 14184 4066 14240
rect 4122 14184 4127 14240
rect 1761 14182 4127 14184
rect 1761 14179 1827 14182
rect 4061 14179 4127 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 24669 13970 24735 13973
rect 27520 13970 28000 14000
rect 24669 13968 28000 13970
rect 24669 13912 24674 13968
rect 24730 13912 28000 13968
rect 24669 13910 28000 13912
rect 24669 13907 24735 13910
rect 27520 13880 28000 13910
rect 13997 13834 14063 13837
rect 10136 13832 14063 13834
rect 10136 13776 14002 13832
rect 14058 13776 14063 13832
rect 10136 13774 14063 13776
rect 0 13698 480 13728
rect 3601 13698 3667 13701
rect 0 13696 3667 13698
rect 0 13640 3606 13696
rect 3662 13640 3667 13696
rect 0 13638 3667 13640
rect 0 13608 480 13638
rect 3601 13635 3667 13638
rect 5257 13698 5323 13701
rect 10136 13698 10196 13774
rect 13997 13771 14063 13774
rect 5257 13696 10196 13698
rect 5257 13640 5262 13696
rect 5318 13640 10196 13696
rect 5257 13638 10196 13640
rect 5257 13635 5323 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 7373 13426 7439 13429
rect 17401 13426 17467 13429
rect 7373 13424 17467 13426
rect 7373 13368 7378 13424
rect 7434 13368 17406 13424
rect 17462 13368 17467 13424
rect 7373 13366 17467 13368
rect 7373 13363 7439 13366
rect 17401 13363 17467 13366
rect 17585 13426 17651 13429
rect 24393 13426 24459 13429
rect 17585 13424 24459 13426
rect 17585 13368 17590 13424
rect 17646 13368 24398 13424
rect 24454 13368 24459 13424
rect 17585 13366 24459 13368
rect 17585 13363 17651 13366
rect 24393 13363 24459 13366
rect 3509 13290 3575 13293
rect 11237 13290 11303 13293
rect 3509 13288 11303 13290
rect 3509 13232 3514 13288
rect 3570 13232 11242 13288
rect 11298 13232 11303 13288
rect 3509 13230 11303 13232
rect 3509 13227 3575 13230
rect 11237 13227 11303 13230
rect 13169 13290 13235 13293
rect 24117 13290 24183 13293
rect 13169 13288 24183 13290
rect 13169 13232 13174 13288
rect 13230 13232 24122 13288
rect 24178 13232 24183 13288
rect 13169 13230 24183 13232
rect 13169 13227 13235 13230
rect 24117 13227 24183 13230
rect 0 13154 480 13184
rect 1301 13154 1367 13157
rect 3693 13154 3759 13157
rect 0 13152 3759 13154
rect 0 13096 1306 13152
rect 1362 13096 3698 13152
rect 3754 13096 3759 13152
rect 0 13094 3759 13096
rect 0 13064 480 13094
rect 1301 13091 1367 13094
rect 3693 13091 3759 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2313 13018 2379 13021
rect 4153 13018 4219 13021
rect 2313 13016 4219 13018
rect 2313 12960 2318 13016
rect 2374 12960 4158 13016
rect 4214 12960 4219 13016
rect 2313 12958 4219 12960
rect 2313 12955 2379 12958
rect 4153 12955 4219 12958
rect 8937 13018 9003 13021
rect 11053 13018 11119 13021
rect 8937 13016 11119 13018
rect 8937 12960 8942 13016
rect 8998 12960 11058 13016
rect 11114 12960 11119 13016
rect 8937 12958 11119 12960
rect 8937 12955 9003 12958
rect 11053 12955 11119 12958
rect 11237 13018 11303 13021
rect 11237 13016 14842 13018
rect 11237 12960 11242 13016
rect 11298 12960 14842 13016
rect 11237 12958 14842 12960
rect 11237 12955 11303 12958
rect 9121 12882 9187 12885
rect 12801 12882 12867 12885
rect 9121 12880 12867 12882
rect 9121 12824 9126 12880
rect 9182 12824 12806 12880
rect 12862 12824 12867 12880
rect 9121 12822 12867 12824
rect 14782 12882 14842 12958
rect 15561 12882 15627 12885
rect 14782 12880 15627 12882
rect 14782 12824 15566 12880
rect 15622 12824 15627 12880
rect 14782 12822 15627 12824
rect 9121 12819 9187 12822
rect 12801 12819 12867 12822
rect 15561 12819 15627 12822
rect 4981 12746 5047 12749
rect 8845 12746 8911 12749
rect 10869 12746 10935 12749
rect 4981 12744 8911 12746
rect 4981 12688 4986 12744
rect 5042 12688 8850 12744
rect 8906 12688 8911 12744
rect 4981 12686 8911 12688
rect 4981 12683 5047 12686
rect 8845 12683 8911 12686
rect 9446 12686 10748 12746
rect 0 12610 480 12640
rect 4613 12610 4679 12613
rect 9305 12610 9371 12613
rect 0 12608 9371 12610
rect 0 12552 4618 12608
rect 4674 12552 9310 12608
rect 9366 12552 9371 12608
rect 0 12550 9371 12552
rect 0 12520 480 12550
rect 4613 12547 4679 12550
rect 9305 12547 9371 12550
rect 4337 12474 4403 12477
rect 6269 12474 6335 12477
rect 9446 12474 9506 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 4337 12472 9506 12474
rect 4337 12416 4342 12472
rect 4398 12416 6274 12472
rect 6330 12416 9506 12472
rect 4337 12414 9506 12416
rect 10688 12474 10748 12686
rect 10869 12744 14290 12746
rect 10869 12688 10874 12744
rect 10930 12688 14290 12744
rect 10869 12686 14290 12688
rect 10869 12683 10935 12686
rect 11053 12610 11119 12613
rect 12985 12610 13051 12613
rect 11053 12608 13051 12610
rect 11053 12552 11058 12608
rect 11114 12552 12990 12608
rect 13046 12552 13051 12608
rect 11053 12550 13051 12552
rect 14230 12610 14290 12686
rect 15469 12610 15535 12613
rect 14230 12608 15535 12610
rect 14230 12552 15474 12608
rect 15530 12552 15535 12608
rect 14230 12550 15535 12552
rect 11053 12547 11119 12550
rect 12985 12547 13051 12550
rect 15469 12547 15535 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 10688 12414 17418 12474
rect 4337 12411 4403 12414
rect 6269 12411 6335 12414
rect 3233 12338 3299 12341
rect 6177 12338 6243 12341
rect 3233 12336 6243 12338
rect 3233 12280 3238 12336
rect 3294 12280 6182 12336
rect 6238 12280 6243 12336
rect 3233 12278 6243 12280
rect 17358 12338 17418 12414
rect 18689 12338 18755 12341
rect 17358 12336 18755 12338
rect 17358 12280 18694 12336
rect 18750 12280 18755 12336
rect 17358 12278 18755 12280
rect 3233 12275 3299 12278
rect 6177 12275 6243 12278
rect 18689 12275 18755 12278
rect 9857 12202 9923 12205
rect 3006 12200 9923 12202
rect 3006 12144 9862 12200
rect 9918 12144 9923 12200
rect 3006 12142 9923 12144
rect 3006 12066 3066 12142
rect 9857 12139 9923 12142
rect 11513 12202 11579 12205
rect 17493 12202 17559 12205
rect 11513 12200 17559 12202
rect 11513 12144 11518 12200
rect 11574 12144 17498 12200
rect 17554 12144 17559 12200
rect 11513 12142 17559 12144
rect 11513 12139 11579 12142
rect 17493 12139 17559 12142
rect 2684 12006 3066 12066
rect 10501 12066 10567 12069
rect 13905 12066 13971 12069
rect 10501 12064 13971 12066
rect 10501 12008 10506 12064
rect 10562 12008 13910 12064
rect 13966 12008 13971 12064
rect 10501 12006 13971 12008
rect 0 11930 480 11960
rect 2684 11930 2744 12006
rect 10501 12003 10567 12006
rect 13905 12003 13971 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11870 2744 11930
rect 15837 11930 15903 11933
rect 20345 11930 20411 11933
rect 15837 11928 20411 11930
rect 15837 11872 15842 11928
rect 15898 11872 20350 11928
rect 20406 11872 20411 11928
rect 15837 11870 20411 11872
rect 0 11840 480 11870
rect 15837 11867 15903 11870
rect 20345 11867 20411 11870
rect 8201 11794 8267 11797
rect 14641 11794 14707 11797
rect 15837 11794 15903 11797
rect 8201 11792 15903 11794
rect 8201 11736 8206 11792
rect 8262 11736 14646 11792
rect 14702 11736 15842 11792
rect 15898 11736 15903 11792
rect 8201 11734 15903 11736
rect 8201 11731 8267 11734
rect 14641 11731 14707 11734
rect 15837 11731 15903 11734
rect 15193 11658 15259 11661
rect 3236 11656 15259 11658
rect 3236 11600 15198 11656
rect 15254 11600 15259 11656
rect 3236 11598 15259 11600
rect 0 11386 480 11416
rect 3236 11386 3296 11598
rect 15193 11595 15259 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3417 11386 3483 11389
rect 5165 11386 5231 11389
rect 0 11326 3296 11386
rect 3374 11384 5231 11386
rect 3374 11328 3422 11384
rect 3478 11328 5170 11384
rect 5226 11328 5231 11384
rect 3374 11326 5231 11328
rect 0 11296 480 11326
rect 3374 11323 3483 11326
rect 5165 11323 5231 11326
rect 9397 11386 9463 11389
rect 12249 11386 12315 11389
rect 9397 11384 10196 11386
rect 9397 11328 9402 11384
rect 9458 11328 10196 11384
rect 9397 11326 10196 11328
rect 9397 11323 9463 11326
rect 2405 11250 2471 11253
rect 3374 11250 3434 11323
rect 9584 11292 9690 11326
rect 10136 11284 10196 11326
rect 12249 11384 13370 11386
rect 12249 11328 12254 11384
rect 12310 11328 13370 11384
rect 12249 11326 13370 11328
rect 12249 11323 12315 11326
rect 10136 11253 10380 11284
rect 13310 11253 13370 11326
rect 8293 11250 8359 11253
rect 2405 11248 3434 11250
rect 2405 11192 2410 11248
rect 2466 11192 3434 11248
rect 2405 11190 3434 11192
rect 6134 11248 8359 11250
rect 6134 11192 8298 11248
rect 8354 11192 8359 11248
rect 10136 11248 10383 11253
rect 10136 11224 10322 11248
rect 6134 11190 8359 11192
rect 2405 11187 2471 11190
rect 2497 11114 2563 11117
rect 3509 11114 3575 11117
rect 6134 11114 6194 11190
rect 8293 11187 8359 11190
rect 10317 11192 10322 11224
rect 10378 11192 10383 11248
rect 10317 11187 10383 11192
rect 13310 11250 13419 11253
rect 15285 11250 15351 11253
rect 13310 11248 15351 11250
rect 13310 11192 13358 11248
rect 13414 11192 15290 11248
rect 15346 11192 15351 11248
rect 13310 11190 15351 11192
rect 13353 11187 13419 11190
rect 15285 11187 15351 11190
rect 2497 11112 6194 11114
rect 2497 11056 2502 11112
rect 2558 11056 3514 11112
rect 3570 11056 6194 11112
rect 2497 11054 6194 11056
rect 6453 11114 6519 11117
rect 7373 11114 7439 11117
rect 6453 11112 7439 11114
rect 6453 11056 6458 11112
rect 6514 11056 7378 11112
rect 7434 11056 7439 11112
rect 6453 11054 7439 11056
rect 2497 11051 2563 11054
rect 3509 11051 3575 11054
rect 6453 11051 6519 11054
rect 7373 11051 7439 11054
rect 9581 11114 9647 11117
rect 11697 11114 11763 11117
rect 9581 11112 11763 11114
rect 9581 11056 9586 11112
rect 9642 11056 11702 11112
rect 11758 11056 11763 11112
rect 9581 11054 11763 11056
rect 9581 11051 9647 11054
rect 11697 11051 11763 11054
rect 14365 11114 14431 11117
rect 14733 11114 14799 11117
rect 16665 11114 16731 11117
rect 14365 11112 16731 11114
rect 14365 11056 14370 11112
rect 14426 11056 14738 11112
rect 14794 11056 16670 11112
rect 16726 11056 16731 11112
rect 14365 11054 16731 11056
rect 14365 11051 14431 11054
rect 14733 11051 14799 11054
rect 16665 11051 16731 11054
rect 7465 10978 7531 10981
rect 12157 10978 12223 10981
rect 12709 10978 12775 10981
rect 7465 10976 11116 10978
rect 7465 10920 7470 10976
rect 7526 10920 11116 10976
rect 7465 10918 11116 10920
rect 7465 10915 7531 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 5441 10842 5507 10845
rect 0 10840 5507 10842
rect 0 10784 5446 10840
rect 5502 10784 5507 10840
rect 0 10782 5507 10784
rect 0 10752 480 10782
rect 5441 10779 5507 10782
rect 6085 10842 6151 10845
rect 10869 10842 10935 10845
rect 6085 10840 10935 10842
rect 6085 10784 6090 10840
rect 6146 10784 10874 10840
rect 10930 10784 10935 10840
rect 6085 10782 10935 10784
rect 11056 10842 11116 10918
rect 12157 10976 12775 10978
rect 12157 10920 12162 10976
rect 12218 10920 12714 10976
rect 12770 10920 12775 10976
rect 12157 10918 12775 10920
rect 12157 10915 12223 10918
rect 12709 10915 12775 10918
rect 15326 10916 15332 10980
rect 15396 10978 15402 10980
rect 16205 10978 16271 10981
rect 15396 10976 16271 10978
rect 15396 10920 16210 10976
rect 16266 10920 16271 10976
rect 15396 10918 16271 10920
rect 15396 10916 15402 10918
rect 16205 10915 16271 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 11056 10782 14842 10842
rect 6085 10779 6151 10782
rect 10869 10779 10935 10782
rect 7097 10706 7163 10709
rect 14365 10706 14431 10709
rect 7097 10704 14431 10706
rect 7097 10648 7102 10704
rect 7158 10648 14370 10704
rect 14426 10648 14431 10704
rect 7097 10646 14431 10648
rect 14782 10706 14842 10782
rect 16113 10706 16179 10709
rect 14782 10704 16179 10706
rect 14782 10648 16118 10704
rect 16174 10648 16179 10704
rect 14782 10646 16179 10648
rect 7097 10643 7163 10646
rect 14365 10643 14431 10646
rect 16113 10643 16179 10646
rect 5533 10570 5599 10573
rect 7833 10570 7899 10573
rect 10869 10570 10935 10573
rect 15009 10570 15075 10573
rect 5533 10568 10748 10570
rect 5533 10512 5538 10568
rect 5594 10512 7838 10568
rect 7894 10512 10748 10568
rect 5533 10510 10748 10512
rect 5533 10507 5599 10510
rect 7833 10507 7899 10510
rect 8017 10434 8083 10437
rect 8661 10434 8727 10437
rect 9673 10434 9739 10437
rect 8017 10432 9739 10434
rect 8017 10376 8022 10432
rect 8078 10376 8666 10432
rect 8722 10376 9678 10432
rect 9734 10376 9739 10432
rect 8017 10374 9739 10376
rect 10688 10434 10748 10510
rect 10869 10568 15075 10570
rect 10869 10512 10874 10568
rect 10930 10512 15014 10568
rect 15070 10512 15075 10568
rect 10869 10510 15075 10512
rect 10869 10507 10935 10510
rect 15009 10507 15075 10510
rect 15193 10570 15259 10573
rect 18781 10570 18847 10573
rect 15193 10568 18847 10570
rect 15193 10512 15198 10568
rect 15254 10512 18786 10568
rect 18842 10512 18847 10568
rect 15193 10510 18847 10512
rect 15193 10507 15259 10510
rect 18781 10507 18847 10510
rect 18321 10434 18387 10437
rect 10688 10432 18387 10434
rect 10688 10376 18326 10432
rect 18382 10376 18387 10432
rect 10688 10374 18387 10376
rect 8017 10371 8083 10374
rect 8661 10371 8727 10374
rect 9673 10371 9739 10374
rect 18321 10371 18387 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 12893 10298 12959 10301
rect 13721 10298 13787 10301
rect 12893 10296 13787 10298
rect 12893 10240 12898 10296
rect 12954 10240 13726 10296
rect 13782 10240 13787 10296
rect 12893 10238 13787 10240
rect 12893 10235 12959 10238
rect 13721 10235 13787 10238
rect 14089 10298 14155 10301
rect 14089 10296 19442 10298
rect 14089 10240 14094 10296
rect 14150 10240 19442 10296
rect 14089 10238 19442 10240
rect 14089 10235 14155 10238
rect 0 10162 480 10192
rect 5625 10162 5691 10165
rect 11237 10162 11303 10165
rect 0 10160 5691 10162
rect 0 10104 5630 10160
rect 5686 10104 5691 10160
rect 0 10102 5691 10104
rect 0 10072 480 10102
rect 5625 10099 5691 10102
rect 8158 10160 11303 10162
rect 8158 10104 11242 10160
rect 11298 10104 11303 10160
rect 8158 10102 11303 10104
rect 19382 10162 19442 10238
rect 21449 10162 21515 10165
rect 19382 10160 21515 10162
rect 19382 10104 21454 10160
rect 21510 10104 21515 10160
rect 19382 10102 21515 10104
rect 3877 10026 3943 10029
rect 8158 10026 8218 10102
rect 11237 10099 11303 10102
rect 21449 10099 21515 10102
rect 3877 10024 8218 10026
rect 3877 9968 3882 10024
rect 3938 9968 8218 10024
rect 3877 9966 8218 9968
rect 8293 10026 8359 10029
rect 14457 10026 14523 10029
rect 15929 10026 15995 10029
rect 8293 10024 14290 10026
rect 8293 9968 8298 10024
rect 8354 9968 14290 10024
rect 8293 9966 14290 9968
rect 3877 9963 3943 9966
rect 8293 9963 8359 9966
rect 12893 9890 12959 9893
rect 6134 9888 12959 9890
rect 6134 9832 12898 9888
rect 12954 9832 12959 9888
rect 6134 9830 12959 9832
rect 14230 9890 14290 9966
rect 14457 10024 15995 10026
rect 14457 9968 14462 10024
rect 14518 9968 15934 10024
rect 15990 9968 15995 10024
rect 14457 9966 15995 9968
rect 14457 9963 14523 9966
rect 15929 9963 15995 9966
rect 14230 9830 14842 9890
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 4337 9754 4403 9757
rect 4337 9752 5458 9754
rect 4337 9696 4342 9752
rect 4398 9696 5458 9752
rect 4337 9694 5458 9696
rect 4337 9691 4403 9694
rect 0 9618 480 9648
rect 2681 9618 2747 9621
rect 3049 9618 3115 9621
rect 0 9558 2514 9618
rect 0 9528 480 9558
rect 2454 9482 2514 9558
rect 2681 9616 3115 9618
rect 2681 9560 2686 9616
rect 2742 9560 3054 9616
rect 3110 9560 3115 9616
rect 2681 9558 3115 9560
rect 5398 9618 5458 9694
rect 6134 9618 6194 9830
rect 12893 9827 12959 9830
rect 10777 9754 10843 9757
rect 12893 9754 12959 9757
rect 10777 9752 12959 9754
rect 10777 9696 10782 9752
rect 10838 9696 12898 9752
rect 12954 9696 12959 9752
rect 10777 9694 12959 9696
rect 10777 9691 10843 9694
rect 12893 9691 12959 9694
rect 5398 9558 6194 9618
rect 9397 9618 9463 9621
rect 12801 9618 12867 9621
rect 9397 9616 12867 9618
rect 9397 9560 9402 9616
rect 9458 9560 12806 9616
rect 12862 9560 12867 9616
rect 9397 9558 12867 9560
rect 14782 9618 14842 9830
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 18413 9754 18479 9757
rect 15334 9752 18479 9754
rect 15334 9696 18418 9752
rect 18474 9696 18479 9752
rect 15334 9694 18479 9696
rect 15334 9618 15394 9694
rect 18413 9691 18479 9694
rect 14782 9558 15394 9618
rect 2681 9555 2747 9558
rect 3049 9555 3115 9558
rect 9397 9555 9463 9558
rect 12801 9555 12867 9558
rect 3417 9482 3483 9485
rect 2454 9480 3483 9482
rect 2454 9424 3422 9480
rect 3478 9424 3483 9480
rect 2454 9422 3483 9424
rect 3417 9419 3483 9422
rect 14089 9482 14155 9485
rect 19057 9482 19123 9485
rect 14089 9480 19123 9482
rect 14089 9424 14094 9480
rect 14150 9424 19062 9480
rect 19118 9424 19123 9480
rect 14089 9422 19123 9424
rect 14089 9419 14155 9422
rect 19057 9419 19123 9422
rect 4429 9346 4495 9349
rect 5349 9346 5415 9349
rect 6361 9346 6427 9349
rect 4429 9344 6427 9346
rect 4429 9288 4434 9344
rect 4490 9288 5354 9344
rect 5410 9288 6366 9344
rect 6422 9288 6427 9344
rect 4429 9286 6427 9288
rect 4429 9283 4495 9286
rect 5349 9283 5415 9286
rect 6361 9283 6427 9286
rect 12341 9346 12407 9349
rect 12985 9346 13051 9349
rect 15929 9346 15995 9349
rect 12341 9344 15995 9346
rect 12341 9288 12346 9344
rect 12402 9288 12990 9344
rect 13046 9288 15934 9344
rect 15990 9288 15995 9344
rect 12341 9286 15995 9288
rect 12341 9283 12407 9286
rect 12985 9283 13051 9286
rect 15929 9283 15995 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 5073 9210 5139 9213
rect 10869 9212 10935 9213
rect 10869 9210 10916 9212
rect 5073 9208 9644 9210
rect 5073 9152 5078 9208
rect 5134 9176 9644 9208
rect 10824 9208 10916 9210
rect 5134 9152 9690 9176
rect 5073 9150 9690 9152
rect 10824 9152 10874 9208
rect 10824 9150 10916 9152
rect 5073 9147 5139 9150
rect 9584 9116 9690 9150
rect 10869 9148 10916 9150
rect 10980 9148 10986 9212
rect 10869 9147 10935 9148
rect 9630 9108 9690 9116
rect 0 9074 480 9104
rect 1853 9074 1919 9077
rect 0 9072 1919 9074
rect 0 9016 1858 9072
rect 1914 9016 1919 9072
rect 9630 9074 9736 9108
rect 10777 9074 10843 9077
rect 9630 9072 10843 9074
rect 9630 9048 10782 9072
rect 0 9014 1919 9016
rect 9676 9016 10782 9048
rect 10838 9016 10843 9072
rect 9676 9014 10843 9016
rect 0 8984 480 9014
rect 1853 9011 1919 9014
rect 10777 9011 10843 9014
rect 8017 8938 8083 8941
rect 13813 8938 13879 8941
rect 15837 8938 15903 8941
rect 8017 8936 13879 8938
rect 8017 8880 8022 8936
rect 8078 8880 13818 8936
rect 13874 8880 13879 8936
rect 8017 8878 13879 8880
rect 8017 8875 8083 8878
rect 13813 8875 13879 8878
rect 14782 8936 15903 8938
rect 14782 8880 15842 8936
rect 15898 8880 15903 8936
rect 14782 8878 15903 8880
rect 7189 8802 7255 8805
rect 14641 8802 14707 8805
rect 14782 8802 14842 8878
rect 15837 8875 15903 8878
rect 7189 8800 14842 8802
rect 7189 8744 7194 8800
rect 7250 8744 14646 8800
rect 14702 8744 14842 8800
rect 7189 8742 14842 8744
rect 7189 8739 7255 8742
rect 14641 8739 14707 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 5073 8666 5139 8669
rect 1948 8664 5139 8666
rect 1948 8608 5078 8664
rect 5134 8608 5139 8664
rect 1948 8606 5139 8608
rect 0 8530 480 8560
rect 1948 8530 2008 8606
rect 5073 8603 5139 8606
rect 0 8470 2008 8530
rect 2129 8530 2195 8533
rect 4429 8530 4495 8533
rect 2129 8528 4495 8530
rect 2129 8472 2134 8528
rect 2190 8472 4434 8528
rect 4490 8472 4495 8528
rect 2129 8470 4495 8472
rect 0 8440 480 8470
rect 2129 8467 2195 8470
rect 4429 8467 4495 8470
rect 8661 8530 8727 8533
rect 14365 8530 14431 8533
rect 16021 8530 16087 8533
rect 8661 8528 16087 8530
rect 8661 8472 8666 8528
rect 8722 8472 14370 8528
rect 14426 8472 16026 8528
rect 16082 8472 16087 8528
rect 8661 8470 16087 8472
rect 8661 8467 8727 8470
rect 14365 8467 14431 8470
rect 16021 8467 16087 8470
rect 3601 8394 3667 8397
rect 7833 8394 7899 8397
rect 8385 8394 8451 8397
rect 3601 8392 8451 8394
rect 3601 8336 3606 8392
rect 3662 8336 7838 8392
rect 7894 8336 8390 8392
rect 8446 8336 8451 8392
rect 3601 8334 8451 8336
rect 3601 8331 3667 8334
rect 7833 8331 7899 8334
rect 8385 8331 8451 8334
rect 17493 8394 17559 8397
rect 19517 8394 19583 8397
rect 17493 8392 19583 8394
rect 17493 8336 17498 8392
rect 17554 8336 19522 8392
rect 19578 8336 19583 8392
rect 17493 8334 19583 8336
rect 17493 8331 17559 8334
rect 19517 8331 19583 8334
rect 3509 8258 3575 8261
rect 5257 8258 5323 8261
rect 7097 8258 7163 8261
rect 3509 8256 7163 8258
rect 3509 8200 3514 8256
rect 3570 8200 5262 8256
rect 5318 8200 7102 8256
rect 7158 8200 7163 8256
rect 3509 8198 7163 8200
rect 3509 8195 3575 8198
rect 5257 8195 5323 8198
rect 7097 8195 7163 8198
rect 7373 8258 7439 8261
rect 9581 8258 9647 8261
rect 7373 8256 9647 8258
rect 7373 8200 7378 8256
rect 7434 8200 9586 8256
rect 9642 8200 9647 8256
rect 7373 8198 9647 8200
rect 7373 8195 7439 8198
rect 9581 8195 9647 8198
rect 11053 8258 11119 8261
rect 17585 8258 17651 8261
rect 11053 8256 17651 8258
rect 11053 8200 11058 8256
rect 11114 8200 17590 8256
rect 17646 8200 17651 8256
rect 11053 8198 17651 8200
rect 11053 8195 11119 8198
rect 17585 8195 17651 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 13721 8122 13787 8125
rect 15193 8122 15259 8125
rect 13721 8120 15259 8122
rect 13721 8064 13726 8120
rect 13782 8064 15198 8120
rect 15254 8064 15259 8120
rect 13721 8062 15259 8064
rect 13721 8059 13787 8062
rect 15193 8059 15259 8062
rect 2681 7986 2747 7989
rect 3969 7986 4035 7989
rect 2681 7984 4035 7986
rect 2681 7928 2686 7984
rect 2742 7928 3974 7984
rect 4030 7928 4035 7984
rect 2681 7926 4035 7928
rect 2681 7923 2747 7926
rect 3969 7923 4035 7926
rect 8569 7986 8635 7989
rect 18873 7986 18939 7989
rect 8569 7984 18939 7986
rect 8569 7928 8574 7984
rect 8630 7928 18878 7984
rect 18934 7928 18939 7984
rect 8569 7926 18939 7928
rect 8569 7923 8635 7926
rect 18873 7923 18939 7926
rect 0 7850 480 7880
rect 3877 7850 3943 7853
rect 0 7848 3943 7850
rect 0 7792 3882 7848
rect 3938 7792 3943 7848
rect 0 7790 3943 7792
rect 0 7760 480 7790
rect 3877 7787 3943 7790
rect 8845 7850 8911 7853
rect 15561 7850 15627 7853
rect 8845 7848 15627 7850
rect 8845 7792 8850 7848
rect 8906 7792 15566 7848
rect 15622 7792 15627 7848
rect 8845 7790 15627 7792
rect 8845 7787 8911 7790
rect 15561 7787 15627 7790
rect 15837 7850 15903 7853
rect 24025 7850 24091 7853
rect 15837 7848 24091 7850
rect 15837 7792 15842 7848
rect 15898 7792 24030 7848
rect 24086 7792 24091 7848
rect 15837 7790 24091 7792
rect 15837 7787 15903 7790
rect 24025 7787 24091 7790
rect 8937 7714 9003 7717
rect 9765 7714 9831 7717
rect 12065 7714 12131 7717
rect 8937 7712 12131 7714
rect 8937 7656 8942 7712
rect 8998 7656 9770 7712
rect 9826 7656 12070 7712
rect 12126 7656 12131 7712
rect 8937 7654 12131 7656
rect 8937 7651 9003 7654
rect 9765 7651 9831 7654
rect 12065 7651 12131 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 12985 7578 13051 7581
rect 6134 7576 13051 7578
rect 6134 7520 12990 7576
rect 13046 7520 13051 7576
rect 6134 7518 13051 7520
rect 0 7306 480 7336
rect 6134 7306 6194 7518
rect 12985 7515 13051 7518
rect 9121 7442 9187 7445
rect 10777 7442 10843 7445
rect 9121 7440 10843 7442
rect 9121 7384 9126 7440
rect 9182 7384 10782 7440
rect 10838 7384 10843 7440
rect 9121 7382 10843 7384
rect 9121 7379 9187 7382
rect 10777 7379 10843 7382
rect 12065 7442 12131 7445
rect 12065 7440 14658 7442
rect 12065 7384 12070 7440
rect 12126 7384 14658 7440
rect 12065 7382 14658 7384
rect 12065 7379 12131 7382
rect 0 7246 6194 7306
rect 8937 7306 9003 7309
rect 11053 7306 11119 7309
rect 8937 7304 11119 7306
rect 8937 7248 8942 7304
rect 8998 7248 11058 7304
rect 11114 7248 11119 7304
rect 8937 7246 11119 7248
rect 0 7216 480 7246
rect 8937 7243 9003 7246
rect 11053 7243 11119 7246
rect 11329 7306 11395 7309
rect 14457 7306 14523 7309
rect 11329 7304 14523 7306
rect 11329 7248 11334 7304
rect 11390 7248 14462 7304
rect 14518 7248 14523 7304
rect 11329 7246 14523 7248
rect 14598 7306 14658 7382
rect 18086 7380 18092 7444
rect 18156 7442 18162 7444
rect 18229 7442 18295 7445
rect 18156 7440 18295 7442
rect 18156 7384 18234 7440
rect 18290 7384 18295 7440
rect 18156 7382 18295 7384
rect 18156 7380 18162 7382
rect 18229 7379 18295 7382
rect 17769 7306 17835 7309
rect 14598 7304 17835 7306
rect 14598 7248 17774 7304
rect 17830 7248 17835 7304
rect 14598 7246 17835 7248
rect 11329 7243 11395 7246
rect 14457 7243 14523 7246
rect 17769 7243 17835 7246
rect 3785 7170 3851 7173
rect 9949 7170 10015 7173
rect 3785 7168 10015 7170
rect 3785 7112 3790 7168
rect 3846 7112 9954 7168
rect 10010 7112 10015 7168
rect 3785 7110 10015 7112
rect 3785 7107 3851 7110
rect 9949 7107 10015 7110
rect 10685 7170 10751 7173
rect 18045 7170 18111 7173
rect 10685 7168 18111 7170
rect 10685 7112 10690 7168
rect 10746 7112 18050 7168
rect 18106 7112 18111 7168
rect 10685 7110 18111 7112
rect 10685 7107 10751 7110
rect 18045 7107 18111 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 3693 7034 3759 7037
rect 5625 7034 5691 7037
rect 3693 7032 5691 7034
rect 3693 6976 3698 7032
rect 3754 6976 5630 7032
rect 5686 6976 5691 7032
rect 3693 6974 5691 6976
rect 3693 6971 3759 6974
rect 5625 6971 5691 6974
rect 6177 7034 6243 7037
rect 9673 7034 9739 7037
rect 6177 7032 9739 7034
rect 6177 6976 6182 7032
rect 6238 6976 9678 7032
rect 9734 6976 9739 7032
rect 6177 6974 9739 6976
rect 6177 6971 6243 6974
rect 9673 6971 9739 6974
rect 11053 7034 11119 7037
rect 17953 7034 18019 7037
rect 11053 7032 18019 7034
rect 11053 6976 11058 7032
rect 11114 6976 17958 7032
rect 18014 6976 18019 7032
rect 11053 6974 18019 6976
rect 11053 6971 11119 6974
rect 17953 6971 18019 6974
rect 3141 6898 3207 6901
rect 4337 6898 4403 6901
rect 3141 6896 4403 6898
rect 3141 6840 3146 6896
rect 3202 6840 4342 6896
rect 4398 6840 4403 6896
rect 3141 6838 4403 6840
rect 3141 6835 3207 6838
rect 4337 6835 4403 6838
rect 11697 6898 11763 6901
rect 12525 6898 12591 6901
rect 11697 6896 12591 6898
rect 11697 6840 11702 6896
rect 11758 6840 12530 6896
rect 12586 6840 12591 6896
rect 11697 6838 12591 6840
rect 11697 6835 11763 6838
rect 12525 6835 12591 6838
rect 17861 6898 17927 6901
rect 20253 6898 20319 6901
rect 17861 6896 20319 6898
rect 17861 6840 17866 6896
rect 17922 6840 20258 6896
rect 20314 6840 20319 6896
rect 17861 6838 20319 6840
rect 17861 6835 17927 6838
rect 20253 6835 20319 6838
rect 0 6762 480 6792
rect 7741 6762 7807 6765
rect 9949 6762 10015 6765
rect 0 6760 10015 6762
rect 0 6704 7746 6760
rect 7802 6704 9954 6760
rect 10010 6704 10015 6760
rect 0 6702 10015 6704
rect 0 6672 480 6702
rect 7741 6699 7807 6702
rect 9949 6699 10015 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 289 6354 355 6357
rect 6545 6354 6611 6357
rect 11053 6354 11119 6357
rect 289 6352 11119 6354
rect 289 6296 294 6352
rect 350 6296 6550 6352
rect 6606 6296 11058 6352
rect 11114 6296 11119 6352
rect 289 6294 11119 6296
rect 289 6291 355 6294
rect 6545 6291 6611 6294
rect 11053 6291 11119 6294
rect 9305 6218 9371 6221
rect 18045 6218 18111 6221
rect 9305 6216 18111 6218
rect 9305 6160 9310 6216
rect 9366 6160 18050 6216
rect 18106 6160 18111 6216
rect 9305 6158 18111 6160
rect 9305 6155 9371 6158
rect 18045 6155 18111 6158
rect 0 6082 480 6112
rect 3877 6082 3943 6085
rect 0 6080 3943 6082
rect 0 6024 3882 6080
rect 3938 6024 3943 6080
rect 0 6022 3943 6024
rect 0 5992 480 6022
rect 3877 6019 3943 6022
rect 11145 6082 11211 6085
rect 12985 6082 13051 6085
rect 11145 6080 13051 6082
rect 11145 6024 11150 6080
rect 11206 6024 12990 6080
rect 13046 6024 13051 6080
rect 11145 6022 13051 6024
rect 11145 6019 11211 6022
rect 12985 6019 13051 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5625 5946 5691 5949
rect 11421 5946 11487 5949
rect 16113 5946 16179 5949
rect 5625 5944 10058 5946
rect 5625 5888 5630 5944
rect 5686 5888 10058 5944
rect 5625 5886 10058 5888
rect 5625 5883 5691 5886
rect 2129 5810 2195 5813
rect 4337 5810 4403 5813
rect 9489 5812 9555 5813
rect 2129 5808 4403 5810
rect 2129 5752 2134 5808
rect 2190 5752 4342 5808
rect 4398 5752 4403 5808
rect 2129 5750 4403 5752
rect 2129 5747 2195 5750
rect 4337 5747 4403 5750
rect 9438 5748 9444 5812
rect 9508 5810 9555 5812
rect 9998 5810 10058 5886
rect 11421 5944 16179 5946
rect 11421 5888 11426 5944
rect 11482 5888 16118 5944
rect 16174 5888 16179 5944
rect 11421 5886 16179 5888
rect 11421 5883 11487 5886
rect 16113 5883 16179 5886
rect 16297 5946 16363 5949
rect 16297 5944 19442 5946
rect 16297 5888 16302 5944
rect 16358 5888 19442 5944
rect 16297 5886 19442 5888
rect 16297 5883 16363 5886
rect 11329 5810 11395 5813
rect 14733 5810 14799 5813
rect 9508 5808 9600 5810
rect 9550 5752 9600 5808
rect 9508 5750 9600 5752
rect 9998 5808 11395 5810
rect 9998 5752 11334 5808
rect 11390 5752 11395 5808
rect 9998 5750 11395 5752
rect 9508 5748 9555 5750
rect 9489 5747 9555 5748
rect 11329 5747 11395 5750
rect 12758 5808 14799 5810
rect 12758 5752 14738 5808
rect 14794 5752 14799 5808
rect 12758 5750 14799 5752
rect 9673 5674 9739 5677
rect 12758 5674 12818 5750
rect 14733 5747 14799 5750
rect 16614 5748 16620 5812
rect 16684 5810 16690 5812
rect 18873 5810 18939 5813
rect 16684 5808 18939 5810
rect 16684 5752 18878 5808
rect 18934 5752 18939 5808
rect 16684 5750 18939 5752
rect 19382 5810 19442 5886
rect 19517 5810 19583 5813
rect 19382 5808 19583 5810
rect 19382 5752 19522 5808
rect 19578 5752 19583 5808
rect 19382 5750 19583 5752
rect 16684 5748 16690 5750
rect 18873 5747 18939 5750
rect 19517 5747 19583 5750
rect 9673 5672 12818 5674
rect 9673 5616 9678 5672
rect 9734 5616 12818 5672
rect 9673 5614 12818 5616
rect 12893 5674 12959 5677
rect 20253 5674 20319 5677
rect 12893 5672 20319 5674
rect 12893 5616 12898 5672
rect 12954 5616 20258 5672
rect 20314 5616 20319 5672
rect 12893 5614 20319 5616
rect 9673 5611 9739 5614
rect 12893 5611 12959 5614
rect 20253 5611 20319 5614
rect 20713 5674 20779 5677
rect 23657 5674 23723 5677
rect 20713 5672 23723 5674
rect 20713 5616 20718 5672
rect 20774 5616 23662 5672
rect 23718 5616 23723 5672
rect 20713 5614 23723 5616
rect 20713 5611 20779 5614
rect 23657 5611 23723 5614
rect 0 5538 480 5568
rect 3601 5538 3667 5541
rect 0 5536 3667 5538
rect 0 5480 3606 5536
rect 3662 5480 3667 5536
rect 0 5478 3667 5480
rect 0 5448 480 5478
rect 3601 5475 3667 5478
rect 6361 5538 6427 5541
rect 7097 5538 7163 5541
rect 6361 5536 7163 5538
rect 6361 5480 6366 5536
rect 6422 5480 7102 5536
rect 7158 5480 7163 5536
rect 6361 5478 7163 5480
rect 6361 5475 6427 5478
rect 7097 5475 7163 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 8293 5402 8359 5405
rect 10593 5402 10659 5405
rect 8293 5400 10659 5402
rect 8293 5344 8298 5400
rect 8354 5344 10598 5400
rect 10654 5344 10659 5400
rect 8293 5342 10659 5344
rect 8293 5339 8359 5342
rect 10593 5339 10659 5342
rect 6453 5266 6519 5269
rect 7741 5266 7807 5269
rect 20069 5266 20135 5269
rect 6453 5264 20135 5266
rect 6453 5208 6458 5264
rect 6514 5208 7746 5264
rect 7802 5208 20074 5264
rect 20130 5208 20135 5264
rect 6453 5206 20135 5208
rect 6453 5203 6519 5206
rect 7741 5203 7807 5206
rect 20069 5203 20135 5206
rect 1853 5132 1919 5133
rect 1853 5130 1900 5132
rect 1808 5128 1900 5130
rect 1808 5072 1858 5128
rect 1808 5070 1900 5072
rect 1853 5068 1900 5070
rect 1964 5068 1970 5132
rect 10910 5130 10916 5132
rect 9630 5070 10916 5130
rect 1853 5067 1919 5068
rect 0 4994 480 5024
rect 1577 4994 1643 4997
rect 0 4992 1643 4994
rect 0 4936 1582 4992
rect 1638 4936 1643 4992
rect 0 4934 1643 4936
rect 0 4904 480 4934
rect 1577 4931 1643 4934
rect 4429 4994 4495 4997
rect 9630 4996 9690 5070
rect 10910 5068 10916 5070
rect 10980 5068 10986 5132
rect 13997 5130 14063 5133
rect 19241 5130 19307 5133
rect 13997 5128 19307 5130
rect 13997 5072 14002 5128
rect 14058 5072 19246 5128
rect 19302 5072 19307 5128
rect 13997 5070 19307 5072
rect 13997 5067 14063 5070
rect 19241 5067 19307 5070
rect 22318 5068 22324 5132
rect 22388 5130 22394 5132
rect 22461 5130 22527 5133
rect 22388 5128 22527 5130
rect 22388 5072 22466 5128
rect 22522 5072 22527 5128
rect 22388 5070 22527 5072
rect 22388 5068 22394 5070
rect 22461 5067 22527 5070
rect 9622 4994 9628 4996
rect 4429 4992 9628 4994
rect 4429 4936 4434 4992
rect 4490 4936 9628 4992
rect 4429 4934 9628 4936
rect 4429 4931 4495 4934
rect 9622 4932 9628 4934
rect 9692 4932 9698 4996
rect 13721 4994 13787 4997
rect 16389 4994 16455 4997
rect 13721 4992 16455 4994
rect 13721 4936 13726 4992
rect 13782 4936 16394 4992
rect 16450 4936 16455 4992
rect 13721 4934 16455 4936
rect 13721 4931 13787 4934
rect 16389 4931 16455 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 12157 4858 12223 4861
rect 17677 4858 17743 4861
rect 12157 4856 17743 4858
rect 12157 4800 12162 4856
rect 12218 4800 17682 4856
rect 17738 4800 17743 4856
rect 12157 4798 17743 4800
rect 12157 4795 12223 4798
rect 17677 4795 17743 4798
rect 20437 4858 20503 4861
rect 22093 4858 22159 4861
rect 20437 4856 22159 4858
rect 20437 4800 20442 4856
rect 20498 4800 22098 4856
rect 22154 4800 22159 4856
rect 20437 4798 22159 4800
rect 20437 4795 20503 4798
rect 22093 4795 22159 4798
rect 2405 4722 2471 4725
rect 4061 4722 4127 4725
rect 2405 4720 4127 4722
rect 2405 4664 2410 4720
rect 2466 4664 4066 4720
rect 4122 4664 4127 4720
rect 2405 4662 4127 4664
rect 2405 4659 2471 4662
rect 4061 4659 4127 4662
rect 13813 4722 13879 4725
rect 17309 4722 17375 4725
rect 13813 4720 17375 4722
rect 13813 4664 13818 4720
rect 13874 4664 17314 4720
rect 17370 4664 17375 4720
rect 13813 4662 17375 4664
rect 13813 4659 13879 4662
rect 17309 4659 17375 4662
rect 18229 4722 18295 4725
rect 22185 4722 22251 4725
rect 18229 4720 22251 4722
rect 18229 4664 18234 4720
rect 18290 4664 22190 4720
rect 22246 4664 22251 4720
rect 18229 4662 22251 4664
rect 18229 4659 18295 4662
rect 22185 4659 22251 4662
rect 24117 4722 24183 4725
rect 27520 4722 28000 4752
rect 24117 4720 28000 4722
rect 24117 4664 24122 4720
rect 24178 4664 28000 4720
rect 24117 4662 28000 4664
rect 24117 4659 24183 4662
rect 27520 4632 28000 4662
rect 1669 4586 1735 4589
rect 5717 4586 5783 4589
rect 1669 4584 5783 4586
rect 1669 4528 1674 4584
rect 1730 4528 5722 4584
rect 5778 4528 5783 4584
rect 1669 4526 5783 4528
rect 1669 4523 1735 4526
rect 5717 4523 5783 4526
rect 11789 4586 11855 4589
rect 17769 4586 17835 4589
rect 11789 4584 17835 4586
rect 11789 4528 11794 4584
rect 11850 4528 17774 4584
rect 17830 4528 17835 4584
rect 11789 4526 17835 4528
rect 11789 4523 11855 4526
rect 17769 4523 17835 4526
rect 18689 4586 18755 4589
rect 25129 4586 25195 4589
rect 18689 4584 25195 4586
rect 18689 4528 18694 4584
rect 18750 4528 25134 4584
rect 25190 4528 25195 4584
rect 18689 4526 25195 4528
rect 18689 4523 18755 4526
rect 25129 4523 25195 4526
rect 0 4450 480 4480
rect 1853 4450 1919 4453
rect 4245 4450 4311 4453
rect 0 4448 4311 4450
rect 0 4392 1858 4448
rect 1914 4392 4250 4448
rect 4306 4392 4311 4448
rect 0 4390 4311 4392
rect 0 4360 480 4390
rect 1853 4387 1919 4390
rect 4245 4387 4311 4390
rect 9949 4450 10015 4453
rect 13997 4450 14063 4453
rect 9949 4448 14063 4450
rect 9949 4392 9954 4448
rect 10010 4392 14002 4448
rect 14058 4392 14063 4448
rect 9949 4390 14063 4392
rect 9949 4387 10015 4390
rect 13997 4387 14063 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 1485 4314 1551 4317
rect 3785 4314 3851 4317
rect 13721 4314 13787 4317
rect 1485 4312 3851 4314
rect 1485 4256 1490 4312
rect 1546 4256 3790 4312
rect 3846 4256 3851 4312
rect 1485 4254 3851 4256
rect 1485 4251 1551 4254
rect 3785 4251 3851 4254
rect 6134 4312 13787 4314
rect 6134 4256 13726 4312
rect 13782 4256 13787 4312
rect 6134 4254 13787 4256
rect 3877 4178 3943 4181
rect 6134 4178 6194 4254
rect 13721 4251 13787 4254
rect 16849 4314 16915 4317
rect 22461 4314 22527 4317
rect 16849 4312 22527 4314
rect 16849 4256 16854 4312
rect 16910 4256 22466 4312
rect 22522 4256 22527 4312
rect 16849 4254 22527 4256
rect 16849 4251 16915 4254
rect 22461 4251 22527 4254
rect 3877 4176 6194 4178
rect 3877 4120 3882 4176
rect 3938 4120 6194 4176
rect 3877 4118 6194 4120
rect 7373 4178 7439 4181
rect 17493 4178 17559 4181
rect 7373 4176 17559 4178
rect 7373 4120 7378 4176
rect 7434 4120 17498 4176
rect 17554 4120 17559 4176
rect 7373 4118 17559 4120
rect 3877 4115 3943 4118
rect 7373 4115 7439 4118
rect 17493 4115 17559 4118
rect 8201 4044 8267 4045
rect 8150 3980 8156 4044
rect 8220 4042 8267 4044
rect 8753 4042 8819 4045
rect 11697 4042 11763 4045
rect 8220 4040 8312 4042
rect 8262 3984 8312 4040
rect 8220 3982 8312 3984
rect 8753 4040 11763 4042
rect 8753 3984 8758 4040
rect 8814 3984 11702 4040
rect 11758 3984 11763 4040
rect 8753 3982 11763 3984
rect 8220 3980 8267 3982
rect 8201 3979 8267 3980
rect 8753 3979 8819 3982
rect 11697 3979 11763 3982
rect 13721 4042 13787 4045
rect 17125 4042 17191 4045
rect 13721 4040 17191 4042
rect 13721 3984 13726 4040
rect 13782 3984 17130 4040
rect 17186 3984 17191 4040
rect 13721 3982 17191 3984
rect 13721 3979 13787 3982
rect 17125 3979 17191 3982
rect 18229 4042 18295 4045
rect 18229 4040 20362 4042
rect 18229 3984 18234 4040
rect 18290 3984 20362 4040
rect 18229 3982 20362 3984
rect 18229 3979 18295 3982
rect 1393 3906 1459 3909
rect 5717 3906 5783 3909
rect 20069 3908 20135 3909
rect 20069 3906 20116 3908
rect 1393 3904 5783 3906
rect 1393 3848 1398 3904
rect 1454 3848 5722 3904
rect 5778 3848 5783 3904
rect 1393 3846 5783 3848
rect 20024 3904 20116 3906
rect 20024 3848 20074 3904
rect 20024 3846 20116 3848
rect 1393 3843 1459 3846
rect 5717 3843 5783 3846
rect 20069 3844 20116 3846
rect 20180 3844 20186 3908
rect 20302 3906 20362 3982
rect 20478 3980 20484 4044
rect 20548 4042 20554 4044
rect 21173 4042 21239 4045
rect 20548 4040 21239 4042
rect 20548 3984 21178 4040
rect 21234 3984 21239 4040
rect 20548 3982 21239 3984
rect 20548 3980 20554 3982
rect 21173 3979 21239 3982
rect 27613 3906 27679 3909
rect 20302 3904 27679 3906
rect 20302 3848 27618 3904
rect 27674 3848 27679 3904
rect 20302 3846 27679 3848
rect 20069 3843 20135 3844
rect 27613 3843 27679 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2957 3770 3023 3773
rect 7005 3770 7071 3773
rect 12985 3770 13051 3773
rect 16757 3770 16823 3773
rect 0 3768 3023 3770
rect 0 3712 2962 3768
rect 3018 3712 3023 3768
rect 0 3710 3023 3712
rect 0 3680 480 3710
rect 2957 3707 3023 3710
rect 5214 3768 10058 3770
rect 5214 3712 7010 3768
rect 7066 3712 10058 3768
rect 5214 3710 10058 3712
rect 841 3634 907 3637
rect 5214 3634 5274 3710
rect 7005 3707 7071 3710
rect 841 3632 5274 3634
rect 841 3576 846 3632
rect 902 3576 5274 3632
rect 841 3574 5274 3576
rect 5441 3634 5507 3637
rect 9857 3634 9923 3637
rect 5441 3632 9923 3634
rect 5441 3576 5446 3632
rect 5502 3576 9862 3632
rect 9918 3576 9923 3632
rect 5441 3574 9923 3576
rect 841 3571 907 3574
rect 5441 3571 5507 3574
rect 9857 3571 9923 3574
rect 4245 3498 4311 3501
rect 9673 3498 9739 3501
rect 4245 3496 9739 3498
rect 4245 3440 4250 3496
rect 4306 3440 9678 3496
rect 9734 3440 9739 3496
rect 4245 3438 9739 3440
rect 9998 3498 10058 3710
rect 12985 3768 16823 3770
rect 12985 3712 12990 3768
rect 13046 3712 16762 3768
rect 16818 3712 16823 3768
rect 12985 3710 16823 3712
rect 12985 3707 13051 3710
rect 16757 3707 16823 3710
rect 17718 3708 17724 3772
rect 17788 3770 17794 3772
rect 17953 3770 18019 3773
rect 17788 3768 18019 3770
rect 17788 3712 17958 3768
rect 18014 3712 18019 3768
rect 17788 3710 18019 3712
rect 17788 3708 17794 3710
rect 17953 3707 18019 3710
rect 10133 3634 10199 3637
rect 22093 3634 22159 3637
rect 10133 3632 22159 3634
rect 10133 3576 10138 3632
rect 10194 3576 22098 3632
rect 22154 3576 22159 3632
rect 10133 3574 22159 3576
rect 10133 3571 10199 3574
rect 22093 3571 22159 3574
rect 11789 3498 11855 3501
rect 9998 3496 11855 3498
rect 9998 3440 11794 3496
rect 11850 3440 11855 3496
rect 9998 3438 11855 3440
rect 4245 3435 4311 3438
rect 9673 3435 9739 3438
rect 11789 3435 11855 3438
rect 19057 3498 19123 3501
rect 22461 3498 22527 3501
rect 19057 3496 22527 3498
rect 19057 3440 19062 3496
rect 19118 3440 22466 3496
rect 22522 3440 22527 3496
rect 19057 3438 22527 3440
rect 19057 3435 19123 3438
rect 22461 3435 22527 3438
rect 6085 3362 6151 3365
rect 14549 3362 14615 3365
rect 6085 3360 14615 3362
rect 6085 3304 6090 3360
rect 6146 3304 14554 3360
rect 14610 3304 14615 3360
rect 6085 3302 14615 3304
rect 6085 3299 6151 3302
rect 14549 3299 14615 3302
rect 15469 3362 15535 3365
rect 20897 3362 20963 3365
rect 15469 3360 20963 3362
rect 15469 3304 15474 3360
rect 15530 3304 20902 3360
rect 20958 3304 20963 3360
rect 15469 3302 20963 3304
rect 15469 3299 15535 3302
rect 20897 3299 20963 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3509 3226 3575 3229
rect 0 3224 3575 3226
rect 0 3168 3514 3224
rect 3570 3168 3575 3224
rect 0 3166 3575 3168
rect 0 3136 480 3166
rect 3509 3163 3575 3166
rect 3785 3226 3851 3229
rect 13537 3226 13603 3229
rect 3785 3224 5090 3226
rect 3785 3168 3790 3224
rect 3846 3168 5090 3224
rect 3785 3166 5090 3168
rect 3785 3163 3851 3166
rect 2129 3090 2195 3093
rect 4889 3090 4955 3093
rect 2129 3088 4955 3090
rect 2129 3032 2134 3088
rect 2190 3032 4894 3088
rect 4950 3032 4955 3088
rect 2129 3030 4955 3032
rect 5030 3090 5090 3166
rect 6088 3224 13603 3226
rect 6088 3168 13542 3224
rect 13598 3168 13603 3224
rect 6088 3166 13603 3168
rect 6088 3090 6148 3166
rect 13537 3163 13603 3166
rect 17585 3226 17651 3229
rect 23565 3226 23631 3229
rect 17585 3224 23631 3226
rect 17585 3168 17590 3224
rect 17646 3168 23570 3224
rect 23626 3168 23631 3224
rect 17585 3166 23631 3168
rect 17585 3163 17651 3166
rect 23565 3163 23631 3166
rect 5030 3030 6148 3090
rect 9489 3090 9555 3093
rect 12157 3090 12223 3093
rect 9489 3088 12223 3090
rect 9489 3032 9494 3088
rect 9550 3032 12162 3088
rect 12218 3032 12223 3088
rect 9489 3030 12223 3032
rect 2129 3027 2195 3030
rect 4889 3027 4955 3030
rect 9489 3027 9555 3030
rect 12157 3027 12223 3030
rect 12893 3090 12959 3093
rect 15469 3090 15535 3093
rect 12893 3088 15535 3090
rect 12893 3032 12898 3088
rect 12954 3032 15474 3088
rect 15530 3032 15535 3088
rect 12893 3030 15535 3032
rect 12893 3027 12959 3030
rect 15469 3027 15535 3030
rect 21081 3090 21147 3093
rect 25957 3090 26023 3093
rect 21081 3088 26023 3090
rect 21081 3032 21086 3088
rect 21142 3032 25962 3088
rect 26018 3032 26023 3088
rect 21081 3030 26023 3032
rect 21081 3027 21147 3030
rect 25957 3027 26023 3030
rect 3325 2954 3391 2957
rect 5349 2954 5415 2957
rect 3325 2952 5415 2954
rect 3325 2896 3330 2952
rect 3386 2896 5354 2952
rect 5410 2896 5415 2952
rect 3325 2894 5415 2896
rect 3325 2891 3391 2894
rect 5349 2891 5415 2894
rect 5993 2954 6059 2957
rect 7189 2954 7255 2957
rect 19517 2954 19583 2957
rect 23289 2954 23355 2957
rect 5993 2952 10748 2954
rect 5993 2896 5998 2952
rect 6054 2896 7194 2952
rect 7250 2896 10748 2952
rect 5993 2894 10748 2896
rect 5993 2891 6059 2894
rect 7189 2891 7255 2894
rect 10688 2818 10748 2894
rect 19517 2952 23355 2954
rect 19517 2896 19522 2952
rect 19578 2896 23294 2952
rect 23350 2896 23355 2952
rect 19517 2894 23355 2896
rect 19517 2891 19583 2894
rect 23289 2891 23355 2894
rect 16573 2818 16639 2821
rect 17677 2818 17743 2821
rect 10688 2816 17743 2818
rect 10688 2760 16578 2816
rect 16634 2760 17682 2816
rect 17738 2760 17743 2816
rect 10688 2758 17743 2760
rect 16573 2755 16639 2758
rect 17677 2755 17743 2758
rect 20253 2818 20319 2821
rect 23841 2818 23907 2821
rect 20253 2816 23907 2818
rect 20253 2760 20258 2816
rect 20314 2760 23846 2816
rect 23902 2760 23907 2816
rect 20253 2758 23907 2760
rect 20253 2755 20319 2758
rect 23841 2755 23907 2758
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4705 2682 4771 2685
rect 6126 2682 6132 2684
rect 0 2622 3986 2682
rect 0 2592 480 2622
rect 3926 2546 3986 2622
rect 4248 2680 6132 2682
rect 4248 2624 4710 2680
rect 4766 2624 6132 2680
rect 4248 2622 6132 2624
rect 4248 2546 4308 2622
rect 4705 2619 4771 2622
rect 6126 2620 6132 2622
rect 6196 2620 6202 2684
rect 10869 2682 10935 2685
rect 13445 2682 13511 2685
rect 10869 2680 13511 2682
rect 10869 2624 10874 2680
rect 10930 2624 13450 2680
rect 13506 2624 13511 2680
rect 10869 2622 13511 2624
rect 10869 2619 10935 2622
rect 13445 2619 13511 2622
rect 14089 2682 14155 2685
rect 17033 2682 17099 2685
rect 14089 2680 17099 2682
rect 14089 2624 14094 2680
rect 14150 2624 17038 2680
rect 17094 2624 17099 2680
rect 14089 2622 17099 2624
rect 14089 2619 14155 2622
rect 17033 2619 17099 2622
rect 17953 2682 18019 2685
rect 18086 2682 18092 2684
rect 17953 2680 18092 2682
rect 17953 2624 17958 2680
rect 18014 2624 18092 2680
rect 17953 2622 18092 2624
rect 17953 2619 18019 2622
rect 18086 2620 18092 2622
rect 18156 2620 18162 2684
rect 3926 2486 4308 2546
rect 8109 2546 8175 2549
rect 11145 2546 11211 2549
rect 8109 2544 11211 2546
rect 8109 2488 8114 2544
rect 8170 2488 11150 2544
rect 11206 2488 11211 2544
rect 8109 2486 11211 2488
rect 8109 2483 8175 2486
rect 11145 2483 11211 2486
rect 13629 2546 13695 2549
rect 16021 2546 16087 2549
rect 13629 2544 16087 2546
rect 13629 2488 13634 2544
rect 13690 2488 16026 2544
rect 16082 2488 16087 2544
rect 13629 2486 16087 2488
rect 13629 2483 13695 2486
rect 16021 2483 16087 2486
rect 16297 2546 16363 2549
rect 23381 2546 23447 2549
rect 16297 2544 23447 2546
rect 16297 2488 16302 2544
rect 16358 2488 23386 2544
rect 23442 2488 23447 2544
rect 16297 2486 23447 2488
rect 16297 2483 16363 2486
rect 23381 2483 23447 2486
rect 15377 2410 15443 2413
rect 19885 2410 19951 2413
rect 15377 2408 19951 2410
rect 15377 2352 15382 2408
rect 15438 2352 19890 2408
rect 19946 2352 19951 2408
rect 15377 2350 19951 2352
rect 15377 2347 15443 2350
rect 19885 2347 19951 2350
rect 1945 2274 2011 2277
rect 5165 2274 5231 2277
rect 1945 2272 5231 2274
rect 1945 2216 1950 2272
rect 2006 2216 5170 2272
rect 5226 2216 5231 2272
rect 1945 2214 5231 2216
rect 1945 2211 2011 2214
rect 5165 2211 5231 2214
rect 8385 2274 8451 2277
rect 14641 2274 14707 2277
rect 8385 2272 14707 2274
rect 8385 2216 8390 2272
rect 8446 2216 14646 2272
rect 14702 2216 14707 2272
rect 8385 2214 14707 2216
rect 8385 2211 8451 2214
rect 14641 2211 14707 2214
rect 15837 2274 15903 2277
rect 19977 2274 20043 2277
rect 15837 2272 20043 2274
rect 15837 2216 15842 2272
rect 15898 2216 19982 2272
rect 20038 2216 20043 2272
rect 15837 2214 20043 2216
rect 15837 2211 15903 2214
rect 19977 2211 20043 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 21173 2138 21239 2141
rect 16990 2136 21239 2138
rect 16990 2080 21178 2136
rect 21234 2080 21239 2136
rect 16990 2078 21239 2080
rect 0 2002 480 2032
rect 3601 2002 3667 2005
rect 0 2000 3667 2002
rect 0 1944 3606 2000
rect 3662 1944 3667 2000
rect 0 1942 3667 1944
rect 0 1912 480 1942
rect 3601 1939 3667 1942
rect 6085 2002 6151 2005
rect 12709 2002 12775 2005
rect 6085 2000 12775 2002
rect 6085 1944 6090 2000
rect 6146 1944 12714 2000
rect 12770 1944 12775 2000
rect 6085 1942 12775 1944
rect 6085 1939 6151 1942
rect 12709 1939 12775 1942
rect 12985 2002 13051 2005
rect 16990 2002 17050 2078
rect 21173 2075 21239 2078
rect 12985 2000 17050 2002
rect 12985 1944 12990 2000
rect 13046 1944 17050 2000
rect 12985 1942 17050 1944
rect 17217 2002 17283 2005
rect 27061 2002 27127 2005
rect 17217 2000 27127 2002
rect 17217 1944 17222 2000
rect 17278 1944 27066 2000
rect 27122 1944 27127 2000
rect 17217 1942 27127 1944
rect 12985 1939 13051 1942
rect 17217 1939 17283 1942
rect 27061 1939 27127 1942
rect 7189 1866 7255 1869
rect 17401 1866 17467 1869
rect 18045 1866 18111 1869
rect 7189 1864 17467 1866
rect 7189 1808 7194 1864
rect 7250 1808 17406 1864
rect 17462 1808 17467 1864
rect 7189 1806 17467 1808
rect 7189 1803 7255 1806
rect 17401 1803 17467 1806
rect 17542 1864 18111 1866
rect 17542 1808 18050 1864
rect 18106 1808 18111 1864
rect 17542 1806 18111 1808
rect 2405 1730 2471 1733
rect 2630 1730 2636 1732
rect 2405 1728 2636 1730
rect 2405 1672 2410 1728
rect 2466 1672 2636 1728
rect 2405 1670 2636 1672
rect 2405 1667 2471 1670
rect 2630 1668 2636 1670
rect 2700 1668 2706 1732
rect 4153 1730 4219 1733
rect 17542 1730 17602 1806
rect 18045 1803 18111 1806
rect 4153 1728 17602 1730
rect 4153 1672 4158 1728
rect 4214 1672 17602 1728
rect 4153 1670 17602 1672
rect 17953 1730 18019 1733
rect 24853 1730 24919 1733
rect 17953 1728 24919 1730
rect 17953 1672 17958 1728
rect 18014 1672 24858 1728
rect 24914 1672 24919 1728
rect 17953 1670 24919 1672
rect 4153 1667 4219 1670
rect 17953 1667 18019 1670
rect 24853 1667 24919 1670
rect 4705 1594 4771 1597
rect 18689 1594 18755 1597
rect 4705 1592 18755 1594
rect 4705 1536 4710 1592
rect 4766 1536 18694 1592
rect 18750 1536 18755 1592
rect 4705 1534 18755 1536
rect 4705 1531 4771 1534
rect 18689 1531 18755 1534
rect 0 1458 480 1488
rect 3049 1458 3115 1461
rect 0 1456 3115 1458
rect 0 1400 3054 1456
rect 3110 1400 3115 1456
rect 0 1398 3115 1400
rect 0 1368 480 1398
rect 3049 1395 3115 1398
rect 3693 1458 3759 1461
rect 7741 1458 7807 1461
rect 20713 1458 20779 1461
rect 3693 1456 4354 1458
rect 3693 1400 3698 1456
rect 3754 1400 4354 1456
rect 3693 1398 4354 1400
rect 3693 1395 3759 1398
rect 4294 1186 4354 1398
rect 7741 1456 20779 1458
rect 7741 1400 7746 1456
rect 7802 1400 20718 1456
rect 20774 1400 20779 1456
rect 7741 1398 20779 1400
rect 7741 1395 7807 1398
rect 20713 1395 20779 1398
rect 21357 1458 21423 1461
rect 23473 1458 23539 1461
rect 21357 1456 23539 1458
rect 21357 1400 21362 1456
rect 21418 1400 23478 1456
rect 23534 1400 23539 1456
rect 21357 1398 23539 1400
rect 21357 1395 21423 1398
rect 23473 1395 23539 1398
rect 9029 1322 9095 1325
rect 22277 1322 22343 1325
rect 9029 1320 22343 1322
rect 9029 1264 9034 1320
rect 9090 1264 22282 1320
rect 22338 1264 22343 1320
rect 9029 1262 22343 1264
rect 9029 1259 9095 1262
rect 22277 1259 22343 1262
rect 18321 1186 18387 1189
rect 4294 1184 18387 1186
rect 4294 1128 18326 1184
rect 18382 1128 18387 1184
rect 4294 1126 18387 1128
rect 18321 1123 18387 1126
rect 5257 1050 5323 1053
rect 19333 1050 19399 1053
rect 5257 1048 19399 1050
rect 5257 992 5262 1048
rect 5318 992 19338 1048
rect 19394 992 19399 1048
rect 5257 990 19399 992
rect 5257 987 5323 990
rect 19333 987 19399 990
rect 0 914 480 944
rect 4705 914 4771 917
rect 0 912 4771 914
rect 0 856 4710 912
rect 4766 856 4771 912
rect 0 854 4771 856
rect 0 824 480 854
rect 4705 851 4771 854
rect 7925 914 7991 917
rect 22001 914 22067 917
rect 7925 912 22067 914
rect 7925 856 7930 912
rect 7986 856 22006 912
rect 22062 856 22067 912
rect 7925 854 22067 856
rect 7925 851 7991 854
rect 22001 851 22067 854
rect 15837 778 15903 781
rect 1166 776 15903 778
rect 1166 720 15842 776
rect 15898 720 15903 776
rect 1166 718 15903 720
rect 0 370 480 400
rect 1166 370 1226 718
rect 15837 715 15903 718
rect 2865 642 2931 645
rect 18137 642 18203 645
rect 2865 640 18203 642
rect 2865 584 2870 640
rect 2926 584 18142 640
rect 18198 584 18203 640
rect 2865 582 18203 584
rect 2865 579 2931 582
rect 18137 579 18203 582
rect 2957 506 3023 509
rect 18229 506 18295 509
rect 2957 504 18295 506
rect 2957 448 2962 504
rect 3018 448 18234 504
rect 18290 448 18295 504
rect 2957 446 18295 448
rect 2957 443 3023 446
rect 18229 443 18295 446
rect 0 310 1226 370
rect 0 280 480 310
rect 10041 234 10107 237
rect 24669 234 24735 237
rect 10041 232 24735 234
rect 10041 176 10046 232
rect 10102 176 24674 232
rect 24730 176 24735 232
rect 10041 174 24735 176
rect 10041 171 10107 174
rect 24669 171 24735 174
rect 8937 98 9003 101
rect 26417 98 26483 101
rect 8937 96 26483 98
rect 8937 40 8942 96
rect 8998 40 26422 96
rect 26478 40 26483 96
rect 8937 38 26483 40
rect 8937 35 9003 38
rect 26417 35 26483 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 9812 24712 9876 24716
rect 9812 24656 9862 24712
rect 9862 24656 9876 24712
rect 9812 24652 9876 24656
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 2636 24108 2700 24172
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 2636 21448 2700 21452
rect 2636 21392 2686 21448
rect 2686 21392 2700 21448
rect 2636 21388 2700 21392
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 9812 20224 9876 20228
rect 9812 20168 9862 20224
rect 9862 20168 9876 20224
rect 9812 20164 9876 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 15332 16008 15396 16012
rect 15332 15952 15346 16008
rect 15346 15952 15396 16008
rect 15332 15948 15396 15952
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 15332 10916 15396 10980
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 10916 9208 10980 9212
rect 10916 9152 10930 9208
rect 10930 9152 10980 9208
rect 10916 9148 10980 9152
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 18092 7380 18156 7444
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 9444 5808 9508 5812
rect 9444 5752 9494 5808
rect 9494 5752 9508 5808
rect 9444 5748 9508 5752
rect 16620 5748 16684 5812
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 1900 5128 1964 5132
rect 1900 5072 1914 5128
rect 1914 5072 1964 5128
rect 1900 5068 1964 5072
rect 10916 5068 10980 5132
rect 22324 5068 22388 5132
rect 9628 4932 9692 4996
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 8156 4040 8220 4044
rect 8156 3984 8206 4040
rect 8206 3984 8220 4040
rect 8156 3980 8220 3984
rect 20116 3904 20180 3908
rect 20116 3848 20130 3904
rect 20130 3848 20180 3904
rect 20116 3844 20180 3848
rect 20484 3980 20548 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 17724 3708 17788 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 6132 2620 6196 2684
rect 18092 2620 18156 2684
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 2636 1668 2700 1732
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 2635 24172 2701 24173
rect 2635 24108 2636 24172
rect 2700 24108 2701 24172
rect 2635 24107 2701 24108
rect 2638 21453 2698 24107
rect 5610 23968 5931 24992
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 9811 24716 9877 24717
rect 9811 24652 9812 24716
rect 9876 24652 9877 24716
rect 9811 24651 9877 24652
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 2635 21452 2701 21453
rect 2635 21388 2636 21452
rect 2700 21388 2701 21452
rect 2635 21387 2701 21388
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 9814 20229 9874 24651
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 9811 20228 9877 20229
rect 9811 20164 9812 20228
rect 9876 20164 9877 20228
rect 9811 20163 9877 20164
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 15331 16012 15397 16013
rect 15331 15948 15332 16012
rect 15396 15948 15397 16012
rect 15331 15947 15397 15948
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 15334 10981 15394 15947
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 15331 10980 15397 10981
rect 15331 10916 15332 10980
rect 15396 10916 15397 10980
rect 15331 10915 15397 10916
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 10915 9212 10981 9213
rect 10915 9148 10916 9212
rect 10980 9148 10981 9212
rect 10915 9147 10981 9148
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 8158 4045 8218 7022
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 9627 4996 9693 4997
rect 9627 4932 9628 4996
rect 9692 4932 9693 4996
rect 9627 4931 9693 4932
rect 9630 4538 9690 4931
rect 10277 4928 10597 5952
rect 10918 5133 10978 9147
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 18091 7444 18157 7445
rect 18091 7380 18092 7444
rect 18156 7380 18157 7444
rect 18091 7379 18157 7380
rect 18094 7258 18154 7379
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 10915 5132 10981 5133
rect 10915 5068 10916 5132
rect 10980 5068 10981 5132
rect 10915 5067 10981 5068
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 8155 4044 8221 4045
rect 8155 3980 8156 4044
rect 8220 3980 8221 4044
rect 8155 3979 8221 3980
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 6134 2685 6194 3622
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 6131 2684 6197 2685
rect 6131 2620 6132 2684
rect 6196 2620 6197 2684
rect 6131 2619 6197 2620
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2128 10597 2688
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 18094 2685 18154 7022
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 20486 4045 20546 4302
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 20115 3908 20181 3909
rect 20115 3844 20116 3908
rect 20180 3844 20181 3908
rect 20115 3843 20181 3844
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 18091 2684 18157 2685
rect 18091 2620 18092 2684
rect 18156 2620 18157 2684
rect 18091 2619 18157 2620
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2128 19930 2688
rect 20118 1818 20178 3843
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 8070 7022 8306 7258
rect 1814 5132 2050 5218
rect 1814 5068 1900 5132
rect 1900 5068 1964 5132
rect 1964 5068 2050 5132
rect 1814 4982 2050 5068
rect 9358 5812 9594 5898
rect 9358 5748 9444 5812
rect 9444 5748 9508 5812
rect 9508 5748 9594 5812
rect 9358 5662 9594 5748
rect 18006 7022 18242 7258
rect 16534 5812 16770 5898
rect 16534 5748 16620 5812
rect 16620 5748 16684 5812
rect 16684 5748 16770 5812
rect 16534 5662 16770 5748
rect 9542 4302 9778 4538
rect 6046 3622 6282 3858
rect 17638 3772 17874 3858
rect 17638 3708 17724 3772
rect 17724 3708 17788 3772
rect 17788 3708 17874 3772
rect 17638 3622 17874 3708
rect 22238 5132 22474 5218
rect 22238 5068 22324 5132
rect 22324 5068 22388 5132
rect 22388 5068 22474 5132
rect 22238 4982 22474 5068
rect 20398 4302 20634 4538
rect 2550 1732 2786 1818
rect 2550 1668 2636 1732
rect 2636 1668 2700 1732
rect 2700 1668 2786 1732
rect 2550 1582 2786 1668
rect 20030 1582 20266 1818
<< metal5 >>
rect 8028 7258 18284 7300
rect 8028 7022 8070 7258
rect 8306 7022 18006 7258
rect 18242 7022 18284 7258
rect 8028 6980 18284 7022
rect 9316 5898 16812 5940
rect 9316 5662 9358 5898
rect 9594 5662 16534 5898
rect 16770 5662 16812 5898
rect 9316 5620 16812 5662
rect 1772 5218 22516 5260
rect 1772 4982 1814 5218
rect 2050 4982 22238 5218
rect 22474 4982 22516 5218
rect 1772 4940 22516 4982
rect 9500 4538 20676 4580
rect 9500 4302 9542 4538
rect 9778 4302 20398 4538
rect 20634 4302 20676 4538
rect 9500 4260 20676 4302
rect 6004 3858 17916 3900
rect 6004 3622 6046 3858
rect 6282 3622 17638 3858
rect 17874 3622 17916 3858
rect 6004 3580 17916 3622
rect 2508 1818 20308 1860
rect 2508 1582 2550 1818
rect 2786 1582 20030 1818
rect 20266 1582 20308 1818
rect 2508 1540 20308 1582
use sky130_fd_sc_hd__fill_2  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_29
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_34
timestamp 1604681595
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37
timestamp 1604681595
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68
timestamp 1604681595
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _103_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1604681595
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1604681595
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12696 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_146
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_176
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_167
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1604681595
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1604681595
transform 1 0 20608 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_217
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1604681595
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_224
timestamp 1604681595
transform 1 0 21712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_229
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_236
timestamp 1604681595
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 1604681595
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1604681595
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_76
timestamp 1604681595
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17112 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18124 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1604681595
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1604681595
transform 1 0 17940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1604681595
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 21804 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_223
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22540 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_231
timestamp 1604681595
transform 1 0 22356 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_235
timestamp 1604681595
transform 1 0 22724 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_259
timestamp 1604681595
transform 1 0 24932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1604681595
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1604681595
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_96
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_100
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1604681595
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1604681595
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_226
timestamp 1604681595
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 22264 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_234
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_238 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1604681595
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_25
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_38
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5428 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1604681595
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_107
timestamp 1604681595
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_125
timestamp 1604681595
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_173
timestamp 1604681595
transform 1 0 17020 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1604681595
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 21160 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_222
timestamp 1604681595
transform 1 0 21528 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_226
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_234
timestamp 1604681595
transform 1 0 22632 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_246
timestamp 1604681595
transform 1 0 23736 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1604681595
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_10
timestamp 1604681595
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3956 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1604681595
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_46
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_84
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1604681595
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12880 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_137
timestamp 1604681595
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17664 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1604681595
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1604681595
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_214
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_218
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_230
timestamp 1604681595
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_234
timestamp 1604681595
transform 1 0 22632 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_242
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_249
timestamp 1604681595
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1604681595
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_265
timestamp 1604681595
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_20
timestamp 1604681595
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1472 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1604681595
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_25
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1604681595
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_31
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_40
timestamp 1604681595
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1604681595
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1604681595
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1604681595
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_107
timestamp 1604681595
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_119
timestamp 1604681595
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1604681595
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12696 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1604681595
transform 1 0 14536 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15732 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1604681595
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1604681595
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_168
timestamp 1604681595
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1604681595
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1604681595
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_209
timestamp 1604681595
transform 1 0 20332 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_221
timestamp 1604681595
transform 1 0 21436 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_231
timestamp 1604681595
transform 1 0 22356 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_238
timestamp 1604681595
transform 1 0 23000 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_250
timestamp 1604681595
transform 1 0 24104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_233
timestamp 1604681595
transform 1 0 22540 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1564 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_25
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1604681595
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_113
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_139
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 18124 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_177
timestamp 1604681595
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1604681595
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1604681595
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1604681595
transform 1 0 3864 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1604681595
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13064 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_146
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_150
timestamp 1604681595
transform 1 0 14904 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_201
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_213
timestamp 1604681595
transform 1 0 20700 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1604681595
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_21
timestamp 1604681595
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 1604681595
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1604681595
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1604681595
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_120
timestamp 1604681595
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_198
timestamp 1604681595
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1604681595
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 5612 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_90
timestamp 1604681595
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_95
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12512 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14168 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1604681595
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_137
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_67
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1604681595
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_111
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_119
timestamp 1604681595
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1604681595
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_136
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_144
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_168
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1604681595
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_192
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_204
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1604681595
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_9
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_14
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6072 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1604681595
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1604681595
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1604681595
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_130
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1604681595
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1604681595
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_168
timestamp 1604681595
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_187
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_175
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_166
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1604681595
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_46
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_74
timestamp 1604681595
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604681595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_142
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1604681595
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_78
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1604681595
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1604681595
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_106
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12696 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_142
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1604681595
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_168
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_173
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_45
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_59
timestamp 1604681595
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1604681595
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_192
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1604681595
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1604681595
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_47
timestamp 1604681595
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604681595
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_109
timestamp 1604681595
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1604681595
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1604681595
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1604681595
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_143
timestamp 1604681595
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_139
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_176
timestamp 1604681595
transform 1 0 17296 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_189
timestamp 1604681595
transform 1 0 18492 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1604681595
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_255
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_6
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1604681595
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1604681595
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_56
timestamp 1604681595
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_52
timestamp 1604681595
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_65
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13156 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_151
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_176
timestamp 1604681595
transform 1 0 17296 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 24380 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1604681595
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_96
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1604681595
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_158
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_162
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16468 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1604681595
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1604681595
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1604681595
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4140 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_24
timestamp 1604681595
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_28
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_49
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_89
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1604681595
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1604681595
transform 1 0 14812 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_153
timestamp 1604681595
transform 1 0 15180 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_205
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_217
timestamp 1604681595
transform 1 0 21068 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1604681595
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1604681595
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8188 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_83
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_87
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 11776 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_147
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_167
timestamp 1604681595
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_186
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_198
timestamp 1604681595
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1604681595
transform 1 0 21436 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1604681595
transform 1 0 22540 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_245
timestamp 1604681595
transform 1 0 23644 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_257
timestamp 1604681595
transform 1 0 24748 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_269
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1564 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_21
timestamp 1604681595
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_25
timestamp 1604681595
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_29
timestamp 1604681595
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_75
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1604681595
transform 1 0 8740 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1604681595
transform 1 0 9108 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1604681595
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_133
timestamp 1604681595
transform 1 0 13340 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1604681595
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_13
timestamp 1604681595
transform 1 0 2300 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1604681595
transform 1 0 4324 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1604681595
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_77
timestamp 1604681595
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8096 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_89
timestamp 1604681595
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1604681595
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_104
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_112
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_112
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_120
timestamp 1604681595
transform 1 0 12144 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_136
timestamp 1604681595
transform 1 0 13616 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_144
timestamp 1604681595
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_140
timestamp 1604681595
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1604681595
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_174
timestamp 1604681595
transform 1 0 17112 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_171
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_187
timestamp 1604681595
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_175
timestamp 1604681595
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_199
timestamp 1604681595
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11960 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1604681595
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_113
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_170
timestamp 1604681595
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_182
timestamp 1604681595
transform 1 0 17848 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_194
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1604681595
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_16
timestamp 1604681595
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_37
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1604681595
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 5244 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1604681595
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5796 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1604681595
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_100
timestamp 1604681595
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_96
timestamp 1604681595
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_120
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_133
timestamp 1604681595
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_175
timestamp 1604681595
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_187
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_199
timestamp 1604681595
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1604681595
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_13
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_16
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1604681595
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1604681595
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_50
timestamp 1604681595
transform 1 0 5704 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_54
timestamp 1604681595
transform 1 0 6072 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_65
timestamp 1604681595
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1604681595
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_103
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_167
timestamp 1604681595
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 1604681595
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1604681595
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_70
timestamp 1604681595
transform 1 0 7544 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_75
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1604681595
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp 1604681595
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_106
timestamp 1604681595
transform 1 0 10856 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_16
timestamp 1604681595
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_12
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1604681595
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_20
timestamp 1604681595
transform 1 0 2944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_24
timestamp 1604681595
transform 1 0 3312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_38
timestamp 1604681595
transform 1 0 4600 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_40
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_46
timestamp 1604681595
transform 1 0 5336 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_42
timestamp 1604681595
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5428 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1604681595
transform 1 0 8648 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_90
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_95
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_113
timestamp 1604681595
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1604681595
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604681595
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_132
timestamp 1604681595
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_128
timestamp 1604681595
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1604681595
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_139
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14076 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_150
timestamp 1604681595
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_157
timestamp 1604681595
transform 1 0 15548 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_158
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_163
timestamp 1604681595
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_164
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 16284 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1604681595
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1604681595
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_192
timestamp 1604681595
transform 1 0 18768 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1604681595
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_12
timestamp 1604681595
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_16
timestamp 1604681595
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_20
timestamp 1604681595
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_24
timestamp 1604681595
transform 1 0 3312 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_38
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8096 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_68
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1604681595
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_92
timestamp 1604681595
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_96
timestamp 1604681595
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 11868 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_109
timestamp 1604681595
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1604681595
transform 1 0 12788 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_133
timestamp 1604681595
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_157
timestamp 1604681595
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_170
timestamp 1604681595
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_174
timestamp 1604681595
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1604681595
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_36
timestamp 1604681595
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4784 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1604681595
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_67
timestamp 1604681595
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_71
timestamp 1604681595
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_102
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11132 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_120
timestamp 1604681595
transform 1 0 12144 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_132
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_170
timestamp 1604681595
transform 1 0 16744 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_182
timestamp 1604681595
transform 1 0 17848 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604681595
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_20
timestamp 1604681595
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3864 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_24
timestamp 1604681595
transform 1 0 3312 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_46
timestamp 1604681595
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_50
timestamp 1604681595
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_54
timestamp 1604681595
transform 1 0 6072 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_58
timestamp 1604681595
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_65
timestamp 1604681595
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 1604681595
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_82
timestamp 1604681595
transform 1 0 8648 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1604681595
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_100
timestamp 1604681595
transform 1 0 10304 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_131
timestamp 1604681595
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 15180 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_151
timestamp 1604681595
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1604681595
transform 1 0 15364 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1604681595
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1604681595
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_173
timestamp 1604681595
transform 1 0 17020 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_181
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_188
timestamp 1604681595
transform 1 0 18400 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1604681595
transform 1 0 19320 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_222
timestamp 1604681595
transform 1 0 21528 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_230
timestamp 1604681595
transform 1 0 22264 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_233
timestamp 1604681595
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_241
timestamp 1604681595
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_13
timestamp 1604681595
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_17
timestamp 1604681595
transform 1 0 2668 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_22
timestamp 1604681595
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_26
timestamp 1604681595
transform 1 0 3496 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_48
timestamp 1604681595
transform 1 0 5520 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_59
timestamp 1604681595
transform 1 0 6532 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7268 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_38_83
timestamp 1604681595
transform 1 0 8740 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_102
timestamp 1604681595
transform 1 0 10488 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_107
timestamp 1604681595
transform 1 0 10948 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1604681595
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_143
timestamp 1604681595
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16284 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_147
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_157
timestamp 1604681595
transform 1 0 15548 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17848 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_171
timestamp 1604681595
transform 1 0 16836 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_179
timestamp 1604681595
transform 1 0 17572 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1604681595
transform 1 0 18400 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_200
timestamp 1604681595
transform 1 0 19504 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 21344 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_222
timestamp 1604681595
transform 1 0 21528 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_230
timestamp 1604681595
transform 1 0 22264 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1604681595
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_249
timestamp 1604681595
transform 1 0 24012 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_261
timestamp 1604681595
transform 1 0 25116 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1604681595
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_16
timestamp 1604681595
transform 1 0 2576 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_12
timestamp 1604681595
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_29
timestamp 1604681595
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_33
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4324 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_40_50
timestamp 1604681595
transform 1 0 5704 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_46
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_58
timestamp 1604681595
transform 1 0 6440 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_65
timestamp 1604681595
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_69
timestamp 1604681595
transform 1 0 7452 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_79
timestamp 1604681595
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_83
timestamp 1604681595
transform 1 0 8740 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_93
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_97
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_111
timestamp 1604681595
transform 1 0 11316 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_123
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_115
timestamp 1604681595
transform 1 0 11684 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_127
timestamp 1604681595
transform 1 0 12788 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13524 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp 1604681595
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_156
timestamp 1604681595
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_160
timestamp 1604681595
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1604681595
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_172
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_168
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_182
timestamp 1604681595
transform 1 0 17848 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_194
timestamp 1604681595
transform 1 0 18952 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_217
timestamp 1604681595
transform 1 0 21068 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_229
timestamp 1604681595
transform 1 0 22172 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_249
timestamp 1604681595
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1604681595
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_25
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_29
timestamp 1604681595
transform 1 0 3772 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_40
timestamp 1604681595
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_73
timestamp 1604681595
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1604681595
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_85
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_97
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1604681595
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_105
timestamp 1604681595
transform 1 0 10764 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 14076 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 12972 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_127
timestamp 1604681595
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_131
timestamp 1604681595
transform 1 0 13156 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_139
timestamp 1604681595
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 15456 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 15272 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_151
timestamp 1604681595
transform 1 0 14996 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_160
timestamp 1604681595
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_164
timestamp 1604681595
transform 1 0 16192 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_170
timestamp 1604681595
transform 1 0 16744 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_175
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1604681595
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_13
timestamp 1604681595
transform 1 0 2300 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_25
timestamp 1604681595
transform 1 0 3404 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_52
timestamp 1604681595
transform 1 0 5888 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_110
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1604681595
transform 1 0 11592 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 13524 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_129
timestamp 1604681595
transform 1 0 12972 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1604681595
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_160
timestamp 1604681595
transform 1 0 15824 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_172
timestamp 1604681595
transform 1 0 16928 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_184
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 27618 0 27674 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 9 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 4360 480 4480 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 139 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
