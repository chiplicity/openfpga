magic
tech sky130A
magscale 1 2
timestamp 1609021633
<< locali >>
rect 23581 20859 23615 22049
rect 12265 18071 12299 18377
rect 4445 16643 4479 16745
rect 12265 15895 12299 16065
rect 23581 9707 23615 19261
rect 23581 9367 23615 9537
<< viali >>
rect 7757 22185 7791 22219
rect 8125 22185 8159 22219
rect 6377 22117 6411 22151
rect 6929 22117 6963 22151
rect 7665 22117 7699 22151
rect 10609 22117 10643 22151
rect 13369 22117 13403 22151
rect 14473 22117 14507 22151
rect 17785 22117 17819 22151
rect 4353 22049 4387 22083
rect 4721 22049 4755 22083
rect 5181 22049 5215 22083
rect 5549 22049 5583 22083
rect 6285 22049 6319 22083
rect 10149 22049 10183 22083
rect 12449 22049 12483 22083
rect 13277 22049 13311 22083
rect 14381 22049 14415 22083
rect 14841 22049 14875 22083
rect 15209 22049 15243 22083
rect 15485 22049 15519 22083
rect 15853 22049 15887 22083
rect 16221 22049 16255 22083
rect 17877 22049 17911 22083
rect 23581 22049 23615 22083
rect 2697 21981 2731 22015
rect 6469 21981 6503 22015
rect 7849 21981 7883 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 13553 21981 13587 22015
rect 14657 21981 14691 22015
rect 17969 21981 18003 22015
rect 4905 21913 4939 21947
rect 12909 21913 12943 21947
rect 2329 21845 2363 21879
rect 4537 21845 4571 21879
rect 5365 21845 5399 21879
rect 5733 21845 5767 21879
rect 5917 21845 5951 21879
rect 7297 21845 7331 21879
rect 9781 21845 9815 21879
rect 14013 21845 14047 21879
rect 15025 21845 15059 21879
rect 15669 21845 15703 21879
rect 16037 21845 16071 21879
rect 17417 21845 17451 21879
rect 18337 21845 18371 21879
rect 2053 21641 2087 21675
rect 4261 21641 4295 21675
rect 6193 21641 6227 21675
rect 6837 21641 6871 21675
rect 7573 21641 7607 21675
rect 13829 21641 13863 21675
rect 17693 21641 17727 21675
rect 22477 21641 22511 21675
rect 2421 21573 2455 21607
rect 12173 21573 12207 21607
rect 22845 21573 22879 21607
rect 4537 21505 4571 21539
rect 8125 21505 8159 21539
rect 8401 21505 8435 21539
rect 15945 21505 15979 21539
rect 17325 21505 17359 21539
rect 18061 21505 18095 21539
rect 18705 21505 18739 21539
rect 1869 21437 1903 21471
rect 2237 21437 2271 21471
rect 2605 21437 2639 21471
rect 4077 21437 4111 21471
rect 6009 21437 6043 21471
rect 6377 21437 6411 21471
rect 7021 21437 7055 21471
rect 9045 21437 9079 21471
rect 10517 21437 10551 21471
rect 11989 21437 12023 21471
rect 12449 21437 12483 21471
rect 13921 21437 13955 21471
rect 15761 21437 15795 21471
rect 16221 21437 16255 21471
rect 17509 21437 17543 21471
rect 18521 21437 18555 21471
rect 19441 21437 19475 21471
rect 22293 21437 22327 21471
rect 22661 21437 22695 21471
rect 23029 21437 23063 21471
rect 2872 21369 2906 21403
rect 4804 21369 4838 21403
rect 7481 21369 7515 21403
rect 9312 21369 9346 21403
rect 10762 21369 10796 21403
rect 12716 21369 12750 21403
rect 14188 21369 14222 21403
rect 3985 21301 4019 21335
rect 5917 21301 5951 21335
rect 6561 21301 6595 21335
rect 7205 21301 7239 21335
rect 7941 21301 7975 21335
rect 8033 21301 8067 21335
rect 10425 21301 10459 21335
rect 11897 21301 11931 21335
rect 15301 21301 15335 21335
rect 15393 21301 15427 21335
rect 15853 21301 15887 21335
rect 16405 21301 16439 21335
rect 16681 21301 16715 21335
rect 17049 21301 17083 21335
rect 17141 21301 17175 21335
rect 22201 21301 22235 21335
rect 1777 21097 1811 21131
rect 3617 21097 3651 21131
rect 3893 21097 3927 21131
rect 5457 21097 5491 21131
rect 5917 21097 5951 21131
rect 6101 21097 6135 21131
rect 7573 21097 7607 21131
rect 9321 21097 9355 21131
rect 11069 21097 11103 21131
rect 11621 21097 11655 21131
rect 13093 21097 13127 21131
rect 14565 21097 14599 21131
rect 16681 21097 16715 21131
rect 18153 21097 18187 21131
rect 22845 21097 22879 21131
rect 4322 21029 4356 21063
rect 5733 21029 5767 21063
rect 6460 21029 6494 21063
rect 7932 21029 7966 21063
rect 11980 21029 12014 21063
rect 13452 21029 13486 21063
rect 14749 21029 14783 21063
rect 17018 21029 17052 21063
rect 18490 21029 18524 21063
rect 22201 21029 22235 21063
rect 1593 20961 1627 20995
rect 1961 20961 1995 20995
rect 2228 20961 2262 20995
rect 3433 20961 3467 20995
rect 5549 20961 5583 20995
rect 9689 20961 9723 20995
rect 9945 20961 9979 20995
rect 11161 20961 11195 20995
rect 14933 20961 14967 20995
rect 15568 20961 15602 20995
rect 22293 20961 22327 20995
rect 22661 20961 22695 20995
rect 4077 20893 4111 20927
rect 6200 20893 6234 20927
rect 7665 20893 7699 20927
rect 11713 20893 11747 20927
rect 13185 20893 13219 20927
rect 15117 20893 15151 20927
rect 15301 20893 15335 20927
rect 16773 20893 16807 20927
rect 18245 20893 18279 20927
rect 3341 20825 3375 20859
rect 22477 20825 22511 20859
rect 23581 20825 23615 20859
rect 1501 20757 1535 20791
rect 9045 20757 9079 20791
rect 11345 20757 11379 20791
rect 19625 20757 19659 20791
rect 23121 20757 23155 20791
rect 2973 20553 3007 20587
rect 4905 20553 4939 20587
rect 6561 20553 6595 20587
rect 10701 20553 10735 20587
rect 13829 20553 13863 20587
rect 15761 20553 15795 20587
rect 16681 20553 16715 20587
rect 19533 20553 19567 20587
rect 22477 20553 22511 20587
rect 1593 20417 1627 20451
rect 3709 20417 3743 20451
rect 4353 20417 4387 20451
rect 4537 20417 4571 20451
rect 5181 20417 5215 20451
rect 6837 20417 6871 20451
rect 9321 20417 9355 20451
rect 11345 20417 11379 20451
rect 16405 20417 16439 20451
rect 17233 20417 17267 20451
rect 18061 20417 18095 20451
rect 20085 20417 20119 20451
rect 3433 20349 3467 20383
rect 4261 20349 4295 20383
rect 4721 20349 4755 20383
rect 5448 20349 5482 20383
rect 7113 20349 7147 20383
rect 7380 20349 7414 20383
rect 8585 20349 8619 20383
rect 9588 20349 9622 20383
rect 11161 20349 11195 20383
rect 11989 20349 12023 20383
rect 12449 20349 12483 20383
rect 12716 20349 12750 20383
rect 13921 20349 13955 20383
rect 14381 20349 14415 20383
rect 16221 20349 16255 20383
rect 17141 20349 17175 20383
rect 17509 20349 17543 20383
rect 18328 20349 18362 20383
rect 22293 20349 22327 20383
rect 1860 20281 1894 20315
rect 3525 20281 3559 20315
rect 9045 20281 9079 20315
rect 11253 20281 11287 20315
rect 14626 20281 14660 20315
rect 16313 20281 16347 20315
rect 17049 20281 17083 20315
rect 19901 20281 19935 20315
rect 3065 20213 3099 20247
rect 3893 20213 3927 20247
rect 8493 20213 8527 20247
rect 8769 20213 8803 20247
rect 10793 20213 10827 20247
rect 12173 20213 12207 20247
rect 14105 20213 14139 20247
rect 15853 20213 15887 20247
rect 17693 20213 17727 20247
rect 19441 20213 19475 20247
rect 19993 20213 20027 20247
rect 22109 20213 22143 20247
rect 22661 20213 22695 20247
rect 22937 20213 22971 20247
rect 2973 20009 3007 20043
rect 4445 20009 4479 20043
rect 4905 20009 4939 20043
rect 5733 20009 5767 20043
rect 8769 20009 8803 20043
rect 9689 20009 9723 20043
rect 13829 20009 13863 20043
rect 14197 20009 14231 20043
rect 14565 20009 14599 20043
rect 15117 20009 15151 20043
rect 15761 20009 15795 20043
rect 16129 20009 16163 20043
rect 22477 20009 22511 20043
rect 22845 20009 22879 20043
rect 1860 19941 1894 19975
rect 4537 19941 4571 19975
rect 6101 19941 6135 19975
rect 7012 19941 7046 19975
rect 10057 19941 10091 19975
rect 10977 19941 11011 19975
rect 16589 19941 16623 19975
rect 17325 19941 17359 19975
rect 17868 19941 17902 19975
rect 21465 19941 21499 19975
rect 1593 19873 1627 19907
rect 3433 19873 3467 19907
rect 5273 19873 5307 19907
rect 6653 19873 6687 19907
rect 8217 19873 8251 19907
rect 9137 19873 9171 19907
rect 10885 19873 10919 19907
rect 12909 19873 12943 19907
rect 13737 19873 13771 19907
rect 15669 19873 15703 19907
rect 16497 19873 16531 19907
rect 16957 19873 16991 19907
rect 19625 19873 19659 19907
rect 21373 19873 21407 19907
rect 21925 19873 21959 19907
rect 22293 19873 22327 19907
rect 22661 19873 22695 19907
rect 3525 19805 3559 19839
rect 3709 19805 3743 19839
rect 4721 19805 4755 19839
rect 5365 19805 5399 19839
rect 5457 19805 5491 19839
rect 6193 19805 6227 19839
rect 6285 19805 6319 19839
rect 6745 19805 6779 19839
rect 9229 19805 9263 19839
rect 9413 19805 9447 19839
rect 10149 19805 10183 19839
rect 10241 19805 10275 19839
rect 11161 19805 11195 19839
rect 13001 19805 13035 19839
rect 13093 19805 13127 19839
rect 13921 19805 13955 19839
rect 14657 19805 14691 19839
rect 14749 19805 14783 19839
rect 15853 19805 15887 19839
rect 16681 19805 16715 19839
rect 17601 19805 17635 19839
rect 19717 19805 19751 19839
rect 19901 19805 19935 19839
rect 21557 19805 21591 19839
rect 8401 19737 8435 19771
rect 8677 19737 8711 19771
rect 11437 19737 11471 19771
rect 13369 19737 13403 19771
rect 15301 19737 15335 19771
rect 3065 19669 3099 19703
rect 4077 19669 4111 19703
rect 8125 19669 8159 19703
rect 10517 19669 10551 19703
rect 12541 19669 12575 19703
rect 17141 19669 17175 19703
rect 18981 19669 19015 19703
rect 19257 19669 19291 19703
rect 21005 19669 21039 19703
rect 22109 19669 22143 19703
rect 23121 19669 23155 19703
rect 2053 19465 2087 19499
rect 13829 19465 13863 19499
rect 22845 19465 22879 19499
rect 2421 19397 2455 19431
rect 15669 19397 15703 19431
rect 3157 19329 3191 19363
rect 3985 19329 4019 19363
rect 5089 19329 5123 19363
rect 5917 19329 5951 19363
rect 7389 19329 7423 19363
rect 7988 19329 8022 19363
rect 8128 19329 8162 19363
rect 14565 19329 14599 19363
rect 15393 19329 15427 19363
rect 16221 19329 16255 19363
rect 1869 19261 1903 19295
rect 2237 19261 2271 19295
rect 3801 19261 3835 19295
rect 5825 19261 5859 19295
rect 6193 19261 6227 19295
rect 7665 19261 7699 19295
rect 8401 19261 8435 19295
rect 9781 19261 9815 19295
rect 10057 19261 10091 19295
rect 10324 19261 10358 19295
rect 12449 19261 12483 19295
rect 15209 19261 15243 19295
rect 16504 19261 16538 19295
rect 16764 19261 16798 19295
rect 18245 19261 18279 19295
rect 19717 19261 19751 19295
rect 21189 19261 21223 19295
rect 22661 19261 22695 19295
rect 23581 19261 23615 19295
rect 5733 19193 5767 19227
rect 11713 19193 11747 19227
rect 12716 19193 12750 19227
rect 14381 19193 14415 19227
rect 16037 19193 16071 19227
rect 18512 19193 18546 19227
rect 19984 19193 20018 19227
rect 21456 19193 21490 19227
rect 2605 19125 2639 19159
rect 2973 19125 3007 19159
rect 3065 19125 3099 19159
rect 3433 19125 3467 19159
rect 3893 19125 3927 19159
rect 4537 19125 4571 19159
rect 4905 19125 4939 19159
rect 4997 19125 5031 19159
rect 5365 19125 5399 19159
rect 6377 19125 6411 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 7297 19125 7331 19159
rect 9505 19125 9539 19159
rect 9689 19125 9723 19159
rect 11437 19125 11471 19159
rect 14013 19125 14047 19159
rect 14473 19125 14507 19159
rect 14841 19125 14875 19159
rect 15301 19125 15335 19159
rect 16129 19125 16163 19159
rect 17877 19125 17911 19159
rect 19625 19125 19659 19159
rect 21097 19125 21131 19159
rect 22569 19125 22603 19159
rect 23029 19125 23063 19159
rect 3065 18921 3099 18955
rect 3157 18921 3191 18955
rect 4261 18921 4295 18955
rect 4905 18921 4939 18955
rect 5273 18921 5307 18955
rect 6561 18921 6595 18955
rect 7021 18921 7055 18955
rect 9229 18921 9263 18955
rect 11529 18921 11563 18955
rect 13001 18921 13035 18955
rect 15301 18921 15335 18955
rect 15669 18921 15703 18955
rect 18521 18921 18555 18955
rect 20361 18921 20395 18955
rect 22293 18921 22327 18955
rect 22753 18921 22787 18955
rect 4813 18853 4847 18887
rect 9413 18853 9447 18887
rect 13338 18853 13372 18887
rect 21158 18853 21192 18887
rect 22845 18853 22879 18887
rect 1685 18785 1719 18819
rect 1952 18785 1986 18819
rect 3525 18785 3559 18819
rect 4077 18785 4111 18819
rect 5641 18785 5675 18819
rect 6101 18785 6135 18819
rect 6929 18785 6963 18819
rect 8125 18785 8159 18819
rect 10425 18785 10459 18819
rect 11621 18785 11655 18819
rect 11888 18785 11922 18819
rect 14565 18785 14599 18819
rect 15761 18785 15795 18819
rect 16129 18785 16163 18819
rect 16589 18785 16623 18819
rect 17325 18785 17359 18819
rect 18981 18785 19015 18819
rect 19248 18785 19282 18819
rect 20453 18785 20487 18819
rect 3617 18717 3651 18751
rect 3709 18717 3743 18751
rect 5089 18717 5123 18751
rect 5733 18717 5767 18751
rect 5825 18717 5859 18751
rect 7113 18717 7147 18751
rect 7389 18717 7423 18751
rect 7712 18717 7746 18751
rect 7895 18717 7929 18751
rect 9689 18717 9723 18751
rect 10012 18717 10046 18751
rect 10195 18717 10229 18751
rect 13093 18717 13127 18751
rect 15945 18717 15979 18751
rect 16912 18717 16946 18751
rect 17095 18717 17129 18751
rect 20913 18717 20947 18751
rect 22937 18717 22971 18751
rect 6285 18649 6319 18683
rect 14749 18649 14783 18683
rect 22385 18649 22419 18683
rect 4445 18581 4479 18615
rect 14473 18581 14507 18615
rect 15117 18581 15151 18615
rect 16313 18581 16347 18615
rect 18429 18581 18463 18615
rect 20637 18581 20671 18615
rect 3157 18377 3191 18411
rect 4629 18377 4663 18411
rect 6469 18377 6503 18411
rect 10793 18377 10827 18411
rect 11621 18377 11655 18411
rect 12265 18377 12299 18411
rect 12449 18377 12483 18411
rect 16313 18377 16347 18411
rect 17785 18377 17819 18411
rect 19993 18377 20027 18411
rect 20085 18377 20119 18411
rect 8309 18241 8343 18275
rect 8585 18241 8619 18275
rect 9324 18241 9358 18275
rect 11253 18241 11287 18275
rect 11345 18241 11379 18275
rect 1777 18173 1811 18207
rect 2044 18173 2078 18207
rect 3249 18173 3283 18207
rect 4813 18173 4847 18207
rect 5080 18173 5114 18207
rect 6285 18173 6319 18207
rect 6837 18173 6871 18207
rect 7104 18173 7138 18207
rect 8861 18173 8895 18207
rect 9597 18173 9631 18207
rect 11161 18173 11195 18207
rect 11805 18173 11839 18207
rect 3516 18105 3550 18139
rect 23029 18309 23063 18343
rect 13093 18241 13127 18275
rect 18613 18241 18647 18275
rect 20545 18241 20579 18275
rect 20637 18241 20671 18275
rect 13277 18173 13311 18207
rect 14933 18173 14967 18207
rect 16405 18173 16439 18207
rect 16661 18173 16695 18207
rect 20453 18173 20487 18207
rect 20913 18173 20947 18207
rect 21373 18173 21407 18207
rect 21640 18173 21674 18207
rect 22845 18173 22879 18207
rect 12817 18105 12851 18139
rect 13544 18105 13578 18139
rect 15200 18105 15234 18139
rect 18880 18105 18914 18139
rect 6193 18037 6227 18071
rect 8217 18037 8251 18071
rect 9327 18037 9361 18071
rect 10701 18037 10735 18071
rect 12265 18037 12299 18071
rect 12909 18037 12943 18071
rect 14657 18037 14691 18071
rect 21097 18037 21131 18071
rect 22753 18037 22787 18071
rect 8953 17833 8987 17867
rect 9689 17833 9723 17867
rect 10057 17833 10091 17867
rect 11805 17833 11839 17867
rect 14013 17833 14047 17867
rect 14105 17833 14139 17867
rect 14473 17833 14507 17867
rect 14933 17833 14967 17867
rect 16681 17833 16715 17867
rect 17509 17833 17543 17867
rect 19441 17833 19475 17867
rect 19809 17833 19843 17867
rect 22937 17833 22971 17867
rect 5080 17765 5114 17799
rect 8861 17765 8895 17799
rect 10149 17765 10183 17799
rect 12265 17765 12299 17799
rect 14565 17765 14599 17799
rect 15546 17765 15580 17799
rect 17601 17765 17635 17799
rect 21005 17765 21039 17799
rect 21097 17765 21131 17799
rect 21281 17765 21315 17799
rect 21824 17765 21858 17799
rect 2145 17697 2179 17731
rect 2412 17697 2446 17731
rect 4813 17697 4847 17731
rect 7288 17697 7322 17731
rect 9505 17697 9539 17731
rect 10885 17697 10919 17731
rect 12173 17697 12207 17731
rect 12900 17697 12934 17731
rect 15117 17697 15151 17731
rect 15301 17697 15335 17731
rect 17969 17697 18003 17731
rect 18236 17697 18270 17731
rect 20269 17697 20303 17731
rect 7021 17629 7055 17663
rect 9045 17629 9079 17663
rect 10241 17629 10275 17663
rect 10977 17629 11011 17663
rect 11069 17629 11103 17663
rect 12449 17629 12483 17663
rect 12633 17629 12667 17663
rect 14657 17629 14691 17663
rect 17785 17629 17819 17663
rect 19901 17629 19935 17663
rect 20085 17629 20119 17663
rect 21557 17629 21591 17663
rect 23121 17629 23155 17663
rect 8493 17561 8527 17595
rect 17141 17561 17175 17595
rect 19349 17561 19383 17595
rect 3525 17493 3559 17527
rect 6193 17493 6227 17527
rect 8401 17493 8435 17527
rect 9321 17493 9355 17527
rect 10517 17493 10551 17527
rect 20453 17493 20487 17527
rect 21465 17493 21499 17527
rect 4721 17289 4755 17323
rect 6285 17289 6319 17323
rect 6561 17289 6595 17323
rect 6837 17289 6871 17323
rect 8033 17289 8067 17323
rect 9597 17289 9631 17323
rect 9873 17289 9907 17323
rect 12081 17289 12115 17323
rect 13829 17289 13863 17323
rect 15393 17289 15427 17323
rect 19441 17289 19475 17323
rect 21557 17289 21591 17323
rect 1869 17153 1903 17187
rect 3341 17153 3375 17187
rect 4813 17153 4847 17187
rect 7389 17153 7423 17187
rect 10517 17153 10551 17187
rect 18061 17153 18095 17187
rect 20177 17153 20211 17187
rect 21189 17153 21223 17187
rect 22109 17153 22143 17187
rect 22845 17153 22879 17187
rect 22937 17153 22971 17187
rect 3608 17085 3642 17119
rect 5080 17085 5114 17119
rect 6469 17085 6503 17119
rect 7665 17085 7699 17119
rect 8217 17085 8251 17119
rect 10241 17085 10275 17119
rect 10701 17085 10735 17119
rect 12449 17085 12483 17119
rect 12716 17085 12750 17119
rect 14013 17085 14047 17119
rect 19901 17085 19935 17119
rect 20913 17085 20947 17119
rect 21925 17085 21959 17119
rect 22753 17085 22787 17119
rect 2136 17017 2170 17051
rect 7297 17017 7331 17051
rect 8484 17017 8518 17051
rect 9689 17017 9723 17051
rect 10968 17017 11002 17051
rect 14280 17017 14314 17051
rect 18328 17017 18362 17051
rect 19993 17017 20027 17051
rect 22017 17017 22051 17051
rect 3249 16949 3283 16983
rect 6193 16949 6227 16983
rect 7205 16949 7239 16983
rect 7849 16949 7883 16983
rect 10333 16949 10367 16983
rect 19533 16949 19567 16983
rect 20545 16949 20579 16983
rect 21005 16949 21039 16983
rect 22385 16949 22419 16983
rect 3065 16745 3099 16779
rect 3617 16745 3651 16779
rect 4445 16745 4479 16779
rect 4537 16745 4571 16779
rect 6653 16745 6687 16779
rect 9413 16745 9447 16779
rect 11161 16745 11195 16779
rect 14933 16745 14967 16779
rect 15301 16745 15335 16779
rect 17417 16745 17451 16779
rect 19073 16745 19107 16779
rect 19165 16745 19199 16779
rect 20453 16745 20487 16779
rect 21373 16745 21407 16779
rect 23121 16745 23155 16779
rect 1952 16677 1986 16711
rect 5080 16677 5114 16711
rect 10048 16677 10082 16711
rect 15936 16677 15970 16711
rect 20361 16677 20395 16711
rect 21802 16677 21836 16711
rect 1685 16609 1719 16643
rect 3525 16609 3559 16643
rect 4445 16609 4479 16643
rect 4721 16609 4755 16643
rect 6285 16609 6319 16643
rect 7196 16609 7230 16643
rect 8769 16609 8803 16643
rect 9229 16609 9263 16643
rect 11713 16609 11747 16643
rect 12173 16609 12207 16643
rect 13553 16609 13587 16643
rect 13820 16609 13854 16643
rect 15485 16609 15519 16643
rect 17601 16609 17635 16643
rect 17693 16609 17727 16643
rect 17960 16609 17994 16643
rect 19533 16609 19567 16643
rect 21189 16609 21223 16643
rect 21557 16609 21591 16643
rect 3709 16541 3743 16575
rect 4813 16541 4847 16575
rect 6929 16541 6963 16575
rect 8861 16541 8895 16575
rect 8953 16541 8987 16575
rect 9781 16541 9815 16575
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 15669 16541 15703 16575
rect 19625 16541 19659 16575
rect 19809 16541 19843 16575
rect 20637 16541 20671 16575
rect 3157 16473 3191 16507
rect 6193 16473 6227 16507
rect 8401 16473 8435 16507
rect 12541 16473 12575 16507
rect 19993 16473 20027 16507
rect 6469 16405 6503 16439
rect 8309 16405 8343 16439
rect 11345 16405 11379 16439
rect 17049 16405 17083 16439
rect 22937 16405 22971 16439
rect 3433 16201 3467 16235
rect 3525 16201 3559 16235
rect 5549 16201 5583 16235
rect 8309 16201 8343 16235
rect 9321 16201 9355 16235
rect 11437 16201 11471 16235
rect 13921 16201 13955 16235
rect 17049 16201 17083 16235
rect 19441 16201 19475 16235
rect 21189 16201 21223 16235
rect 4537 16133 4571 16167
rect 11345 16133 11379 16167
rect 3985 16065 4019 16099
rect 4077 16065 4111 16099
rect 5273 16065 5307 16099
rect 6193 16065 6227 16099
rect 8861 16065 8895 16099
rect 9828 16065 9862 16099
rect 10011 16065 10045 16099
rect 10241 16065 10275 16099
rect 11897 16065 11931 16099
rect 11989 16065 12023 16099
rect 12265 16065 12299 16099
rect 14473 16065 14507 16099
rect 15672 16065 15706 16099
rect 17693 16065 17727 16099
rect 20177 16065 20211 16099
rect 20913 16065 20947 16099
rect 21649 16065 21683 16099
rect 21833 16065 21867 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 2053 15997 2087 16031
rect 2320 15997 2354 16031
rect 3893 15997 3927 16031
rect 4353 15997 4387 16031
rect 5181 15997 5215 16031
rect 5917 15997 5951 16031
rect 6377 15997 6411 16031
rect 6837 15997 6871 16031
rect 8677 15997 8711 16031
rect 9137 15997 9171 16031
rect 9505 15997 9539 16031
rect 6009 15929 6043 15963
rect 7082 15929 7116 15963
rect 12449 15997 12483 16031
rect 15209 15997 15243 16031
rect 15945 15997 15979 16031
rect 17509 15997 17543 16031
rect 18061 15997 18095 16031
rect 22845 15997 22879 16031
rect 12694 15929 12728 15963
rect 14289 15929 14323 15963
rect 14749 15929 14783 15963
rect 17601 15929 17635 15963
rect 18328 15929 18362 15963
rect 20729 15929 20763 15963
rect 22385 15929 22419 15963
rect 4721 15861 4755 15895
rect 5089 15861 5123 15895
rect 6561 15861 6595 15895
rect 8217 15861 8251 15895
rect 8769 15861 8803 15895
rect 11805 15861 11839 15895
rect 12265 15861 12299 15895
rect 13829 15861 13863 15895
rect 14381 15861 14415 15895
rect 15117 15861 15151 15895
rect 15675 15861 15709 15895
rect 17141 15861 17175 15895
rect 19533 15861 19567 15895
rect 19901 15861 19935 15895
rect 19993 15861 20027 15895
rect 20361 15861 20395 15895
rect 20821 15861 20855 15895
rect 21557 15861 21591 15895
rect 22017 15861 22051 15895
rect 23029 15861 23063 15895
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 9965 15657 9999 15691
rect 12173 15657 12207 15691
rect 12731 15657 12765 15691
rect 14197 15657 14231 15691
rect 14657 15657 14691 15691
rect 18705 15657 18739 15691
rect 20361 15657 20395 15691
rect 20637 15657 20671 15691
rect 23029 15657 23063 15691
rect 7113 15589 7147 15623
rect 7297 15589 7331 15623
rect 7840 15589 7874 15623
rect 10425 15589 10459 15623
rect 15568 15589 15602 15623
rect 17592 15589 17626 15623
rect 21640 15589 21674 15623
rect 1593 15521 1627 15555
rect 1860 15521 1894 15555
rect 3433 15521 3467 15555
rect 4344 15521 4378 15555
rect 5549 15521 5583 15555
rect 5816 15521 5850 15555
rect 7481 15521 7515 15555
rect 9505 15521 9539 15555
rect 10333 15521 10367 15555
rect 11060 15521 11094 15555
rect 13001 15521 13035 15555
rect 14565 15521 14599 15555
rect 15301 15521 15335 15555
rect 17233 15521 17267 15555
rect 18981 15521 19015 15555
rect 19248 15521 19282 15555
rect 20453 15521 20487 15555
rect 22845 15521 22879 15555
rect 3525 15453 3559 15487
rect 3709 15453 3743 15487
rect 4077 15453 4111 15487
rect 7573 15453 7607 15487
rect 10517 15453 10551 15487
rect 10793 15453 10827 15487
rect 12265 15453 12299 15487
rect 12771 15453 12805 15487
rect 14749 15453 14783 15487
rect 16773 15453 16807 15487
rect 17325 15453 17359 15487
rect 21373 15453 21407 15487
rect 8953 15385 8987 15419
rect 9321 15385 9355 15419
rect 2973 15317 3007 15351
rect 3065 15317 3099 15351
rect 5457 15317 5491 15351
rect 6929 15317 6963 15351
rect 14105 15317 14139 15351
rect 16681 15317 16715 15351
rect 17049 15317 17083 15351
rect 22753 15317 22787 15351
rect 6377 15113 6411 15147
rect 6469 15113 6503 15147
rect 7665 15113 7699 15147
rect 8677 15113 8711 15147
rect 8861 15113 8895 15147
rect 9321 15113 9355 15147
rect 11529 15113 11563 15147
rect 12817 15113 12851 15147
rect 14565 15113 14599 15147
rect 15669 15113 15703 15147
rect 17785 15113 17819 15147
rect 20085 15113 20119 15147
rect 20177 15113 20211 15147
rect 23029 15113 23063 15147
rect 4905 15045 4939 15079
rect 6837 15045 6871 15079
rect 11713 15045 11747 15079
rect 17509 15045 17543 15079
rect 7389 14977 7423 15011
rect 8125 14977 8159 15011
rect 8217 14977 8251 15011
rect 9965 14977 9999 15011
rect 15301 14977 15335 15011
rect 16313 14977 16347 15011
rect 17049 14977 17083 15011
rect 18705 14977 18739 15011
rect 20729 14977 20763 15011
rect 2053 14909 2087 14943
rect 3525 14909 3559 14943
rect 4997 14909 5031 14943
rect 5264 14909 5298 14943
rect 6653 14909 6687 14943
rect 8033 14909 8067 14943
rect 8493 14909 8527 14943
rect 9045 14909 9079 14943
rect 10149 14909 10183 14943
rect 11805 14909 11839 14943
rect 12173 14909 12207 14943
rect 12449 14909 12483 14943
rect 13001 14909 13035 14943
rect 13185 14909 13219 14943
rect 13452 14909 13486 14943
rect 16037 14909 16071 14943
rect 17325 14909 17359 14943
rect 18061 14909 18095 14943
rect 21373 14909 21407 14943
rect 21640 14909 21674 14943
rect 22845 14909 22879 14943
rect 2320 14841 2354 14875
rect 3770 14841 3804 14875
rect 7297 14841 7331 14875
rect 10416 14841 10450 14875
rect 11989 14841 12023 14875
rect 16129 14841 16163 14875
rect 18972 14841 19006 14875
rect 20545 14841 20579 14875
rect 3433 14773 3467 14807
rect 7205 14773 7239 14807
rect 9137 14773 9171 14807
rect 9689 14773 9723 14807
rect 9781 14773 9815 14807
rect 12633 14773 12667 14807
rect 14657 14773 14691 14807
rect 15025 14773 15059 14807
rect 15117 14773 15151 14807
rect 16497 14773 16531 14807
rect 16865 14773 16899 14807
rect 16957 14773 16991 14807
rect 18245 14773 18279 14807
rect 18521 14773 18555 14807
rect 20637 14773 20671 14807
rect 21097 14773 21131 14807
rect 22753 14773 22787 14807
rect 3157 14569 3191 14603
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 4905 14569 4939 14603
rect 5273 14569 5307 14603
rect 5733 14569 5767 14603
rect 6193 14569 6227 14603
rect 9413 14569 9447 14603
rect 11069 14569 11103 14603
rect 13001 14569 13035 14603
rect 15301 14569 15335 14603
rect 15669 14569 15703 14603
rect 19809 14569 19843 14603
rect 20269 14569 20303 14603
rect 2044 14501 2078 14535
rect 4537 14501 4571 14535
rect 5365 14501 5399 14535
rect 6101 14501 6135 14535
rect 7564 14501 7598 14535
rect 9956 14501 9990 14535
rect 13636 14501 13670 14535
rect 1777 14433 1811 14467
rect 3525 14433 3559 14467
rect 7297 14433 7331 14467
rect 8861 14433 8895 14467
rect 9229 14433 9263 14467
rect 11345 14433 11379 14467
rect 11612 14433 11646 14467
rect 12817 14433 12851 14467
rect 13185 14433 13219 14467
rect 14841 14433 14875 14467
rect 16313 14433 16347 14467
rect 16580 14433 16614 14467
rect 17785 14433 17819 14467
rect 18337 14433 18371 14467
rect 18429 14433 18463 14467
rect 18696 14433 18730 14467
rect 20085 14433 20119 14467
rect 20913 14433 20947 14467
rect 21916 14433 21950 14467
rect 4721 14365 4755 14399
rect 5549 14365 5583 14399
rect 6377 14365 6411 14399
rect 9689 14365 9723 14399
rect 11161 14365 11195 14399
rect 13369 14365 13403 14399
rect 15761 14365 15795 14399
rect 15853 14365 15887 14399
rect 21649 14365 21683 14399
rect 3709 14297 3743 14331
rect 18153 14297 18187 14331
rect 8677 14229 8711 14263
rect 9045 14229 9079 14263
rect 12725 14229 12759 14263
rect 14749 14229 14783 14263
rect 15025 14229 15059 14263
rect 17693 14229 17727 14263
rect 17969 14229 18003 14263
rect 19901 14229 19935 14263
rect 20361 14229 20395 14263
rect 21097 14229 21131 14263
rect 23029 14229 23063 14263
rect 2973 14025 3007 14059
rect 4813 14025 4847 14059
rect 7021 14025 7055 14059
rect 10517 14025 10551 14059
rect 13461 14025 13495 14059
rect 15117 14025 15151 14059
rect 19441 14025 19475 14059
rect 21833 14025 21867 14059
rect 2881 13957 2915 13991
rect 3801 13957 3835 13991
rect 5089 13957 5123 13991
rect 8861 13957 8895 13991
rect 11345 13957 11379 13991
rect 17693 13957 17727 13991
rect 19901 13957 19935 13991
rect 21925 13957 21959 13991
rect 1501 13889 1535 13923
rect 3433 13889 3467 13923
rect 3617 13889 3651 13923
rect 4445 13889 4479 13923
rect 5733 13889 5767 13923
rect 6561 13889 6595 13923
rect 9413 13889 9447 13923
rect 10241 13889 10275 13923
rect 11069 13889 11103 13923
rect 11805 13889 11839 13923
rect 11897 13889 11931 13923
rect 13001 13889 13035 13923
rect 20499 13889 20533 13923
rect 22385 13889 22419 13923
rect 22569 13889 22603 13923
rect 4629 13821 4663 13855
rect 6837 13821 6871 13855
rect 7389 13821 7423 13855
rect 7656 13821 7690 13855
rect 9321 13821 9355 13855
rect 10149 13821 10183 13855
rect 10977 13821 11011 13855
rect 12817 13821 12851 13855
rect 13277 13821 13311 13855
rect 13829 13821 13863 13855
rect 15669 13821 15703 13855
rect 15925 13821 15959 13855
rect 17141 13821 17175 13855
rect 17509 13821 17543 13855
rect 18061 13821 18095 13855
rect 18328 13821 18362 13855
rect 19533 13821 19567 13855
rect 19993 13821 20027 13855
rect 20729 13821 20763 13855
rect 22293 13821 22327 13855
rect 1768 13753 1802 13787
rect 3341 13753 3375 13787
rect 4261 13753 4295 13787
rect 5457 13753 5491 13787
rect 6285 13753 6319 13787
rect 9229 13753 9263 13787
rect 11713 13753 11747 13787
rect 12909 13753 12943 13787
rect 19717 13753 19751 13787
rect 4169 13685 4203 13719
rect 5549 13685 5583 13719
rect 5917 13685 5951 13719
rect 6377 13685 6411 13719
rect 8769 13685 8803 13719
rect 9689 13685 9723 13719
rect 10057 13685 10091 13719
rect 10885 13685 10919 13719
rect 12449 13685 12483 13719
rect 17049 13685 17083 13719
rect 17325 13685 17359 13719
rect 20459 13685 20493 13719
rect 22753 13685 22787 13719
rect 2881 13481 2915 13515
rect 4077 13481 4111 13515
rect 6469 13481 6503 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 12357 13481 12391 13515
rect 14565 13481 14599 13515
rect 16681 13481 16715 13515
rect 19809 13481 19843 13515
rect 20361 13481 20395 13515
rect 3249 13413 3283 13447
rect 6929 13413 6963 13447
rect 7656 13413 7690 13447
rect 15568 13413 15602 13447
rect 17040 13413 17074 13447
rect 20453 13413 20487 13447
rect 21180 13413 21214 13447
rect 22753 13413 22787 13447
rect 4445 13345 4479 13379
rect 4997 13345 5031 13379
rect 5264 13345 5298 13379
rect 6837 13345 6871 13379
rect 8861 13345 8895 13379
rect 9229 13345 9263 13379
rect 10057 13345 10091 13379
rect 10517 13345 10551 13379
rect 11152 13345 11186 13379
rect 12725 13345 12759 13379
rect 13185 13345 13219 13379
rect 13452 13345 13486 13379
rect 14841 13345 14875 13379
rect 15301 13345 15335 13379
rect 16773 13345 16807 13379
rect 18501 13345 18535 13379
rect 22845 13345 22879 13379
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 4537 13277 4571 13311
rect 4721 13277 4755 13311
rect 7021 13277 7055 13311
rect 7389 13277 7423 13311
rect 10241 13277 10275 13311
rect 10885 13277 10919 13311
rect 12817 13277 12851 13311
rect 12909 13277 12943 13311
rect 18245 13277 18279 13311
rect 20637 13277 20671 13311
rect 20913 13277 20947 13311
rect 22937 13277 22971 13311
rect 9045 13209 9079 13243
rect 12265 13209 12299 13243
rect 6377 13141 6411 13175
rect 8769 13141 8803 13175
rect 9413 13141 9447 13175
rect 10701 13141 10735 13175
rect 15025 13141 15059 13175
rect 18153 13141 18187 13175
rect 19625 13141 19659 13175
rect 19993 13141 20027 13175
rect 22293 13141 22327 13175
rect 22385 13141 22419 13175
rect 3985 12937 4019 12971
rect 6101 12937 6135 12971
rect 9689 12937 9723 12971
rect 11989 12937 12023 12971
rect 12633 12937 12667 12971
rect 14381 12937 14415 12971
rect 15301 12937 15335 12971
rect 16957 12937 16991 12971
rect 17785 12937 17819 12971
rect 19717 12937 19751 12971
rect 22017 12937 22051 12971
rect 4077 12869 4111 12903
rect 8769 12869 8803 12903
rect 12081 12869 12115 12903
rect 16129 12869 16163 12903
rect 4721 12801 4755 12835
rect 9321 12801 9355 12835
rect 10241 12801 10275 12835
rect 13001 12801 13035 12835
rect 15025 12801 15059 12835
rect 15853 12801 15887 12835
rect 16681 12801 16715 12835
rect 17509 12801 17543 12835
rect 20177 12801 20211 12835
rect 20361 12801 20395 12835
rect 22477 12801 22511 12835
rect 22661 12801 22695 12835
rect 2605 12733 2639 12767
rect 4261 12733 4295 12767
rect 4988 12733 5022 12767
rect 6653 12733 6687 12767
rect 7205 12733 7239 12767
rect 7297 12733 7331 12767
rect 7564 12733 7598 12767
rect 9229 12733 9263 12767
rect 10609 12733 10643 12767
rect 12265 12733 12299 12767
rect 12449 12733 12483 12767
rect 14933 12733 14967 12767
rect 15669 12733 15703 12767
rect 16497 12733 16531 12767
rect 17325 12733 17359 12767
rect 18061 12733 18095 12767
rect 18328 12733 18362 12767
rect 20545 12733 20579 12767
rect 20812 12733 20846 12767
rect 22385 12733 22419 12767
rect 2872 12665 2906 12699
rect 9137 12665 9171 12699
rect 10149 12665 10183 12699
rect 10876 12665 10910 12699
rect 13268 12665 13302 12699
rect 14841 12665 14875 12699
rect 17417 12665 17451 12699
rect 22845 12665 22879 12699
rect 6469 12597 6503 12631
rect 7021 12597 7055 12631
rect 8677 12597 8711 12631
rect 10057 12597 10091 12631
rect 14473 12597 14507 12631
rect 15761 12597 15795 12631
rect 16589 12597 16623 12631
rect 19441 12597 19475 12631
rect 20085 12597 20119 12631
rect 21925 12597 21959 12631
rect 3433 12393 3467 12427
rect 5457 12393 5491 12427
rect 6929 12393 6963 12427
rect 9321 12393 9355 12427
rect 9689 12393 9723 12427
rect 11529 12393 11563 12427
rect 14841 12393 14875 12427
rect 15301 12393 15335 12427
rect 16773 12393 16807 12427
rect 17233 12393 17267 12427
rect 17601 12393 17635 12427
rect 2320 12325 2354 12359
rect 4344 12325 4378 12359
rect 5816 12325 5850 12359
rect 7288 12325 7322 12359
rect 13369 12325 13403 12359
rect 17693 12325 17727 12359
rect 20453 12325 20487 12359
rect 21434 12325 21468 12359
rect 4077 12257 4111 12291
rect 5549 12257 5583 12291
rect 8861 12257 8895 12291
rect 9505 12257 9539 12291
rect 10149 12257 10183 12291
rect 10416 12257 10450 12291
rect 11621 12257 11655 12291
rect 13728 12257 13762 12291
rect 15117 12257 15151 12291
rect 15485 12257 15519 12291
rect 15945 12257 15979 12291
rect 18613 12257 18647 12291
rect 19441 12257 19475 12291
rect 20361 12257 20395 12291
rect 2053 12189 2087 12223
rect 7021 12189 7055 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 13461 12189 13495 12223
rect 16037 12189 16071 12223
rect 16129 12189 16163 12223
rect 16865 12189 16899 12223
rect 17049 12189 17083 12223
rect 17785 12189 17819 12223
rect 18705 12189 18739 12223
rect 18797 12189 18831 12223
rect 19533 12189 19567 12223
rect 19625 12189 19659 12223
rect 20545 12189 20579 12223
rect 21189 12189 21223 12223
rect 8401 12121 8435 12155
rect 8493 12121 8527 12155
rect 14933 12121 14967 12155
rect 15577 12053 15611 12087
rect 16405 12053 16439 12087
rect 18245 12053 18279 12087
rect 19073 12053 19107 12087
rect 19993 12053 20027 12087
rect 22569 12053 22603 12087
rect 4537 11849 4571 11883
rect 8401 11849 8435 11883
rect 10241 11849 10275 11883
rect 11805 11849 11839 11883
rect 12633 11849 12667 11883
rect 14289 11849 14323 11883
rect 15485 11849 15519 11883
rect 15669 11849 15703 11883
rect 16497 11849 16531 11883
rect 17785 11849 17819 11883
rect 22109 11849 22143 11883
rect 22017 11781 22051 11815
rect 3157 11713 3191 11747
rect 10425 11713 10459 11747
rect 15025 11713 15059 11747
rect 16221 11713 16255 11747
rect 17049 11713 17083 11747
rect 20640 11713 20674 11747
rect 22661 11713 22695 11747
rect 22937 11713 22971 11747
rect 3424 11645 3458 11679
rect 7021 11645 7055 11679
rect 8585 11645 8619 11679
rect 10057 11645 10091 11679
rect 12817 11645 12851 11679
rect 12909 11645 12943 11679
rect 14749 11645 14783 11679
rect 15301 11645 15335 11679
rect 17601 11645 17635 11679
rect 18061 11645 18095 11679
rect 18328 11645 18362 11679
rect 19533 11645 19567 11679
rect 20177 11645 20211 11679
rect 20500 11645 20534 11679
rect 20913 11645 20947 11679
rect 22569 11645 22603 11679
rect 7288 11577 7322 11611
rect 8852 11577 8886 11611
rect 10692 11577 10726 11611
rect 13176 11577 13210 11611
rect 14841 11577 14875 11611
rect 16037 11577 16071 11611
rect 19993 11577 20027 11611
rect 22477 11577 22511 11611
rect 9965 11509 9999 11543
rect 14381 11509 14415 11543
rect 16129 11509 16163 11543
rect 16865 11509 16899 11543
rect 16957 11509 16991 11543
rect 19441 11509 19475 11543
rect 19717 11509 19751 11543
rect 2789 11305 2823 11339
rect 8217 11305 8251 11339
rect 11345 11305 11379 11339
rect 11713 11305 11747 11339
rect 11805 11305 11839 11339
rect 16773 11305 16807 11339
rect 20913 11305 20947 11339
rect 1654 11237 1688 11271
rect 7104 11237 7138 11271
rect 17408 11237 17442 11271
rect 19064 11237 19098 11271
rect 20269 11237 20303 11271
rect 21373 11237 21407 11271
rect 22008 11237 22042 11271
rect 6837 11169 6871 11203
rect 8677 11169 8711 11203
rect 9321 11169 9355 11203
rect 9873 11169 9907 11203
rect 10140 11169 10174 11203
rect 12817 11169 12851 11203
rect 13176 11169 13210 11203
rect 14749 11169 14783 11203
rect 15393 11169 15427 11203
rect 15660 11169 15694 11203
rect 17141 11169 17175 11203
rect 18797 11169 18831 11203
rect 21281 11169 21315 11203
rect 21741 11169 21775 11203
rect 1409 11101 1443 11135
rect 8769 11101 8803 11135
rect 8861 11101 8895 11135
rect 11897 11101 11931 11135
rect 12909 11101 12943 11135
rect 14841 11101 14875 11135
rect 15025 11101 15059 11135
rect 21557 11101 21591 11135
rect 8309 11033 8343 11067
rect 9137 11033 9171 11067
rect 12633 11033 12667 11067
rect 14289 11033 14323 11067
rect 18521 11033 18555 11067
rect 18705 11033 18739 11067
rect 23121 11033 23155 11067
rect 11253 10965 11287 10999
rect 14381 10965 14415 10999
rect 20177 10965 20211 10999
rect 8677 10761 8711 10795
rect 10701 10761 10735 10795
rect 12173 10761 12207 10795
rect 14105 10761 14139 10795
rect 14197 10761 14231 10795
rect 16405 10761 16439 10795
rect 18245 10761 18279 10795
rect 21281 10761 21315 10795
rect 22753 10761 22787 10795
rect 7297 10625 7331 10659
rect 14657 10625 14691 10659
rect 14841 10625 14875 10659
rect 19073 10625 19107 10659
rect 19441 10625 19475 10659
rect 19947 10625 19981 10659
rect 7564 10557 7598 10591
rect 9321 10557 9355 10591
rect 9588 10557 9622 10591
rect 10793 10557 10827 10591
rect 11060 10557 11094 10591
rect 12725 10557 12759 10591
rect 14565 10557 14599 10591
rect 15025 10557 15059 10591
rect 16497 10557 16531 10591
rect 18061 10557 18095 10591
rect 18981 10557 19015 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 12992 10489 13026 10523
rect 15292 10489 15326 10523
rect 16764 10489 16798 10523
rect 18889 10489 18923 10523
rect 21640 10489 21674 10523
rect 1409 10421 1443 10455
rect 17877 10421 17911 10455
rect 18521 10421 18555 10455
rect 19907 10421 19941 10455
rect 22845 10421 22879 10455
rect 9321 10217 9355 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 10517 10217 10551 10251
rect 10885 10217 10919 10251
rect 14381 10217 14415 10251
rect 19349 10217 19383 10251
rect 19993 10217 20027 10251
rect 22293 10217 22327 10251
rect 22753 10217 22787 10251
rect 8208 10149 8242 10183
rect 10149 10149 10183 10183
rect 10977 10149 11011 10183
rect 13176 10149 13210 10183
rect 14749 10149 14783 10183
rect 17233 10149 17267 10183
rect 7941 10081 7975 10115
rect 12449 10081 12483 10115
rect 12541 10081 12575 10115
rect 14841 10081 14875 10115
rect 15568 10081 15602 10115
rect 17509 10081 17543 10115
rect 19901 10081 19935 10115
rect 20913 10081 20947 10115
rect 21180 10081 21214 10115
rect 22845 10081 22879 10115
rect 10241 10013 10275 10047
rect 11069 10013 11103 10047
rect 12909 10013 12943 10047
rect 15025 10013 15059 10047
rect 15301 10013 15335 10047
rect 17141 10013 17175 10047
rect 17832 10013 17866 10047
rect 17972 10013 18006 10047
rect 18245 10013 18279 10047
rect 20177 10013 20211 10047
rect 20545 10013 20579 10047
rect 22937 10013 22971 10047
rect 14289 9945 14323 9979
rect 16681 9945 16715 9979
rect 12725 9877 12759 9911
rect 19533 9877 19567 9911
rect 22385 9877 22419 9911
rect 21189 9673 21223 9707
rect 23581 9673 23615 9707
rect 9689 9605 9723 9639
rect 16313 9605 16347 9639
rect 19441 9605 19475 9639
rect 21281 9605 21315 9639
rect 22937 9605 22971 9639
rect 12081 9537 12115 9571
rect 16957 9537 16991 9571
rect 17693 9537 17727 9571
rect 21833 9537 21867 9571
rect 22753 9537 22787 9571
rect 23581 9537 23615 9571
rect 9873 9469 9907 9503
rect 12449 9469 12483 9503
rect 14197 9469 14231 9503
rect 14464 9469 14498 9503
rect 15853 9469 15887 9503
rect 16681 9469 16715 9503
rect 18061 9469 18095 9503
rect 18328 9469 18362 9503
rect 19717 9469 19751 9503
rect 19809 9469 19843 9503
rect 21649 9469 21683 9503
rect 22293 9469 22327 9503
rect 11897 9401 11931 9435
rect 12716 9401 12750 9435
rect 16773 9401 16807 9435
rect 20076 9401 20110 9435
rect 21741 9401 21775 9435
rect 11529 9333 11563 9367
rect 11989 9333 12023 9367
rect 13829 9333 13863 9367
rect 15577 9333 15611 9367
rect 15669 9333 15703 9367
rect 17141 9333 17175 9367
rect 17509 9333 17543 9367
rect 17601 9333 17635 9367
rect 19533 9333 19567 9367
rect 22477 9333 22511 9367
rect 23029 9333 23063 9367
rect 23581 9333 23615 9367
rect 14657 9129 14691 9163
rect 21557 9129 21591 9163
rect 13544 9061 13578 9095
rect 17316 9061 17350 9095
rect 9689 8993 9723 9027
rect 9956 8993 9990 9027
rect 11437 8993 11471 9027
rect 11805 8993 11839 9027
rect 12072 8993 12106 9027
rect 13277 8993 13311 9027
rect 14933 8993 14967 9027
rect 15301 8993 15335 9027
rect 15557 8993 15591 9027
rect 16957 8993 16991 9027
rect 18788 8993 18822 9027
rect 20361 8993 20395 9027
rect 21649 8993 21683 9027
rect 21916 8993 21950 9027
rect 17049 8925 17083 8959
rect 18521 8925 18555 8959
rect 20453 8925 20487 8959
rect 20545 8925 20579 8959
rect 19993 8857 20027 8891
rect 11069 8789 11103 8823
rect 11621 8789 11655 8823
rect 13185 8789 13219 8823
rect 14749 8789 14783 8823
rect 15117 8789 15151 8823
rect 16681 8789 16715 8823
rect 16773 8789 16807 8823
rect 18429 8789 18463 8823
rect 19901 8789 19935 8823
rect 21005 8789 21039 8823
rect 23029 8789 23063 8823
rect 10609 8585 10643 8619
rect 11529 8585 11563 8619
rect 13829 8585 13863 8619
rect 13921 8585 13955 8619
rect 17141 8585 17175 8619
rect 19901 8585 19935 8619
rect 16957 8517 16991 8551
rect 21925 8517 21959 8551
rect 2053 8449 2087 8483
rect 9229 8449 9263 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 12173 8449 12207 8483
rect 14565 8449 14599 8483
rect 15212 8449 15246 8483
rect 16681 8449 16715 8483
rect 17601 8449 17635 8483
rect 17785 8449 17819 8483
rect 18061 8449 18095 8483
rect 18521 8449 18555 8483
rect 19993 8449 20027 8483
rect 20499 8449 20533 8483
rect 22477 8449 22511 8483
rect 1777 8381 1811 8415
rect 2421 8381 2455 8415
rect 9496 8381 9530 8415
rect 11069 8381 11103 8415
rect 11897 8381 11931 8415
rect 12449 8381 12483 8415
rect 12716 8381 12750 8415
rect 14757 8381 14791 8415
rect 15485 8381 15519 8415
rect 18788 8381 18822 8415
rect 20729 8381 20763 8415
rect 22753 8381 22787 8415
rect 14289 8313 14323 8347
rect 17509 8313 17543 8347
rect 22293 8313 22327 8347
rect 10701 8245 10735 8279
rect 11989 8245 12023 8279
rect 14381 8245 14415 8279
rect 15215 8245 15249 8279
rect 16589 8245 16623 8279
rect 18337 8245 18371 8279
rect 20459 8245 20493 8279
rect 21833 8245 21867 8279
rect 22385 8245 22419 8279
rect 22937 8245 22971 8279
rect 9321 8041 9355 8075
rect 12265 8041 12299 8075
rect 12633 8041 12667 8075
rect 14381 8041 14415 8075
rect 15485 8041 15519 8075
rect 16503 8041 16537 8075
rect 17877 8041 17911 8075
rect 20453 8041 20487 8075
rect 22569 8041 22603 8075
rect 8585 7973 8619 8007
rect 9956 7973 9990 8007
rect 13461 7973 13495 8007
rect 14749 7973 14783 8007
rect 18245 7973 18279 8007
rect 22937 7973 22971 8007
rect 7757 7905 7791 7939
rect 8861 7905 8895 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 11529 7905 11563 7939
rect 12725 7905 12759 7939
rect 13553 7905 13587 7939
rect 14013 7905 14047 7939
rect 15301 7905 15335 7939
rect 16037 7905 16071 7939
rect 16773 7905 16807 7939
rect 17969 7905 18003 7939
rect 18521 7905 18555 7939
rect 18844 7905 18878 7939
rect 21456 7905 21490 7939
rect 22661 7905 22695 7939
rect 11621 7837 11655 7871
rect 11805 7837 11839 7871
rect 12817 7837 12851 7871
rect 13737 7837 13771 7871
rect 14841 7837 14875 7871
rect 15025 7837 15059 7871
rect 15669 7837 15703 7871
rect 16500 7837 16534 7871
rect 19027 7837 19061 7871
rect 19257 7837 19291 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 20361 7769 20395 7803
rect 11069 7701 11103 7735
rect 11161 7701 11195 7735
rect 13093 7701 13127 7735
rect 14197 7701 14231 7735
rect 10701 7497 10735 7531
rect 11805 7497 11839 7531
rect 12449 7497 12483 7531
rect 14105 7497 14139 7531
rect 17693 7497 17727 7531
rect 19441 7497 19475 7531
rect 21833 7497 21867 7531
rect 10793 7429 10827 7463
rect 12265 7429 12299 7463
rect 19625 7429 19659 7463
rect 9321 7361 9355 7395
rect 11253 7361 11287 7395
rect 11437 7361 11471 7395
rect 13093 7361 13127 7395
rect 14841 7361 14875 7395
rect 17417 7361 17451 7395
rect 18061 7361 18095 7395
rect 20085 7361 20119 7395
rect 20269 7361 20303 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 9588 7293 9622 7327
rect 11161 7293 11195 7327
rect 11621 7293 11655 7327
rect 13277 7293 13311 7327
rect 13737 7293 13771 7327
rect 14657 7293 14691 7327
rect 15025 7293 15059 7327
rect 15393 7293 15427 7327
rect 17325 7293 17359 7327
rect 17877 7293 17911 7327
rect 20453 7293 20487 7327
rect 22753 7293 22787 7327
rect 12817 7225 12851 7259
rect 13921 7225 13955 7259
rect 15660 7225 15694 7259
rect 17233 7225 17267 7259
rect 18306 7225 18340 7259
rect 20720 7225 20754 7259
rect 12909 7157 12943 7191
rect 13461 7157 13495 7191
rect 14197 7157 14231 7191
rect 14565 7157 14599 7191
rect 15209 7157 15243 7191
rect 16773 7157 16807 7191
rect 16865 7157 16899 7191
rect 19993 7157 20027 7191
rect 21925 7157 21959 7191
rect 22293 7157 22327 7191
rect 22937 7157 22971 7191
rect 13185 6953 13219 6987
rect 13553 6953 13587 6987
rect 14749 6953 14783 6987
rect 18153 6953 18187 6987
rect 18613 6953 18647 6987
rect 19349 6953 19383 6987
rect 22293 6953 22327 6987
rect 9956 6885 9990 6919
rect 9689 6817 9723 6851
rect 11529 6817 11563 6851
rect 11989 6817 12023 6851
rect 12725 6817 12759 6851
rect 14013 6817 14047 6851
rect 15568 6817 15602 6851
rect 16773 6817 16807 6851
rect 17040 6817 17074 6851
rect 20177 6817 20211 6851
rect 20913 6817 20947 6851
rect 21281 6817 21315 6851
rect 21649 6817 21683 6851
rect 22385 6817 22419 6851
rect 22753 6817 22787 6851
rect 11621 6749 11655 6783
rect 11805 6749 11839 6783
rect 12817 6749 12851 6783
rect 13001 6749 13035 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 14841 6749 14875 6783
rect 15025 6749 15059 6783
rect 15301 6749 15335 6783
rect 18245 6749 18279 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 22477 6749 22511 6783
rect 12357 6681 12391 6715
rect 14197 6681 14231 6715
rect 16681 6681 16715 6715
rect 18981 6681 19015 6715
rect 11069 6613 11103 6647
rect 11161 6613 11195 6647
rect 12173 6613 12207 6647
rect 14381 6613 14415 6647
rect 19809 6613 19843 6647
rect 20729 6613 20763 6647
rect 21097 6613 21131 6647
rect 21465 6613 21499 6647
rect 21925 6613 21959 6647
rect 22937 6613 22971 6647
rect 10333 6409 10367 6443
rect 15577 6409 15611 6443
rect 17049 6409 17083 6443
rect 23121 6409 23155 6443
rect 18521 6341 18555 6375
rect 18705 6341 18739 6375
rect 20913 6341 20947 6375
rect 8953 6273 8987 6307
rect 10425 6273 10459 6307
rect 17601 6273 17635 6307
rect 17785 6273 17819 6307
rect 19165 6273 19199 6307
rect 19349 6273 19383 6307
rect 21557 6273 21591 6307
rect 22477 6273 22511 6307
rect 9220 6205 9254 6239
rect 12725 6205 12759 6239
rect 14197 6205 14231 6239
rect 15669 6205 15703 6239
rect 15925 6205 15959 6239
rect 17509 6205 17543 6239
rect 18337 6205 18371 6239
rect 19540 6205 19574 6239
rect 19800 6205 19834 6239
rect 21373 6205 21407 6239
rect 21833 6205 21867 6239
rect 22201 6205 22235 6239
rect 22753 6205 22787 6239
rect 10692 6137 10726 6171
rect 12992 6137 13026 6171
rect 14442 6137 14476 6171
rect 18061 6137 18095 6171
rect 19073 6137 19107 6171
rect 21465 6137 21499 6171
rect 22937 6137 22971 6171
rect 11805 6069 11839 6103
rect 14105 6069 14139 6103
rect 17141 6069 17175 6103
rect 21005 6069 21039 6103
rect 22017 6069 22051 6103
rect 11345 5865 11379 5899
rect 12817 5865 12851 5899
rect 14289 5865 14323 5899
rect 14381 5865 14415 5899
rect 14749 5865 14783 5899
rect 15301 5865 15335 5899
rect 15669 5865 15703 5899
rect 20361 5865 20395 5899
rect 20637 5865 20671 5899
rect 20913 5865 20947 5899
rect 21281 5865 21315 5899
rect 23121 5865 23155 5899
rect 10232 5797 10266 5831
rect 11704 5797 11738 5831
rect 13154 5797 13188 5831
rect 14841 5797 14875 5831
rect 15761 5797 15795 5831
rect 19248 5797 19282 5831
rect 9965 5729 9999 5763
rect 11437 5729 11471 5763
rect 12909 5729 12943 5763
rect 16672 5729 16706 5763
rect 18245 5729 18279 5763
rect 18981 5729 19015 5763
rect 20453 5729 20487 5763
rect 22008 5729 22042 5763
rect 14933 5661 14967 5695
rect 15945 5661 15979 5695
rect 16405 5661 16439 5695
rect 18337 5661 18371 5695
rect 18521 5661 18555 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 21741 5661 21775 5695
rect 17785 5525 17819 5559
rect 17877 5525 17911 5559
rect 13829 5321 13863 5355
rect 14197 5321 14231 5355
rect 17325 5321 17359 5355
rect 18061 5321 18095 5355
rect 18889 5321 18923 5355
rect 20729 5321 20763 5355
rect 22937 5321 22971 5355
rect 19717 5253 19751 5287
rect 23029 5253 23063 5287
rect 11437 5185 11471 5219
rect 11621 5185 11655 5219
rect 18521 5185 18555 5219
rect 18705 5185 18739 5219
rect 19533 5185 19567 5219
rect 20269 5185 20303 5219
rect 21281 5185 21315 5219
rect 12449 5117 12483 5151
rect 14381 5117 14415 5151
rect 15945 5117 15979 5151
rect 17601 5117 17635 5151
rect 19257 5117 19291 5151
rect 21557 5117 21591 5151
rect 11345 5049 11379 5083
rect 12716 5049 12750 5083
rect 16212 5049 16246 5083
rect 19349 5049 19383 5083
rect 21097 5049 21131 5083
rect 21824 5049 21858 5083
rect 10977 4981 11011 5015
rect 17785 4981 17819 5015
rect 18429 4981 18463 5015
rect 20085 4981 20119 5015
rect 20177 4981 20211 5015
rect 21189 4981 21223 5015
rect 11253 4777 11287 4811
rect 17877 4777 17911 4811
rect 19533 4777 19567 4811
rect 20545 4777 20579 4811
rect 21465 4777 21499 4811
rect 22937 4777 22971 4811
rect 11161 4709 11195 4743
rect 16672 4709 16706 4743
rect 23029 4709 23063 4743
rect 16405 4641 16439 4675
rect 18245 4641 18279 4675
rect 19073 4641 19107 4675
rect 19901 4641 19935 4675
rect 20361 4641 20395 4675
rect 20913 4641 20947 4675
rect 21557 4641 21591 4675
rect 21824 4641 21858 4675
rect 11437 4573 11471 4607
rect 18337 4573 18371 4607
rect 18521 4573 18555 4607
rect 19165 4573 19199 4607
rect 19257 4573 19291 4607
rect 19993 4573 20027 4607
rect 20085 4573 20119 4607
rect 10793 4505 10827 4539
rect 18705 4505 18739 4539
rect 17785 4437 17819 4471
rect 21097 4437 21131 4471
rect 19625 4233 19659 4267
rect 22845 4233 22879 4267
rect 21465 4097 21499 4131
rect 23029 4097 23063 4131
rect 16313 4029 16347 4063
rect 16580 4029 16614 4063
rect 18245 4029 18279 4063
rect 19717 4029 19751 4063
rect 19984 4029 20018 4063
rect 18512 3961 18546 3995
rect 21732 3961 21766 3995
rect 17693 3893 17727 3927
rect 21097 3893 21131 3927
rect 3525 3689 3559 3723
rect 19441 3689 19475 3723
rect 19809 3689 19843 3723
rect 20453 3689 20487 3723
rect 22293 3689 22327 3723
rect 22845 3689 22879 3723
rect 3157 3621 3191 3655
rect 16764 3621 16798 3655
rect 2329 3553 2363 3587
rect 18225 3553 18259 3587
rect 20269 3553 20303 3587
rect 20913 3553 20947 3587
rect 21169 3553 21203 3587
rect 22753 3553 22787 3587
rect 16497 3485 16531 3519
rect 17969 3485 18003 3519
rect 19901 3485 19935 3519
rect 20085 3485 20119 3519
rect 22937 3485 22971 3519
rect 19349 3417 19383 3451
rect 22385 3417 22419 3451
rect 17877 3349 17911 3383
rect 2329 3145 2363 3179
rect 2973 3145 3007 3179
rect 17877 3145 17911 3179
rect 18061 3145 18095 3179
rect 22201 3145 22235 3179
rect 22293 3145 22327 3179
rect 2697 3077 2731 3111
rect 1961 3009 1995 3043
rect 18705 3009 18739 3043
rect 22937 3009 22971 3043
rect 1777 2941 1811 2975
rect 2501 2941 2535 2975
rect 6101 2941 6135 2975
rect 16497 2941 16531 2975
rect 18429 2941 18463 2975
rect 19349 2941 19383 2975
rect 19616 2941 19650 2975
rect 20821 2941 20855 2975
rect 22661 2941 22695 2975
rect 22753 2941 22787 2975
rect 16764 2873 16798 2907
rect 18521 2873 18555 2907
rect 21066 2873 21100 2907
rect 20729 2805 20763 2839
rect 19717 2601 19751 2635
rect 20269 2601 20303 2635
rect 20729 2601 20763 2635
rect 22569 2601 22603 2635
rect 18604 2533 18638 2567
rect 20637 2533 20671 2567
rect 21456 2533 21490 2567
rect 18337 2465 18371 2499
rect 21189 2465 21223 2499
rect 22661 2465 22695 2499
rect 20821 2397 20855 2431
rect 22845 2397 22879 2431
<< metal1 >>
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 6914 22488 6920 22500
rect 5592 22460 6920 22488
rect 5592 22448 5598 22460
rect 6914 22448 6920 22460
rect 6972 22488 6978 22500
rect 8662 22488 8668 22500
rect 6972 22460 8668 22488
rect 6972 22448 6978 22460
rect 8662 22448 8668 22460
rect 8720 22448 8726 22500
rect 5442 22380 5448 22432
rect 5500 22420 5506 22432
rect 6638 22420 6644 22432
rect 5500 22392 6644 22420
rect 5500 22380 5506 22392
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14826 22420 14832 22432
rect 13872 22392 14832 22420
rect 13872 22380 13878 22392
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 1104 22330 23460 22352
rect 1104 22278 8446 22330
rect 8498 22278 8510 22330
rect 8562 22278 8574 22330
rect 8626 22278 8638 22330
rect 8690 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 23460 22330
rect 1104 22256 23460 22278
rect 5092 22188 7052 22216
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4709 22083 4767 22089
rect 4709 22080 4721 22083
rect 4387 22052 4721 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4709 22049 4721 22052
rect 4755 22080 4767 22083
rect 5092 22080 5120 22188
rect 5350 22108 5356 22160
rect 5408 22148 5414 22160
rect 6365 22151 6423 22157
rect 6365 22148 6377 22151
rect 5408 22120 6377 22148
rect 5408 22108 5414 22120
rect 6365 22117 6377 22120
rect 6411 22117 6423 22151
rect 6914 22148 6920 22160
rect 6875 22120 6920 22148
rect 6365 22111 6423 22117
rect 6914 22108 6920 22120
rect 6972 22108 6978 22160
rect 4755 22052 5120 22080
rect 5169 22083 5227 22089
rect 4755 22049 4767 22052
rect 4709 22043 4767 22049
rect 5169 22049 5181 22083
rect 5215 22080 5227 22083
rect 5258 22080 5264 22092
rect 5215 22052 5264 22080
rect 5215 22049 5227 22052
rect 5169 22043 5227 22049
rect 5258 22040 5264 22052
rect 5316 22040 5322 22092
rect 5534 22040 5540 22092
rect 5592 22080 5598 22092
rect 6270 22080 6276 22092
rect 5592 22052 5637 22080
rect 6231 22052 6276 22080
rect 5592 22040 5598 22052
rect 6270 22040 6276 22052
rect 6328 22040 6334 22092
rect 7024 22080 7052 22188
rect 7558 22176 7564 22228
rect 7616 22216 7622 22228
rect 7745 22219 7803 22225
rect 7745 22216 7757 22219
rect 7616 22188 7757 22216
rect 7616 22176 7622 22188
rect 7745 22185 7757 22188
rect 7791 22185 7803 22219
rect 7745 22179 7803 22185
rect 8018 22176 8024 22228
rect 8076 22216 8082 22228
rect 8113 22219 8171 22225
rect 8113 22216 8125 22219
rect 8076 22188 8125 22216
rect 8076 22176 8082 22188
rect 8113 22185 8125 22188
rect 8159 22185 8171 22219
rect 8113 22179 8171 22185
rect 12360 22188 15332 22216
rect 7653 22151 7711 22157
rect 7653 22117 7665 22151
rect 7699 22148 7711 22151
rect 8386 22148 8392 22160
rect 7699 22120 8392 22148
rect 7699 22117 7711 22120
rect 7653 22111 7711 22117
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 10594 22148 10600 22160
rect 9968 22120 10272 22148
rect 10555 22120 10600 22148
rect 7024 22052 7972 22080
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 2685 22015 2743 22021
rect 2685 22012 2697 22015
rect 2464 21984 2697 22012
rect 2464 21972 2470 21984
rect 2685 21981 2697 21984
rect 2731 22012 2743 22015
rect 5902 22012 5908 22024
rect 2731 21984 5908 22012
rect 2731 21981 2743 21984
rect 2685 21975 2743 21981
rect 5902 21972 5908 21984
rect 5960 21972 5966 22024
rect 6454 21972 6460 22024
rect 6512 22012 6518 22024
rect 7834 22012 7840 22024
rect 6512 21984 6557 22012
rect 7795 21984 7840 22012
rect 6512 21972 6518 21984
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 7944 22012 7972 22052
rect 9968 22012 9996 22120
rect 10134 22080 10140 22092
rect 10095 22052 10140 22080
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 10244 22080 10272 22120
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 12360 22080 12388 22188
rect 13078 22108 13084 22160
rect 13136 22148 13142 22160
rect 13357 22151 13415 22157
rect 13357 22148 13369 22151
rect 13136 22120 13369 22148
rect 13136 22108 13142 22120
rect 13357 22117 13369 22120
rect 13403 22117 13415 22151
rect 13357 22111 13415 22117
rect 14182 22108 14188 22160
rect 14240 22148 14246 22160
rect 14461 22151 14519 22157
rect 14461 22148 14473 22151
rect 14240 22120 14473 22148
rect 14240 22108 14246 22120
rect 14461 22117 14473 22120
rect 14507 22117 14519 22151
rect 14461 22111 14519 22117
rect 15304 22092 15332 22188
rect 17773 22151 17831 22157
rect 15764 22120 15976 22148
rect 10244 22052 12388 22080
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22080 12495 22083
rect 12618 22080 12624 22092
rect 12483 22052 12624 22080
rect 12483 22049 12495 22052
rect 12437 22043 12495 22049
rect 12618 22040 12624 22052
rect 12676 22080 12682 22092
rect 13170 22080 13176 22092
rect 12676 22052 13176 22080
rect 12676 22040 12682 22052
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22080 13323 22083
rect 13722 22080 13728 22092
rect 13311 22052 13728 22080
rect 13311 22049 13323 22052
rect 13265 22043 13323 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 14369 22083 14427 22089
rect 14369 22049 14381 22083
rect 14415 22080 14427 22083
rect 14826 22080 14832 22092
rect 14415 22052 14504 22080
rect 14787 22052 14832 22080
rect 14415 22049 14427 22052
rect 14369 22043 14427 22049
rect 14476 22024 14504 22052
rect 14826 22040 14832 22052
rect 14884 22080 14890 22092
rect 15197 22083 15255 22089
rect 15197 22080 15209 22083
rect 14884 22052 15209 22080
rect 14884 22040 14890 22052
rect 15197 22049 15209 22052
rect 15243 22049 15255 22083
rect 15197 22043 15255 22049
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 15473 22083 15531 22089
rect 15473 22049 15485 22083
rect 15519 22080 15531 22083
rect 15764 22080 15792 22120
rect 15519 22052 15792 22080
rect 15841 22083 15899 22089
rect 15519 22049 15531 22052
rect 15473 22043 15531 22049
rect 15841 22049 15853 22083
rect 15887 22049 15899 22083
rect 15948 22080 15976 22120
rect 17773 22117 17785 22151
rect 17819 22148 17831 22151
rect 18046 22148 18052 22160
rect 17819 22120 18052 22148
rect 17819 22117 17831 22120
rect 17773 22111 17831 22117
rect 18046 22108 18052 22120
rect 18104 22108 18110 22160
rect 16209 22083 16267 22089
rect 16209 22080 16221 22083
rect 15948 22052 16221 22080
rect 15841 22043 15899 22049
rect 16209 22049 16221 22052
rect 16255 22049 16267 22083
rect 16209 22043 16267 22049
rect 17865 22083 17923 22089
rect 17865 22049 17877 22083
rect 17911 22080 17923 22083
rect 19426 22080 19432 22092
rect 17911 22052 19432 22080
rect 17911 22049 17923 22052
rect 17865 22043 17923 22049
rect 10226 22012 10232 22024
rect 7944 21984 9996 22012
rect 10187 21984 10232 22012
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10413 22015 10471 22021
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 11054 22012 11060 22024
rect 10459 21984 11060 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 13354 22012 13360 22024
rect 12032 21984 13360 22012
rect 12032 21972 12038 21984
rect 13354 21972 13360 21984
rect 13412 22012 13418 22024
rect 13541 22015 13599 22021
rect 13541 22012 13553 22015
rect 13412 21984 13553 22012
rect 13412 21972 13418 21984
rect 13541 21981 13553 21984
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 4154 21904 4160 21956
rect 4212 21944 4218 21956
rect 4893 21947 4951 21953
rect 4893 21944 4905 21947
rect 4212 21916 4905 21944
rect 4212 21904 4218 21916
rect 4893 21913 4905 21916
rect 4939 21913 4951 21947
rect 4893 21907 4951 21913
rect 5258 21904 5264 21956
rect 5316 21944 5322 21956
rect 5810 21944 5816 21956
rect 5316 21916 5816 21944
rect 5316 21904 5322 21916
rect 5810 21904 5816 21916
rect 5868 21904 5874 21956
rect 12894 21944 12900 21956
rect 12855 21916 12900 21944
rect 12894 21904 12900 21916
rect 12952 21904 12958 21956
rect 13556 21944 13584 21975
rect 14458 21972 14464 22024
rect 14516 21972 14522 22024
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 14660 21944 14688 21975
rect 14918 21972 14924 22024
rect 14976 22012 14982 22024
rect 15488 22012 15516 22043
rect 14976 21984 15516 22012
rect 14976 21972 14982 21984
rect 13556 21916 14688 21944
rect 15194 21904 15200 21956
rect 15252 21944 15258 21956
rect 15856 21944 15884 22043
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 23566 22080 23572 22092
rect 23527 22052 23572 22080
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 17957 22015 18015 22021
rect 17957 22012 17969 22015
rect 17880 21984 17969 22012
rect 17880 21956 17908 21984
rect 17957 21981 17969 21984
rect 18003 21981 18015 22015
rect 17957 21975 18015 21981
rect 15252 21916 15884 21944
rect 15252 21904 15258 21916
rect 17862 21904 17868 21956
rect 17920 21904 17926 21956
rect 24118 21944 24124 21956
rect 17972 21916 24124 21944
rect 2314 21876 2320 21888
rect 2275 21848 2320 21876
rect 2314 21836 2320 21848
rect 2372 21836 2378 21888
rect 4522 21876 4528 21888
rect 4483 21848 4528 21876
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 5353 21879 5411 21885
rect 5353 21845 5365 21879
rect 5399 21876 5411 21879
rect 5534 21876 5540 21888
rect 5399 21848 5540 21876
rect 5399 21845 5411 21848
rect 5353 21839 5411 21845
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 5718 21876 5724 21888
rect 5679 21848 5724 21876
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 5905 21879 5963 21885
rect 5905 21845 5917 21879
rect 5951 21876 5963 21879
rect 7190 21876 7196 21888
rect 5951 21848 7196 21876
rect 5951 21845 5963 21848
rect 5905 21839 5963 21845
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 7285 21879 7343 21885
rect 7285 21845 7297 21879
rect 7331 21876 7343 21879
rect 7650 21876 7656 21888
rect 7331 21848 7656 21876
rect 7331 21845 7343 21848
rect 7285 21839 7343 21845
rect 7650 21836 7656 21848
rect 7708 21836 7714 21888
rect 7834 21836 7840 21888
rect 7892 21876 7898 21888
rect 9769 21879 9827 21885
rect 9769 21876 9781 21879
rect 7892 21848 9781 21876
rect 7892 21836 7898 21848
rect 9769 21845 9781 21848
rect 9815 21876 9827 21879
rect 13814 21876 13820 21888
rect 9815 21848 13820 21876
rect 9815 21845 9827 21848
rect 9769 21839 9827 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 13998 21876 14004 21888
rect 13959 21848 14004 21876
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 14734 21836 14740 21888
rect 14792 21876 14798 21888
rect 14918 21876 14924 21888
rect 14792 21848 14924 21876
rect 14792 21836 14798 21848
rect 14918 21836 14924 21848
rect 14976 21876 14982 21888
rect 15013 21879 15071 21885
rect 15013 21876 15025 21879
rect 14976 21848 15025 21876
rect 14976 21836 14982 21848
rect 15013 21845 15025 21848
rect 15059 21845 15071 21879
rect 15654 21876 15660 21888
rect 15615 21848 15660 21876
rect 15013 21839 15071 21845
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 16025 21879 16083 21885
rect 16025 21845 16037 21879
rect 16071 21876 16083 21879
rect 16298 21876 16304 21888
rect 16071 21848 16304 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 17402 21876 17408 21888
rect 17363 21848 17408 21876
rect 17402 21836 17408 21848
rect 17460 21876 17466 21888
rect 17972 21876 18000 21916
rect 24118 21904 24124 21916
rect 24176 21904 24182 21956
rect 17460 21848 18000 21876
rect 17460 21836 17466 21848
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 18325 21879 18383 21885
rect 18325 21876 18337 21879
rect 18288 21848 18337 21876
rect 18288 21836 18294 21848
rect 18325 21845 18337 21848
rect 18371 21845 18383 21879
rect 18325 21839 18383 21845
rect 1104 21786 23460 21808
rect 1104 21734 4714 21786
rect 4766 21734 4778 21786
rect 4830 21734 4842 21786
rect 4894 21734 4906 21786
rect 4958 21734 12178 21786
rect 12230 21734 12242 21786
rect 12294 21734 12306 21786
rect 12358 21734 12370 21786
rect 12422 21734 19642 21786
rect 19694 21734 19706 21786
rect 19758 21734 19770 21786
rect 19822 21734 19834 21786
rect 19886 21734 23460 21786
rect 1104 21712 23460 21734
rect 290 21632 296 21684
rect 348 21672 354 21684
rect 2041 21675 2099 21681
rect 2041 21672 2053 21675
rect 348 21644 2053 21672
rect 348 21632 354 21644
rect 2041 21641 2053 21644
rect 2087 21641 2099 21675
rect 2041 21635 2099 21641
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 4249 21675 4307 21681
rect 4249 21672 4261 21675
rect 2924 21644 4261 21672
rect 2924 21632 2930 21644
rect 4249 21641 4261 21644
rect 4295 21641 4307 21675
rect 4249 21635 4307 21641
rect 5166 21632 5172 21684
rect 5224 21672 5230 21684
rect 6181 21675 6239 21681
rect 6181 21672 6193 21675
rect 5224 21644 6193 21672
rect 5224 21632 5230 21644
rect 6181 21641 6193 21644
rect 6227 21641 6239 21675
rect 6181 21635 6239 21641
rect 6730 21632 6736 21684
rect 6788 21672 6794 21684
rect 6825 21675 6883 21681
rect 6825 21672 6837 21675
rect 6788 21644 6837 21672
rect 6788 21632 6794 21644
rect 6825 21641 6837 21644
rect 6871 21641 6883 21675
rect 7558 21672 7564 21684
rect 7519 21644 7564 21672
rect 6825 21635 6883 21641
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 11790 21672 11796 21684
rect 7708 21644 11796 21672
rect 7708 21632 7714 21644
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12618 21672 12624 21684
rect 11992 21644 12624 21672
rect 934 21564 940 21616
rect 992 21604 998 21616
rect 2409 21607 2467 21613
rect 2409 21604 2421 21607
rect 992 21576 2421 21604
rect 992 21564 998 21576
rect 2409 21573 2421 21576
rect 2455 21573 2467 21607
rect 7668 21604 7696 21632
rect 2409 21567 2467 21573
rect 5552 21576 7696 21604
rect 2314 21536 2320 21548
rect 1872 21508 2320 21536
rect 1872 21477 1900 21508
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 4525 21539 4583 21545
rect 4525 21505 4537 21539
rect 4571 21536 4583 21539
rect 4571 21508 4660 21536
rect 4571 21505 4583 21508
rect 4525 21499 4583 21505
rect 4632 21480 4660 21508
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 2225 21471 2283 21477
rect 2225 21437 2237 21471
rect 2271 21468 2283 21471
rect 2406 21468 2412 21480
rect 2271 21440 2412 21468
rect 2271 21437 2283 21440
rect 2225 21431 2283 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 2590 21468 2596 21480
rect 2551 21440 2596 21468
rect 2590 21428 2596 21440
rect 2648 21428 2654 21480
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 4111 21440 4568 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 4540 21412 4568 21440
rect 4614 21428 4620 21480
rect 4672 21428 4678 21480
rect 5074 21428 5080 21480
rect 5132 21468 5138 21480
rect 5552 21468 5580 21576
rect 5902 21496 5908 21548
rect 5960 21536 5966 21548
rect 7834 21536 7840 21548
rect 5960 21508 7840 21536
rect 5960 21496 5966 21508
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 8110 21536 8116 21548
rect 8071 21508 8116 21536
rect 8110 21496 8116 21508
rect 8168 21496 8174 21548
rect 8386 21536 8392 21548
rect 8347 21508 8392 21536
rect 8386 21496 8392 21508
rect 8444 21496 8450 21548
rect 5132 21440 5580 21468
rect 5997 21471 6055 21477
rect 5132 21428 5138 21440
rect 5997 21437 6009 21471
rect 6043 21437 6055 21471
rect 5997 21431 6055 21437
rect 6365 21471 6423 21477
rect 6365 21437 6377 21471
rect 6411 21468 6423 21471
rect 6730 21468 6736 21480
rect 6411 21440 6736 21468
rect 6411 21437 6423 21440
rect 6365 21431 6423 21437
rect 2860 21403 2918 21409
rect 2860 21369 2872 21403
rect 2906 21400 2918 21403
rect 4338 21400 4344 21412
rect 2906 21372 4344 21400
rect 2906 21369 2918 21372
rect 2860 21363 2918 21369
rect 4338 21360 4344 21372
rect 4396 21360 4402 21412
rect 4522 21360 4528 21412
rect 4580 21360 4586 21412
rect 4792 21403 4850 21409
rect 4792 21369 4804 21403
rect 4838 21400 4850 21403
rect 5442 21400 5448 21412
rect 4838 21372 5448 21400
rect 4838 21369 4850 21372
rect 4792 21363 4850 21369
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 6012 21400 6040 21431
rect 6730 21428 6736 21440
rect 6788 21428 6794 21480
rect 7009 21471 7067 21477
rect 7009 21437 7021 21471
rect 7055 21468 7067 21471
rect 8018 21468 8024 21480
rect 7055 21440 8024 21468
rect 7055 21437 7067 21440
rect 7009 21431 7067 21437
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 9030 21468 9036 21480
rect 8991 21440 9036 21468
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 10042 21468 10048 21480
rect 9140 21440 10048 21468
rect 7469 21403 7527 21409
rect 7469 21400 7481 21403
rect 6012 21372 7481 21400
rect 7469 21369 7481 21372
rect 7515 21400 7527 21403
rect 9140 21400 9168 21440
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 10502 21468 10508 21480
rect 10463 21440 10508 21468
rect 10502 21428 10508 21440
rect 10560 21428 10566 21480
rect 11992 21477 12020 21644
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 13817 21675 13875 21681
rect 13817 21672 13829 21675
rect 13780 21644 13829 21672
rect 13780 21632 13786 21644
rect 13817 21641 13829 21644
rect 13863 21641 13875 21675
rect 13817 21635 13875 21641
rect 13906 21632 13912 21684
rect 13964 21672 13970 21684
rect 13964 21644 14872 21672
rect 13964 21632 13970 21644
rect 12066 21564 12072 21616
rect 12124 21604 12130 21616
rect 12161 21607 12219 21613
rect 12161 21604 12173 21607
rect 12124 21576 12173 21604
rect 12124 21564 12130 21576
rect 12161 21573 12173 21576
rect 12207 21573 12219 21607
rect 14844 21604 14872 21644
rect 14918 21632 14924 21684
rect 14976 21672 14982 21684
rect 17678 21672 17684 21684
rect 14976 21644 15976 21672
rect 17639 21644 17684 21672
rect 14976 21632 14982 21644
rect 14844 21576 15884 21604
rect 12161 21567 12219 21573
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21437 12035 21471
rect 11977 21431 12035 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21437 12495 21471
rect 13906 21468 13912 21480
rect 13867 21440 13912 21468
rect 12437 21431 12495 21437
rect 7515 21372 9168 21400
rect 9300 21403 9358 21409
rect 7515 21369 7527 21372
rect 7469 21363 7527 21369
rect 9300 21369 9312 21403
rect 9346 21400 9358 21403
rect 9346 21372 10548 21400
rect 9346 21369 9358 21372
rect 9300 21363 9358 21369
rect 3973 21335 4031 21341
rect 3973 21301 3985 21335
rect 4019 21332 4031 21335
rect 4154 21332 4160 21344
rect 4019 21304 4160 21332
rect 4019 21301 4031 21304
rect 3973 21295 4031 21301
rect 4154 21292 4160 21304
rect 4212 21292 4218 21344
rect 5902 21332 5908 21344
rect 5863 21304 5908 21332
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 6546 21332 6552 21344
rect 6507 21304 6552 21332
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7193 21335 7251 21341
rect 7193 21332 7205 21335
rect 6972 21304 7205 21332
rect 6972 21292 6978 21304
rect 7193 21301 7205 21304
rect 7239 21301 7251 21335
rect 7193 21295 7251 21301
rect 7282 21292 7288 21344
rect 7340 21332 7346 21344
rect 7742 21332 7748 21344
rect 7340 21304 7748 21332
rect 7340 21292 7346 21304
rect 7742 21292 7748 21304
rect 7800 21332 7806 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7800 21304 7941 21332
rect 7800 21292 7806 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 7929 21295 7987 21301
rect 8021 21335 8079 21341
rect 8021 21301 8033 21335
rect 8067 21332 8079 21335
rect 8202 21332 8208 21344
rect 8067 21304 8208 21332
rect 8067 21301 8079 21304
rect 8021 21295 8079 21301
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 10042 21332 10048 21344
rect 8352 21304 10048 21332
rect 8352 21292 8358 21304
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 10410 21332 10416 21344
rect 10371 21304 10416 21332
rect 10410 21292 10416 21304
rect 10468 21292 10474 21344
rect 10520 21332 10548 21372
rect 10686 21360 10692 21412
rect 10744 21409 10750 21412
rect 10744 21403 10808 21409
rect 10744 21369 10762 21403
rect 10796 21369 10808 21403
rect 12452 21400 12480 21431
rect 13906 21428 13912 21440
rect 13964 21428 13970 21480
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 15749 21471 15807 21477
rect 15749 21468 15761 21471
rect 14056 21440 15761 21468
rect 14056 21428 14062 21440
rect 15749 21437 15761 21440
rect 15795 21437 15807 21471
rect 15856 21468 15884 21576
rect 15948 21545 15976 21644
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 21910 21632 21916 21684
rect 21968 21672 21974 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 21968 21644 22477 21672
rect 21968 21632 21974 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 20254 21604 20260 21616
rect 16040 21576 20260 21604
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 16040 21468 16068 21576
rect 20254 21564 20260 21576
rect 20312 21564 20318 21616
rect 21818 21564 21824 21616
rect 21876 21604 21882 21616
rect 22833 21607 22891 21613
rect 22833 21604 22845 21607
rect 21876 21576 22845 21604
rect 21876 21564 21882 21576
rect 22833 21573 22845 21576
rect 22879 21573 22891 21607
rect 22833 21567 22891 21573
rect 17310 21536 17316 21548
rect 17271 21508 17316 21536
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 18046 21536 18052 21548
rect 18007 21508 18052 21536
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 18598 21496 18604 21548
rect 18656 21536 18662 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18656 21508 18705 21536
rect 18656 21496 18662 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 16206 21468 16212 21480
rect 15856 21440 16068 21468
rect 16167 21440 16212 21468
rect 15749 21431 15807 21437
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 17497 21471 17555 21477
rect 17497 21437 17509 21471
rect 17543 21468 17555 21471
rect 18230 21468 18236 21480
rect 17543 21440 18236 21468
rect 17543 21437 17555 21440
rect 17497 21431 17555 21437
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 18380 21440 18521 21468
rect 18380 21428 18386 21440
rect 18509 21437 18521 21440
rect 18555 21468 18567 21471
rect 19429 21471 19487 21477
rect 19429 21468 19441 21471
rect 18555 21440 19441 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 19429 21437 19441 21440
rect 19475 21437 19487 21471
rect 19429 21431 19487 21437
rect 22281 21471 22339 21477
rect 22281 21437 22293 21471
rect 22327 21437 22339 21471
rect 22281 21431 22339 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21468 22707 21471
rect 23017 21471 23075 21477
rect 23017 21468 23029 21471
rect 22695 21440 23029 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 23017 21437 23029 21440
rect 23063 21468 23075 21471
rect 23290 21468 23296 21480
rect 23063 21440 23296 21468
rect 23063 21437 23075 21440
rect 23017 21431 23075 21437
rect 12526 21400 12532 21412
rect 12452 21372 12532 21400
rect 10744 21363 10808 21369
rect 10744 21360 10750 21363
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 12704 21403 12762 21409
rect 12704 21369 12716 21403
rect 12750 21400 12762 21403
rect 13078 21400 13084 21412
rect 12750 21372 13084 21400
rect 12750 21369 12762 21372
rect 12704 21363 12762 21369
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 14182 21409 14188 21412
rect 14176 21400 14188 21409
rect 14143 21372 14188 21400
rect 14176 21363 14188 21372
rect 14182 21360 14188 21363
rect 14240 21360 14246 21412
rect 18248 21400 18276 21428
rect 19242 21400 19248 21412
rect 18248 21372 19248 21400
rect 19242 21360 19248 21372
rect 19300 21360 19306 21412
rect 11054 21332 11060 21344
rect 10520 21304 11060 21332
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11146 21292 11152 21344
rect 11204 21332 11210 21344
rect 11885 21335 11943 21341
rect 11885 21332 11897 21335
rect 11204 21304 11897 21332
rect 11204 21292 11210 21304
rect 11885 21301 11897 21304
rect 11931 21301 11943 21335
rect 11885 21295 11943 21301
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 14516 21304 15301 21332
rect 14516 21292 14522 21304
rect 15289 21301 15301 21304
rect 15335 21301 15347 21335
rect 15289 21295 15347 21301
rect 15378 21292 15384 21344
rect 15436 21332 15442 21344
rect 15436 21304 15481 21332
rect 15436 21292 15442 21304
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 15841 21335 15899 21341
rect 15841 21332 15853 21335
rect 15804 21304 15853 21332
rect 15804 21292 15810 21304
rect 15841 21301 15853 21304
rect 15887 21301 15899 21335
rect 15841 21295 15899 21301
rect 16393 21335 16451 21341
rect 16393 21301 16405 21335
rect 16439 21332 16451 21335
rect 16574 21332 16580 21344
rect 16439 21304 16580 21332
rect 16439 21301 16451 21304
rect 16393 21295 16451 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 16669 21335 16727 21341
rect 16669 21301 16681 21335
rect 16715 21332 16727 21335
rect 16850 21332 16856 21344
rect 16715 21304 16856 21332
rect 16715 21301 16727 21304
rect 16669 21295 16727 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 17034 21332 17040 21344
rect 16995 21304 17040 21332
rect 17034 21292 17040 21304
rect 17092 21292 17098 21344
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 22189 21335 22247 21341
rect 17184 21304 17229 21332
rect 17184 21292 17190 21304
rect 22189 21301 22201 21335
rect 22235 21332 22247 21335
rect 22296 21332 22324 21431
rect 23290 21428 23296 21440
rect 23348 21428 23354 21480
rect 22554 21332 22560 21344
rect 22235 21304 22560 21332
rect 22235 21301 22247 21304
rect 22189 21295 22247 21301
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 1104 21242 23460 21264
rect 1104 21190 8446 21242
rect 8498 21190 8510 21242
rect 8562 21190 8574 21242
rect 8626 21190 8638 21242
rect 8690 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 23460 21242
rect 1104 21168 23460 21190
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 1765 21131 1823 21137
rect 1765 21128 1777 21131
rect 1636 21100 1777 21128
rect 1636 21088 1642 21100
rect 1765 21097 1777 21100
rect 1811 21097 1823 21131
rect 1765 21091 1823 21097
rect 2222 21088 2228 21140
rect 2280 21128 2286 21140
rect 3605 21131 3663 21137
rect 3605 21128 3617 21131
rect 2280 21100 3617 21128
rect 2280 21088 2286 21100
rect 3605 21097 3617 21100
rect 3651 21097 3663 21131
rect 3605 21091 3663 21097
rect 3881 21131 3939 21137
rect 3881 21097 3893 21131
rect 3927 21128 3939 21131
rect 5074 21128 5080 21140
rect 3927 21100 5080 21128
rect 3927 21097 3939 21100
rect 3881 21091 3939 21097
rect 2590 21060 2596 21072
rect 1964 21032 2596 21060
rect 1964 21001 1992 21032
rect 2590 21020 2596 21032
rect 2648 21060 2654 21072
rect 2648 21032 3372 21060
rect 2648 21020 2654 21032
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20961 1639 20995
rect 1581 20955 1639 20961
rect 1949 20995 2007 21001
rect 1949 20961 1961 20995
rect 1995 20961 2007 20995
rect 1949 20955 2007 20961
rect 2216 20995 2274 21001
rect 2216 20961 2228 20995
rect 2262 20992 2274 20995
rect 2958 20992 2964 21004
rect 2262 20964 2964 20992
rect 2262 20961 2274 20964
rect 2216 20955 2274 20961
rect 1489 20791 1547 20797
rect 1489 20757 1501 20791
rect 1535 20788 1547 20791
rect 1596 20788 1624 20955
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 3344 20924 3372 21032
rect 3421 20995 3479 21001
rect 3421 20961 3433 20995
rect 3467 20992 3479 20995
rect 3896 20992 3924 21091
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 5442 21088 5448 21100
rect 5500 21128 5506 21140
rect 5500 21100 5764 21128
rect 5500 21088 5506 21100
rect 4154 21020 4160 21072
rect 4212 21060 4218 21072
rect 4310 21063 4368 21069
rect 4310 21060 4322 21063
rect 4212 21032 4322 21060
rect 4212 21020 4218 21032
rect 4310 21029 4322 21032
rect 4356 21029 4368 21063
rect 4310 21023 4368 21029
rect 4522 21020 4528 21072
rect 4580 21060 4586 21072
rect 5736 21069 5764 21100
rect 5810 21088 5816 21140
rect 5868 21128 5874 21140
rect 5905 21131 5963 21137
rect 5905 21128 5917 21131
rect 5868 21100 5917 21128
rect 5868 21088 5874 21100
rect 5905 21097 5917 21100
rect 5951 21097 5963 21131
rect 5905 21091 5963 21097
rect 5994 21088 6000 21140
rect 6052 21128 6058 21140
rect 6089 21131 6147 21137
rect 6089 21128 6101 21131
rect 6052 21100 6101 21128
rect 6052 21088 6058 21100
rect 6089 21097 6101 21100
rect 6135 21128 6147 21131
rect 6638 21128 6644 21140
rect 6135 21100 6644 21128
rect 6135 21097 6147 21100
rect 6089 21091 6147 21097
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 7561 21131 7619 21137
rect 7561 21097 7573 21131
rect 7607 21097 7619 21131
rect 7561 21091 7619 21097
rect 9309 21131 9367 21137
rect 9309 21097 9321 21131
rect 9355 21128 9367 21131
rect 10134 21128 10140 21140
rect 9355 21100 10140 21128
rect 9355 21097 9367 21100
rect 9309 21091 9367 21097
rect 6454 21069 6460 21072
rect 5721 21063 5779 21069
rect 4580 21032 5672 21060
rect 4580 21020 4586 21032
rect 5166 20992 5172 21004
rect 3467 20964 3924 20992
rect 4080 20964 5172 20992
rect 3467 20961 3479 20964
rect 3421 20955 3479 20961
rect 3970 20924 3976 20936
rect 3344 20896 3976 20924
rect 3970 20884 3976 20896
rect 4028 20924 4034 20936
rect 4080 20933 4108 20964
rect 5166 20952 5172 20964
rect 5224 20952 5230 21004
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20961 5595 20995
rect 5644 20992 5672 21032
rect 5721 21029 5733 21063
rect 5767 21029 5779 21063
rect 6448 21060 6460 21069
rect 6415 21032 6460 21060
rect 5721 21023 5779 21029
rect 6448 21023 6460 21032
rect 6454 21020 6460 21023
rect 6512 21020 6518 21072
rect 7576 21060 7604 21091
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 11054 21128 11060 21140
rect 11015 21100 11060 21128
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 11609 21131 11667 21137
rect 11609 21097 11621 21131
rect 11655 21128 11667 21131
rect 11882 21128 11888 21140
rect 11655 21100 11888 21128
rect 11655 21097 11667 21100
rect 11609 21091 11667 21097
rect 7920 21063 7978 21069
rect 7920 21060 7932 21063
rect 7576 21032 7932 21060
rect 7920 21029 7932 21032
rect 7966 21060 7978 21063
rect 8110 21060 8116 21072
rect 7966 21032 8116 21060
rect 7966 21029 7978 21032
rect 7920 21023 7978 21029
rect 8110 21020 8116 21032
rect 8168 21020 8174 21072
rect 9030 21020 9036 21072
rect 9088 21060 9094 21072
rect 9214 21060 9220 21072
rect 9088 21032 9220 21060
rect 9088 21020 9094 21032
rect 9214 21020 9220 21032
rect 9272 21060 9278 21072
rect 9272 21032 10548 21060
rect 9272 21020 9278 21032
rect 9692 21001 9720 21032
rect 10520 21004 10548 21032
rect 9677 20995 9735 21001
rect 5644 20964 9168 20992
rect 5537 20955 5595 20961
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 4028 20896 4077 20924
rect 4028 20884 4034 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 5552 20924 5580 20955
rect 5810 20924 5816 20936
rect 5552 20896 5816 20924
rect 4065 20887 4123 20893
rect 5810 20884 5816 20896
rect 5868 20884 5874 20936
rect 6178 20884 6184 20936
rect 6236 20933 6242 20936
rect 6236 20924 6246 20933
rect 6236 20896 6281 20924
rect 6236 20887 6246 20896
rect 6236 20884 6242 20887
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7653 20927 7711 20933
rect 7653 20924 7665 20927
rect 7248 20896 7665 20924
rect 7248 20884 7254 20896
rect 7653 20893 7665 20896
rect 7699 20893 7711 20927
rect 7653 20887 7711 20893
rect 3329 20859 3387 20865
rect 3329 20825 3341 20859
rect 3375 20856 3387 20859
rect 3375 20828 3924 20856
rect 3375 20825 3387 20828
rect 3329 20819 3387 20825
rect 3786 20788 3792 20800
rect 1535 20760 3792 20788
rect 1535 20757 1547 20760
rect 1489 20751 1547 20757
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 3896 20788 3924 20828
rect 4338 20788 4344 20800
rect 3896 20760 4344 20788
rect 4338 20748 4344 20760
rect 4396 20748 4402 20800
rect 5166 20748 5172 20800
rect 5224 20788 5230 20800
rect 6178 20788 6184 20800
rect 5224 20760 6184 20788
rect 5224 20748 5230 20760
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 8386 20748 8392 20800
rect 8444 20788 8450 20800
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8444 20760 9045 20788
rect 8444 20748 8450 20760
rect 9033 20757 9045 20760
rect 9079 20757 9091 20791
rect 9140 20788 9168 20964
rect 9677 20961 9689 20995
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 9933 20995 9991 21001
rect 9933 20992 9945 20995
rect 9824 20964 9945 20992
rect 9824 20952 9830 20964
rect 9933 20961 9945 20964
rect 9979 20961 9991 20995
rect 9933 20955 9991 20961
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 11149 20995 11207 21001
rect 10560 20964 10732 20992
rect 10560 20952 10566 20964
rect 10704 20924 10732 20964
rect 11149 20961 11161 20995
rect 11195 20992 11207 20995
rect 11624 20992 11652 21091
rect 11882 21088 11888 21100
rect 11940 21088 11946 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 14182 21088 14188 21140
rect 14240 21128 14246 21140
rect 14553 21131 14611 21137
rect 14553 21128 14565 21131
rect 14240 21100 14565 21128
rect 14240 21088 14246 21100
rect 14553 21097 14565 21100
rect 14599 21097 14611 21131
rect 16669 21131 16727 21137
rect 14553 21091 14611 21097
rect 14660 21100 15700 21128
rect 11968 21063 12026 21069
rect 11968 21029 11980 21063
rect 12014 21060 12026 21063
rect 13170 21060 13176 21072
rect 12014 21032 13176 21060
rect 12014 21029 12026 21032
rect 11968 21023 12026 21029
rect 13170 21020 13176 21032
rect 13228 21020 13234 21072
rect 13440 21063 13498 21069
rect 13440 21029 13452 21063
rect 13486 21060 13498 21063
rect 13722 21060 13728 21072
rect 13486 21032 13728 21060
rect 13486 21029 13498 21032
rect 13440 21023 13498 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 11195 20964 11652 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 14660 20992 14688 21100
rect 14737 21063 14795 21069
rect 14737 21029 14749 21063
rect 14783 21060 14795 21063
rect 15102 21060 15108 21072
rect 14783 21032 15108 21060
rect 14783 21029 14795 21032
rect 14737 21023 14795 21029
rect 15102 21020 15108 21032
rect 15160 21020 15166 21072
rect 15562 21001 15568 21004
rect 11848 20964 14688 20992
rect 14921 20995 14979 21001
rect 11848 20952 11854 20964
rect 14921 20961 14933 20995
rect 14967 20992 14979 20995
rect 15556 20992 15568 21001
rect 14967 20964 15568 20992
rect 14967 20961 14979 20964
rect 14921 20955 14979 20961
rect 15556 20955 15568 20964
rect 15562 20952 15568 20955
rect 15620 20952 15626 21004
rect 15672 20992 15700 21100
rect 16669 21097 16681 21131
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 16684 21060 16712 21091
rect 17310 21088 17316 21140
rect 17368 21128 17374 21140
rect 18141 21131 18199 21137
rect 18141 21128 18153 21131
rect 17368 21100 18153 21128
rect 17368 21088 17374 21100
rect 18141 21097 18153 21100
rect 18187 21097 18199 21131
rect 18141 21091 18199 21097
rect 17006 21063 17064 21069
rect 17006 21060 17018 21063
rect 16684 21032 17018 21060
rect 17006 21029 17018 21032
rect 17052 21060 17064 21063
rect 17218 21060 17224 21072
rect 17052 21032 17224 21060
rect 17052 21029 17064 21032
rect 17006 21023 17064 21029
rect 17218 21020 17224 21032
rect 17276 21020 17282 21072
rect 18156 21060 18184 21091
rect 22002 21088 22008 21140
rect 22060 21128 22066 21140
rect 22833 21131 22891 21137
rect 22833 21128 22845 21131
rect 22060 21100 22845 21128
rect 22060 21088 22066 21100
rect 22833 21097 22845 21100
rect 22879 21097 22891 21131
rect 22833 21091 22891 21097
rect 18478 21063 18536 21069
rect 18478 21060 18490 21063
rect 18156 21032 18490 21060
rect 18478 21029 18490 21032
rect 18524 21029 18536 21063
rect 18478 21023 18536 21029
rect 22189 21063 22247 21069
rect 22189 21029 22201 21063
rect 22235 21060 22247 21063
rect 22235 21032 22692 21060
rect 22235 21029 22247 21032
rect 22189 21023 22247 21029
rect 21542 20992 21548 21004
rect 15672 20964 21548 20992
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 22664 21001 22692 21032
rect 22281 20995 22339 21001
rect 22281 20961 22293 20995
rect 22327 20961 22339 20995
rect 22281 20955 22339 20961
rect 22649 20995 22707 21001
rect 22649 20961 22661 20995
rect 22695 20992 22707 20995
rect 23658 20992 23664 21004
rect 22695 20964 23664 20992
rect 22695 20961 22707 20964
rect 22649 20955 22707 20961
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 10704 20896 11713 20924
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 15105 20927 15163 20933
rect 15105 20893 15117 20927
rect 15151 20924 15163 20927
rect 15194 20924 15200 20936
rect 15151 20896 15200 20924
rect 15151 20893 15163 20896
rect 15105 20887 15163 20893
rect 11606 20856 11612 20868
rect 10612 20828 11612 20856
rect 10612 20788 10640 20828
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 11330 20788 11336 20800
rect 9140 20760 10640 20788
rect 11291 20760 11336 20788
rect 9033 20751 9091 20757
rect 11330 20748 11336 20760
rect 11388 20748 11394 20800
rect 11716 20788 11744 20887
rect 12618 20788 12624 20800
rect 11716 20760 12624 20788
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13188 20788 13216 20887
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15289 20927 15347 20933
rect 15289 20893 15301 20927
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 16761 20927 16819 20933
rect 16761 20893 16773 20927
rect 16807 20893 16819 20927
rect 18046 20924 18052 20936
rect 16761 20887 16819 20893
rect 17788 20896 18052 20924
rect 15304 20856 15332 20887
rect 14384 20828 15332 20856
rect 14384 20800 14412 20828
rect 13906 20788 13912 20800
rect 13188 20760 13912 20788
rect 13906 20748 13912 20760
rect 13964 20788 13970 20800
rect 14366 20788 14372 20800
rect 13964 20760 14372 20788
rect 13964 20748 13970 20760
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 16776 20788 16804 20887
rect 17402 20788 17408 20800
rect 16776 20760 17408 20788
rect 17402 20748 17408 20760
rect 17460 20788 17466 20800
rect 17788 20788 17816 20896
rect 18046 20884 18052 20896
rect 18104 20924 18110 20936
rect 18233 20927 18291 20933
rect 18233 20924 18245 20927
rect 18104 20896 18245 20924
rect 18104 20884 18110 20896
rect 18233 20893 18245 20896
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 17460 20760 17816 20788
rect 17460 20748 17466 20760
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19613 20791 19671 20797
rect 19613 20788 19625 20791
rect 19576 20760 19625 20788
rect 19576 20748 19582 20760
rect 19613 20757 19625 20760
rect 19659 20757 19671 20791
rect 22296 20788 22324 20955
rect 23658 20952 23664 20964
rect 23716 20952 23722 21004
rect 22465 20859 22523 20865
rect 22465 20825 22477 20859
rect 22511 20856 22523 20859
rect 23569 20859 23627 20865
rect 23569 20856 23581 20859
rect 22511 20828 23581 20856
rect 22511 20825 22523 20828
rect 22465 20819 22523 20825
rect 23569 20825 23581 20828
rect 23615 20825 23627 20859
rect 23569 20819 23627 20825
rect 23109 20791 23167 20797
rect 23109 20788 23121 20791
rect 22296 20760 23121 20788
rect 19613 20751 19671 20757
rect 23109 20757 23121 20760
rect 23155 20788 23167 20791
rect 23198 20788 23204 20800
rect 23155 20760 23204 20788
rect 23155 20757 23167 20760
rect 23109 20751 23167 20757
rect 23198 20748 23204 20760
rect 23256 20748 23262 20800
rect 1104 20698 23460 20720
rect 1104 20646 4714 20698
rect 4766 20646 4778 20698
rect 4830 20646 4842 20698
rect 4894 20646 4906 20698
rect 4958 20646 12178 20698
rect 12230 20646 12242 20698
rect 12294 20646 12306 20698
rect 12358 20646 12370 20698
rect 12422 20646 19642 20698
rect 19694 20646 19706 20698
rect 19758 20646 19770 20698
rect 19822 20646 19834 20698
rect 19886 20646 23460 20698
rect 1104 20624 23460 20646
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3510 20544 3516 20596
rect 3568 20584 3574 20596
rect 4893 20587 4951 20593
rect 4893 20584 4905 20587
rect 3568 20556 4905 20584
rect 3568 20544 3574 20556
rect 4893 20553 4905 20556
rect 4939 20553 4951 20587
rect 4893 20547 4951 20553
rect 5000 20556 6132 20584
rect 3712 20488 4568 20516
rect 3712 20460 3740 20488
rect 1578 20448 1584 20460
rect 1539 20420 1584 20448
rect 1578 20408 1584 20420
rect 1636 20408 1642 20460
rect 3142 20408 3148 20460
rect 3200 20448 3206 20460
rect 3694 20448 3700 20460
rect 3200 20420 3700 20448
rect 3200 20408 3206 20420
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 4338 20448 4344 20460
rect 4299 20420 4344 20448
rect 4338 20408 4344 20420
rect 4396 20408 4402 20460
rect 4540 20457 4568 20488
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20448 4583 20451
rect 5000 20448 5028 20556
rect 6104 20516 6132 20556
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6512 20556 6561 20584
rect 6512 20544 6518 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 6638 20544 6644 20596
rect 6696 20584 6702 20596
rect 10686 20584 10692 20596
rect 6696 20556 8064 20584
rect 6696 20544 6702 20556
rect 6914 20516 6920 20528
rect 6104 20488 6920 20516
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 8036 20516 8064 20556
rect 9324 20556 10272 20584
rect 10647 20556 10692 20584
rect 9324 20516 9352 20556
rect 8036 20488 9352 20516
rect 10244 20516 10272 20556
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 13078 20584 13084 20596
rect 10836 20556 13084 20584
rect 10836 20544 10842 20556
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13722 20584 13728 20596
rect 13228 20556 13728 20584
rect 13228 20544 13234 20556
rect 13722 20544 13728 20556
rect 13780 20584 13786 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13780 20556 13829 20584
rect 13780 20544 13786 20556
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 15378 20584 15384 20596
rect 13817 20547 13875 20553
rect 13924 20556 15384 20584
rect 11882 20516 11888 20528
rect 10244 20488 11888 20516
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 5166 20448 5172 20460
rect 4571 20420 5028 20448
rect 5127 20420 5172 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 6270 20408 6276 20460
rect 6328 20448 6334 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6328 20420 6837 20448
rect 6328 20408 6334 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 9214 20408 9220 20460
rect 9272 20448 9278 20460
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 9272 20420 9321 20448
rect 9272 20408 9278 20420
rect 9309 20417 9321 20420
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 11333 20451 11391 20457
rect 11333 20448 11345 20451
rect 10928 20420 11345 20448
rect 10928 20408 10934 20420
rect 11333 20417 11345 20420
rect 11379 20417 11391 20451
rect 13924 20448 13952 20556
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15620 20556 15761 20584
rect 15620 20544 15626 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 16669 20587 16727 20593
rect 16669 20553 16681 20587
rect 16715 20584 16727 20587
rect 17126 20584 17132 20596
rect 16715 20556 17132 20584
rect 16715 20553 16727 20556
rect 16669 20547 16727 20553
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19484 20556 19533 20584
rect 19484 20544 19490 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 22462 20584 22468 20596
rect 22423 20556 22468 20584
rect 19521 20547 19579 20553
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 16850 20476 16856 20528
rect 16908 20516 16914 20528
rect 17678 20516 17684 20528
rect 16908 20488 17684 20516
rect 16908 20476 16914 20488
rect 17678 20476 17684 20488
rect 17736 20516 17742 20528
rect 17736 20488 18000 20516
rect 17736 20476 17742 20488
rect 11333 20411 11391 20417
rect 13648 20420 13952 20448
rect 2958 20340 2964 20392
rect 3016 20380 3022 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3016 20352 3433 20380
rect 3016 20340 3022 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 4154 20340 4160 20392
rect 4212 20380 4218 20392
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 4212 20352 4261 20380
rect 4212 20340 4218 20352
rect 4249 20349 4261 20352
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 4982 20380 4988 20392
rect 4755 20352 4988 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 5436 20383 5494 20389
rect 5436 20349 5448 20383
rect 5482 20380 5494 20383
rect 5902 20380 5908 20392
rect 5482 20352 5908 20380
rect 5482 20349 5494 20352
rect 5436 20343 5494 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 6730 20380 6736 20392
rect 6236 20352 6736 20380
rect 6236 20340 6242 20352
rect 6730 20340 6736 20352
rect 6788 20380 6794 20392
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 6788 20352 7113 20380
rect 6788 20340 6794 20352
rect 7101 20349 7113 20352
rect 7147 20380 7159 20383
rect 7190 20380 7196 20392
rect 7147 20352 7196 20380
rect 7147 20349 7159 20352
rect 7101 20343 7159 20349
rect 7190 20340 7196 20352
rect 7248 20340 7254 20392
rect 7368 20383 7426 20389
rect 7368 20349 7380 20383
rect 7414 20380 7426 20383
rect 7926 20380 7932 20392
rect 7414 20352 7932 20380
rect 7414 20349 7426 20352
rect 7368 20343 7426 20349
rect 7926 20340 7932 20352
rect 7984 20380 7990 20392
rect 8386 20380 8392 20392
rect 7984 20352 8392 20380
rect 7984 20340 7990 20352
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20380 8631 20383
rect 9576 20383 9634 20389
rect 8619 20352 9076 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 1848 20315 1906 20321
rect 1848 20281 1860 20315
rect 1894 20312 1906 20315
rect 3513 20315 3571 20321
rect 3513 20312 3525 20315
rect 1894 20284 3525 20312
rect 1894 20281 1906 20284
rect 1848 20275 1906 20281
rect 2976 20256 3004 20284
rect 3513 20281 3525 20284
rect 3559 20281 3571 20315
rect 3513 20275 3571 20281
rect 5626 20272 5632 20324
rect 5684 20312 5690 20324
rect 9048 20321 9076 20352
rect 9576 20349 9588 20383
rect 9622 20380 9634 20383
rect 10410 20380 10416 20392
rect 9622 20352 10416 20380
rect 9622 20349 9634 20352
rect 9576 20343 9634 20349
rect 9692 20324 9720 20352
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10594 20340 10600 20392
rect 10652 20380 10658 20392
rect 11149 20383 11207 20389
rect 11149 20380 11161 20383
rect 10652 20352 11161 20380
rect 10652 20340 10658 20352
rect 11149 20349 11161 20352
rect 11195 20349 11207 20383
rect 11149 20343 11207 20349
rect 11977 20383 12035 20389
rect 11977 20349 11989 20383
rect 12023 20349 12035 20383
rect 11977 20343 12035 20349
rect 9033 20315 9091 20321
rect 5684 20284 8800 20312
rect 5684 20272 5690 20284
rect 2958 20204 2964 20256
rect 3016 20204 3022 20256
rect 3050 20204 3056 20256
rect 3108 20244 3114 20256
rect 3878 20244 3884 20256
rect 3108 20216 3153 20244
rect 3839 20216 3884 20244
rect 3108 20204 3114 20216
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 8772 20253 8800 20284
rect 9033 20281 9045 20315
rect 9079 20312 9091 20315
rect 9306 20312 9312 20324
rect 9079 20284 9312 20312
rect 9079 20281 9091 20284
rect 9033 20275 9091 20281
rect 9306 20272 9312 20284
rect 9364 20272 9370 20324
rect 9674 20272 9680 20324
rect 9732 20272 9738 20324
rect 11241 20315 11299 20321
rect 11241 20312 11253 20315
rect 9784 20284 11253 20312
rect 8481 20247 8539 20253
rect 8481 20244 8493 20247
rect 7064 20216 8493 20244
rect 7064 20204 7070 20216
rect 8481 20213 8493 20216
rect 8527 20213 8539 20247
rect 8481 20207 8539 20213
rect 8757 20247 8815 20253
rect 8757 20213 8769 20247
rect 8803 20213 8815 20247
rect 8757 20207 8815 20213
rect 8846 20204 8852 20256
rect 8904 20244 8910 20256
rect 9784 20244 9812 20284
rect 11241 20281 11253 20284
rect 11287 20281 11299 20315
rect 11992 20312 12020 20343
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12704 20383 12762 20389
rect 12492 20352 12537 20380
rect 12492 20340 12498 20352
rect 12704 20349 12716 20383
rect 12750 20380 12762 20383
rect 13538 20380 13544 20392
rect 12750 20352 13544 20380
rect 12750 20349 12762 20352
rect 12704 20343 12762 20349
rect 13538 20340 13544 20352
rect 13596 20340 13602 20392
rect 13648 20312 13676 20420
rect 15654 20408 15660 20460
rect 15712 20448 15718 20460
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 15712 20420 16405 20448
rect 15712 20408 15718 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 16393 20411 16451 20417
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20380 13967 20383
rect 14182 20380 14188 20392
rect 13955 20352 14188 20380
rect 13955 20349 13967 20352
rect 13909 20343 13967 20349
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 14366 20380 14372 20392
rect 14327 20352 14372 20380
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 16209 20383 16267 20389
rect 16209 20380 16221 20383
rect 14476 20352 16221 20380
rect 14476 20312 14504 20352
rect 16209 20349 16221 20352
rect 16255 20349 16267 20383
rect 16209 20343 16267 20349
rect 16574 20340 16580 20392
rect 16632 20380 16638 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16632 20352 17141 20380
rect 16632 20340 16638 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17494 20380 17500 20392
rect 17455 20352 17500 20380
rect 17129 20343 17187 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 11992 20284 13676 20312
rect 13740 20284 14504 20312
rect 11241 20275 11299 20281
rect 8904 20216 9812 20244
rect 8904 20204 8910 20216
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 10778 20244 10784 20256
rect 10100 20216 10784 20244
rect 10100 20204 10106 20216
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 12161 20247 12219 20253
rect 12161 20213 12173 20247
rect 12207 20244 12219 20247
rect 13740 20244 13768 20284
rect 14550 20272 14556 20324
rect 14608 20321 14614 20324
rect 14608 20315 14672 20321
rect 14608 20281 14626 20315
rect 14660 20281 14672 20315
rect 16301 20315 16359 20321
rect 16301 20312 16313 20315
rect 14608 20275 14672 20281
rect 15212 20284 16313 20312
rect 14608 20272 14614 20275
rect 12207 20216 13768 20244
rect 14093 20247 14151 20253
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 14093 20213 14105 20247
rect 14139 20244 14151 20247
rect 15212 20244 15240 20284
rect 16301 20281 16313 20284
rect 16347 20281 16359 20315
rect 16301 20275 16359 20281
rect 17037 20315 17095 20321
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17972 20312 18000 20488
rect 19058 20476 19064 20528
rect 19116 20516 19122 20528
rect 23474 20516 23480 20528
rect 19116 20488 23480 20516
rect 19116 20476 19122 20488
rect 23474 20476 23480 20488
rect 23532 20476 23538 20528
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 20073 20451 20131 20457
rect 18104 20420 18149 20448
rect 18104 20408 18110 20420
rect 20073 20417 20085 20451
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 18316 20383 18374 20389
rect 18316 20349 18328 20383
rect 18362 20380 18374 20383
rect 19518 20380 19524 20392
rect 18362 20352 19524 20380
rect 18362 20349 18374 20352
rect 18316 20343 18374 20349
rect 19518 20340 19524 20352
rect 19576 20380 19582 20392
rect 20088 20380 20116 20411
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22922 20448 22928 20460
rect 22428 20420 22928 20448
rect 22428 20408 22434 20420
rect 22922 20408 22928 20420
rect 22980 20408 22986 20460
rect 19576 20352 20116 20380
rect 22281 20383 22339 20389
rect 19576 20340 19582 20352
rect 22281 20349 22293 20383
rect 22327 20380 22339 20383
rect 22327 20352 22968 20380
rect 22327 20349 22339 20352
rect 22281 20343 22339 20349
rect 19889 20315 19947 20321
rect 19889 20312 19901 20315
rect 17083 20284 17172 20312
rect 17972 20284 19901 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 14139 20216 15240 20244
rect 15841 20247 15899 20253
rect 14139 20213 14151 20216
rect 14093 20207 14151 20213
rect 15841 20213 15853 20247
rect 15887 20244 15899 20247
rect 16482 20244 16488 20256
rect 15887 20216 16488 20244
rect 15887 20213 15899 20216
rect 15841 20207 15899 20213
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 17144 20244 17172 20284
rect 19889 20281 19901 20284
rect 19935 20281 19947 20315
rect 19889 20275 19947 20281
rect 22186 20272 22192 20324
rect 22244 20312 22250 20324
rect 22738 20312 22744 20324
rect 22244 20284 22744 20312
rect 22244 20272 22250 20284
rect 22738 20272 22744 20284
rect 22796 20272 22802 20324
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17144 20216 17693 20244
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 17920 20216 19441 20244
rect 17920 20204 17926 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 20036 20216 20081 20244
rect 20036 20204 20042 20216
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 22646 20244 22652 20256
rect 22152 20216 22197 20244
rect 22607 20216 22652 20244
rect 22152 20204 22158 20216
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 22940 20253 22968 20352
rect 22925 20247 22983 20253
rect 22925 20213 22937 20247
rect 22971 20244 22983 20247
rect 23566 20244 23572 20256
rect 22971 20216 23572 20244
rect 22971 20213 22983 20216
rect 22925 20207 22983 20213
rect 23566 20204 23572 20216
rect 23624 20204 23630 20256
rect 1104 20154 23460 20176
rect 1104 20102 8446 20154
rect 8498 20102 8510 20154
rect 8562 20102 8574 20154
rect 8626 20102 8638 20154
rect 8690 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 23460 20154
rect 1104 20080 23460 20102
rect 2958 20040 2964 20052
rect 2919 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 3936 20012 4445 20040
rect 3936 20000 3942 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 4893 20043 4951 20049
rect 4893 20009 4905 20043
rect 4939 20009 4951 20043
rect 4893 20003 4951 20009
rect 5721 20043 5779 20049
rect 5721 20009 5733 20043
rect 5767 20040 5779 20043
rect 8757 20043 8815 20049
rect 5767 20012 8248 20040
rect 5767 20009 5779 20012
rect 5721 20003 5779 20009
rect 1848 19975 1906 19981
rect 1848 19941 1860 19975
rect 1894 19972 1906 19975
rect 2866 19972 2872 19984
rect 1894 19944 2872 19972
rect 1894 19941 1906 19944
rect 1848 19935 1906 19941
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3050 19932 3056 19984
rect 3108 19972 3114 19984
rect 4525 19975 4583 19981
rect 4525 19972 4537 19975
rect 3108 19944 4537 19972
rect 3108 19932 3114 19944
rect 4525 19941 4537 19944
rect 4571 19941 4583 19975
rect 4908 19972 4936 20003
rect 6086 19972 6092 19984
rect 4908 19944 6092 19972
rect 4525 19935 4583 19941
rect 6086 19932 6092 19944
rect 6144 19932 6150 19984
rect 7006 19981 7012 19984
rect 7000 19972 7012 19981
rect 6967 19944 7012 19972
rect 7000 19935 7012 19944
rect 7006 19932 7012 19935
rect 7064 19932 7070 19984
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 3421 19907 3479 19913
rect 3421 19904 3433 19907
rect 2832 19876 3433 19904
rect 2832 19864 2838 19876
rect 3421 19873 3433 19876
rect 3467 19873 3479 19907
rect 3421 19867 3479 19873
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 5258 19904 5264 19916
rect 3660 19876 4835 19904
rect 5219 19876 5264 19904
rect 3660 19864 3666 19876
rect 3510 19836 3516 19848
rect 3471 19808 3516 19836
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 3697 19839 3755 19845
rect 3697 19805 3709 19839
rect 3743 19836 3755 19839
rect 3970 19836 3976 19848
rect 3743 19808 3976 19836
rect 3743 19805 3755 19808
rect 3697 19799 3755 19805
rect 3970 19796 3976 19808
rect 4028 19836 4034 19848
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 4028 19808 4721 19836
rect 4028 19796 4034 19808
rect 4709 19805 4721 19808
rect 4755 19805 4767 19839
rect 4807 19836 4835 19876
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5534 19864 5540 19916
rect 5592 19904 5598 19916
rect 8220 19913 8248 20012
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 8846 20040 8852 20052
rect 8803 20012 8852 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9677 20043 9735 20049
rect 9677 20009 9689 20043
rect 9723 20040 9735 20043
rect 10226 20040 10232 20052
rect 9723 20012 10232 20040
rect 9723 20009 9735 20012
rect 9677 20003 9735 20009
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 13814 20040 13820 20052
rect 13596 20012 13820 20040
rect 13596 20000 13602 20012
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14182 20040 14188 20052
rect 14143 20012 14188 20040
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 14550 20040 14556 20052
rect 14511 20012 14556 20040
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15252 20012 15761 20040
rect 15252 20000 15258 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 16206 20040 16212 20052
rect 16163 20012 16212 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 22278 20040 22284 20052
rect 16316 20012 22284 20040
rect 10045 19975 10103 19981
rect 10045 19972 10057 19975
rect 8864 19944 10057 19972
rect 8864 19916 8892 19944
rect 10045 19941 10057 19944
rect 10091 19972 10103 19975
rect 10965 19975 11023 19981
rect 10965 19972 10977 19975
rect 10091 19944 10977 19972
rect 10091 19941 10103 19944
rect 10045 19935 10103 19941
rect 10965 19941 10977 19944
rect 11011 19941 11023 19975
rect 10965 19935 11023 19941
rect 12526 19932 12532 19984
rect 12584 19972 12590 19984
rect 16316 19972 16344 20012
rect 22278 20000 22284 20012
rect 22336 20000 22342 20052
rect 22462 20040 22468 20052
rect 22423 20012 22468 20040
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 22830 20040 22836 20052
rect 22791 20012 22836 20040
rect 22830 20000 22836 20012
rect 22888 20000 22894 20052
rect 16574 19972 16580 19984
rect 12584 19944 16344 19972
rect 16535 19944 16580 19972
rect 12584 19932 12590 19944
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 17862 19981 17868 19984
rect 17313 19975 17371 19981
rect 17313 19972 17325 19975
rect 17092 19944 17325 19972
rect 17092 19932 17098 19944
rect 17313 19941 17325 19944
rect 17359 19941 17371 19975
rect 17856 19972 17868 19981
rect 17823 19944 17868 19972
rect 17313 19935 17371 19941
rect 17856 19935 17868 19944
rect 17862 19932 17868 19935
rect 17920 19932 17926 19984
rect 18046 19932 18052 19984
rect 18104 19972 18110 19984
rect 20898 19972 20904 19984
rect 18104 19944 20904 19972
rect 18104 19932 18110 19944
rect 20898 19932 20904 19944
rect 20956 19932 20962 19984
rect 21453 19975 21511 19981
rect 21453 19941 21465 19975
rect 21499 19972 21511 19975
rect 22370 19972 22376 19984
rect 21499 19944 22376 19972
rect 21499 19941 21511 19944
rect 21453 19935 21511 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 6641 19907 6699 19913
rect 5592 19876 6316 19904
rect 5592 19864 5598 19876
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 4807 19808 5365 19836
rect 4709 19799 4767 19805
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 5626 19836 5632 19848
rect 5491 19808 5632 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 3786 19728 3792 19780
rect 3844 19768 3850 19780
rect 4724 19768 4752 19799
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 6178 19836 6184 19848
rect 6139 19808 6184 19836
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 6288 19845 6316 19876
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 8205 19907 8263 19913
rect 6687 19876 7788 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 6273 19799 6331 19805
rect 5534 19768 5540 19780
rect 3844 19740 4292 19768
rect 4724 19740 5540 19768
rect 3844 19728 3850 19740
rect 3050 19660 3056 19712
rect 3108 19700 3114 19712
rect 4062 19700 4068 19712
rect 3108 19672 3153 19700
rect 4023 19672 4068 19700
rect 3108 19660 3114 19672
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4264 19700 4292 19740
rect 5534 19728 5540 19740
rect 5592 19768 5598 19780
rect 5718 19768 5724 19780
rect 5592 19740 5724 19768
rect 5592 19728 5598 19740
rect 5718 19728 5724 19740
rect 5776 19728 5782 19780
rect 5810 19728 5816 19780
rect 5868 19768 5874 19780
rect 6656 19768 6684 19867
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 7760 19836 7788 19876
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 8846 19864 8852 19916
rect 8904 19864 8910 19916
rect 9125 19907 9183 19913
rect 9125 19873 9137 19907
rect 9171 19904 9183 19907
rect 9306 19904 9312 19916
rect 9171 19876 9312 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 9214 19836 9220 19848
rect 6788 19808 6833 19836
rect 7760 19808 8524 19836
rect 9175 19808 9220 19836
rect 6788 19796 6794 19808
rect 5868 19740 6684 19768
rect 5868 19728 5874 19740
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 8389 19771 8447 19777
rect 8389 19768 8401 19771
rect 7892 19740 8401 19768
rect 7892 19728 7898 19740
rect 8389 19737 8401 19740
rect 8435 19737 8447 19771
rect 8389 19731 8447 19737
rect 6730 19700 6736 19712
rect 4264 19672 6736 19700
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7098 19660 7104 19712
rect 7156 19700 7162 19712
rect 8113 19703 8171 19709
rect 8113 19700 8125 19703
rect 7156 19672 8125 19700
rect 7156 19660 7162 19672
rect 8113 19669 8125 19672
rect 8159 19669 8171 19703
rect 8496 19700 8524 19808
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9674 19836 9680 19848
rect 9447 19808 9680 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10137 19839 10195 19845
rect 10137 19836 10149 19839
rect 10008 19808 10149 19836
rect 10008 19796 10014 19808
rect 10137 19805 10149 19808
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 8665 19771 8723 19777
rect 8665 19737 8677 19771
rect 8711 19768 8723 19771
rect 9122 19768 9128 19780
rect 8711 19740 9128 19768
rect 8711 19737 8723 19740
rect 8665 19731 8723 19737
rect 9122 19728 9128 19740
rect 9180 19728 9186 19780
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 10244 19768 10272 19799
rect 9824 19740 10272 19768
rect 10888 19768 10916 19867
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 12897 19907 12955 19913
rect 12897 19904 12909 19907
rect 12768 19876 12909 19904
rect 12768 19864 12774 19876
rect 12897 19873 12909 19876
rect 12943 19873 12955 19907
rect 13354 19904 13360 19916
rect 12897 19867 12955 19873
rect 13096 19876 13360 19904
rect 11146 19836 11152 19848
rect 11107 19808 11152 19836
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 12802 19836 12808 19848
rect 11296 19808 12808 19836
rect 11296 19796 11302 19808
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13096 19845 13124 19876
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13722 19904 13728 19916
rect 13683 19876 13728 19904
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 15470 19904 15476 19916
rect 13832 19876 15476 19904
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13832 19836 13860 19876
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15654 19904 15660 19916
rect 15615 19876 15660 19904
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 16482 19904 16488 19916
rect 16443 19876 16488 19904
rect 16482 19864 16488 19876
rect 16540 19904 16546 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 16540 19876 16957 19904
rect 16540 19864 16546 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 19058 19904 19064 19916
rect 16945 19867 17003 19873
rect 17052 19876 19064 19904
rect 13081 19799 13139 19805
rect 13188 19808 13860 19836
rect 11425 19771 11483 19777
rect 11425 19768 11437 19771
rect 10888 19740 11437 19768
rect 9824 19728 9830 19740
rect 11425 19737 11437 19740
rect 11471 19768 11483 19771
rect 13188 19768 13216 19808
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14645 19839 14703 19845
rect 13964 19808 14009 19836
rect 13964 19796 13970 19808
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 11471 19740 13216 19768
rect 13357 19771 13415 19777
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 13357 19737 13369 19771
rect 13403 19768 13415 19771
rect 14550 19768 14556 19780
rect 13403 19740 14556 19768
rect 13403 19737 13415 19740
rect 13357 19731 13415 19737
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 9858 19700 9864 19712
rect 8496 19672 9864 19700
rect 8113 19663 8171 19669
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 10505 19703 10563 19709
rect 10505 19669 10517 19703
rect 10551 19700 10563 19703
rect 11238 19700 11244 19712
rect 10551 19672 11244 19700
rect 10551 19669 10563 19672
rect 10505 19663 10563 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 14660 19700 14688 19799
rect 14734 19796 14740 19848
rect 14792 19836 14798 19848
rect 15838 19836 15844 19848
rect 14792 19808 14837 19836
rect 15799 19808 15844 19836
rect 14792 19796 14798 19808
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 16574 19836 16580 19848
rect 16224 19808 16580 19836
rect 15289 19771 15347 19777
rect 15289 19737 15301 19771
rect 15335 19768 15347 19771
rect 16224 19768 16252 19808
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 15335 19740 16252 19768
rect 15335 19737 15347 19740
rect 15289 19731 15347 19737
rect 16298 19728 16304 19780
rect 16356 19768 16362 19780
rect 16684 19768 16712 19799
rect 17052 19768 17080 19876
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 19613 19907 19671 19913
rect 19613 19873 19625 19907
rect 19659 19904 19671 19907
rect 20070 19904 20076 19916
rect 19659 19876 20076 19904
rect 19659 19873 19671 19876
rect 19613 19867 19671 19873
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 21358 19904 21364 19916
rect 21319 19876 21364 19904
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 22278 19904 22284 19916
rect 21959 19876 22140 19904
rect 22239 19876 22284 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 17402 19796 17408 19848
rect 17460 19836 17466 19848
rect 17586 19836 17592 19848
rect 17460 19808 17592 19836
rect 17460 19796 17466 19808
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 19426 19796 19432 19848
rect 19484 19836 19490 19848
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 19484 19808 19717 19836
rect 19484 19796 19490 19808
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 19935 19808 21557 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 16356 19740 16712 19768
rect 16776 19740 17080 19768
rect 21560 19768 21588 19799
rect 21910 19768 21916 19780
rect 21560 19740 21916 19768
rect 16356 19728 16362 19740
rect 12575 19672 14688 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 16776 19700 16804 19740
rect 21910 19728 21916 19740
rect 21968 19728 21974 19780
rect 22112 19768 22140 19876
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 22646 19904 22652 19916
rect 22559 19876 22652 19904
rect 22646 19864 22652 19876
rect 22704 19904 22710 19916
rect 23382 19904 23388 19916
rect 22704 19876 23388 19904
rect 22704 19864 22710 19876
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 22112 19740 23152 19768
rect 23124 19712 23152 19740
rect 17126 19700 17132 19712
rect 15896 19672 16804 19700
rect 17087 19672 17132 19700
rect 15896 19660 15902 19672
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18969 19703 19027 19709
rect 18969 19700 18981 19703
rect 18012 19672 18981 19700
rect 18012 19660 18018 19672
rect 18969 19669 18981 19672
rect 19015 19669 19027 19703
rect 18969 19663 19027 19669
rect 19245 19703 19303 19709
rect 19245 19669 19257 19703
rect 19291 19700 19303 19703
rect 20438 19700 20444 19712
rect 19291 19672 20444 19700
rect 19291 19669 19303 19672
rect 19245 19663 19303 19669
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 20990 19700 20996 19712
rect 20951 19672 20996 19700
rect 20990 19660 20996 19672
rect 21048 19660 21054 19712
rect 22097 19703 22155 19709
rect 22097 19669 22109 19703
rect 22143 19700 22155 19703
rect 22278 19700 22284 19712
rect 22143 19672 22284 19700
rect 22143 19669 22155 19672
rect 22097 19663 22155 19669
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 23106 19700 23112 19712
rect 23067 19672 23112 19700
rect 23106 19660 23112 19672
rect 23164 19660 23170 19712
rect 1104 19610 23460 19632
rect 1104 19558 4714 19610
rect 4766 19558 4778 19610
rect 4830 19558 4842 19610
rect 4894 19558 4906 19610
rect 4958 19558 12178 19610
rect 12230 19558 12242 19610
rect 12294 19558 12306 19610
rect 12358 19558 12370 19610
rect 12422 19558 19642 19610
rect 19694 19558 19706 19610
rect 19758 19558 19770 19610
rect 19822 19558 19834 19610
rect 19886 19558 23460 19610
rect 1104 19536 23460 19558
rect 2041 19499 2099 19505
rect 2041 19465 2053 19499
rect 2087 19496 2099 19499
rect 5258 19496 5264 19508
rect 2087 19468 5264 19496
rect 2087 19465 2099 19468
rect 2041 19459 2099 19465
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 10686 19496 10692 19508
rect 6788 19468 10692 19496
rect 6788 19456 6794 19468
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 10778 19456 10784 19508
rect 10836 19496 10842 19508
rect 10836 19468 12480 19496
rect 10836 19456 10842 19468
rect 12452 19440 12480 19468
rect 13078 19456 13084 19508
rect 13136 19496 13142 19508
rect 13814 19496 13820 19508
rect 13136 19468 13400 19496
rect 13775 19468 13820 19496
rect 13136 19456 13142 19468
rect 2409 19431 2467 19437
rect 2409 19397 2421 19431
rect 2455 19428 2467 19431
rect 3602 19428 3608 19440
rect 2455 19400 3608 19428
rect 2455 19397 2467 19400
rect 2409 19391 2467 19397
rect 3602 19388 3608 19400
rect 3660 19388 3666 19440
rect 3786 19388 3792 19440
rect 3844 19388 3850 19440
rect 12434 19388 12440 19440
rect 12492 19388 12498 19440
rect 13372 19428 13400 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 15010 19496 15016 19508
rect 14424 19468 15016 19496
rect 14424 19456 14430 19468
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 18046 19496 18052 19508
rect 15120 19468 18052 19496
rect 15120 19428 15148 19468
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 18966 19496 18972 19508
rect 18196 19468 18972 19496
rect 18196 19456 18202 19468
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 22830 19496 22836 19508
rect 19208 19468 22140 19496
rect 22791 19468 22836 19496
rect 19208 19456 19214 19468
rect 13372 19400 15148 19428
rect 15286 19388 15292 19440
rect 15344 19428 15350 19440
rect 15657 19431 15715 19437
rect 15657 19428 15669 19431
rect 15344 19400 15669 19428
rect 15344 19388 15350 19400
rect 15657 19397 15669 19400
rect 15703 19428 15715 19431
rect 15838 19428 15844 19440
rect 15703 19400 15844 19428
rect 15703 19397 15715 19400
rect 15657 19391 15715 19397
rect 15838 19388 15844 19400
rect 15896 19388 15902 19440
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 22112 19428 22140 19468
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 22738 19428 22744 19440
rect 17644 19400 18276 19428
rect 22112 19400 22744 19428
rect 17644 19388 17650 19400
rect 3142 19360 3148 19372
rect 3103 19332 3148 19360
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19261 1915 19295
rect 1857 19255 1915 19261
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19292 2283 19295
rect 3050 19292 3056 19304
rect 2271 19264 3056 19292
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 1872 19224 1900 19255
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 3804 19301 3832 19388
rect 3970 19360 3976 19372
rect 3931 19332 3976 19360
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19360 5135 19363
rect 5626 19360 5632 19372
rect 5123 19332 5632 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 5902 19360 5908 19372
rect 5863 19332 5908 19360
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 6104 19332 6408 19360
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19261 3847 19295
rect 3789 19255 3847 19261
rect 5813 19295 5871 19301
rect 5813 19261 5825 19295
rect 5859 19292 5871 19295
rect 6104 19292 6132 19332
rect 5859 19264 6132 19292
rect 5859 19261 5871 19264
rect 5813 19255 5871 19261
rect 6178 19252 6184 19304
rect 6236 19292 6242 19304
rect 6380 19292 6408 19332
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 7064 19332 7389 19360
rect 7064 19320 7070 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7834 19360 7840 19372
rect 7377 19323 7435 19329
rect 7484 19332 7840 19360
rect 7484 19292 7512 19332
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 8018 19369 8024 19372
rect 7976 19363 8024 19369
rect 7976 19329 7988 19363
rect 8022 19329 8024 19363
rect 7976 19323 8024 19329
rect 8018 19320 8024 19323
rect 8076 19320 8082 19372
rect 8116 19363 8174 19369
rect 8116 19329 8128 19363
rect 8162 19329 8174 19363
rect 8116 19323 8174 19329
rect 7650 19292 7656 19304
rect 6236 19264 6281 19292
rect 6380 19264 7512 19292
rect 7611 19264 7656 19292
rect 6236 19252 6242 19264
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 8128 19292 8156 19323
rect 14366 19320 14372 19372
rect 14424 19360 14430 19372
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 14424 19332 14565 19360
rect 14424 19320 14430 19332
rect 14553 19329 14565 19332
rect 14599 19360 14611 19363
rect 14734 19360 14740 19372
rect 14599 19332 14740 19360
rect 14599 19329 14611 19332
rect 14553 19323 14611 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15378 19360 15384 19372
rect 15339 19332 15384 19360
rect 15378 19320 15384 19332
rect 15436 19360 15442 19372
rect 15746 19360 15752 19372
rect 15436 19332 15752 19360
rect 15436 19320 15442 19332
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 16206 19360 16212 19372
rect 16167 19332 16212 19360
rect 16206 19320 16212 19332
rect 16264 19360 16270 19372
rect 16264 19332 16620 19360
rect 16264 19320 16270 19332
rect 7760 19264 8156 19292
rect 4062 19224 4068 19236
rect 1872 19196 4068 19224
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 5721 19227 5779 19233
rect 4540 19196 5672 19224
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2774 19156 2780 19168
rect 2639 19128 2780 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 2961 19159 3019 19165
rect 2961 19156 2973 19159
rect 2924 19128 2973 19156
rect 2924 19116 2930 19128
rect 2961 19125 2973 19128
rect 3007 19125 3019 19159
rect 2961 19119 3019 19125
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 3418 19156 3424 19168
rect 3108 19128 3153 19156
rect 3379 19128 3424 19156
rect 3108 19116 3114 19128
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 3602 19116 3608 19168
rect 3660 19156 3666 19168
rect 4540 19165 4568 19196
rect 3881 19159 3939 19165
rect 3881 19156 3893 19159
rect 3660 19128 3893 19156
rect 3660 19116 3666 19128
rect 3881 19125 3893 19128
rect 3927 19125 3939 19159
rect 3881 19119 3939 19125
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19125 4583 19159
rect 4525 19119 4583 19125
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 4893 19159 4951 19165
rect 4893 19156 4905 19159
rect 4672 19128 4905 19156
rect 4672 19116 4678 19128
rect 4893 19125 4905 19128
rect 4939 19125 4951 19159
rect 4893 19119 4951 19125
rect 4985 19159 5043 19165
rect 4985 19125 4997 19159
rect 5031 19156 5043 19159
rect 5166 19156 5172 19168
rect 5031 19128 5172 19156
rect 5031 19125 5043 19128
rect 4985 19119 5043 19125
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 5350 19156 5356 19168
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 5644 19156 5672 19196
rect 5721 19193 5733 19227
rect 5767 19224 5779 19227
rect 7760 19224 7788 19264
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8260 19264 8401 19292
rect 8260 19252 8266 19264
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19292 9827 19295
rect 10045 19295 10103 19301
rect 9815 19264 10002 19292
rect 9815 19261 9827 19264
rect 9769 19255 9827 19261
rect 9858 19224 9864 19236
rect 5767 19196 6408 19224
rect 5767 19193 5779 19196
rect 5721 19187 5779 19193
rect 6178 19156 6184 19168
rect 5644 19128 6184 19156
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 6380 19165 6408 19196
rect 7208 19196 7788 19224
rect 9508 19196 9864 19224
rect 7208 19168 7236 19196
rect 6365 19159 6423 19165
rect 6365 19125 6377 19159
rect 6411 19125 6423 19159
rect 6365 19119 6423 19125
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19156 6883 19159
rect 7006 19156 7012 19168
rect 6871 19128 7012 19156
rect 6871 19125 6883 19128
rect 6825 19119 6883 19125
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 9508 19165 9536 19196
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 7285 19159 7343 19165
rect 7285 19125 7297 19159
rect 7331 19156 7343 19159
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 7331 19128 9505 19156
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 9493 19119 9551 19125
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9974 19156 10002 19264
rect 10045 19261 10057 19295
rect 10091 19261 10103 19295
rect 10045 19255 10103 19261
rect 10312 19295 10370 19301
rect 10312 19261 10324 19295
rect 10358 19292 10370 19295
rect 11146 19292 11152 19304
rect 10358 19264 11152 19292
rect 10358 19261 10370 19264
rect 10312 19255 10370 19261
rect 10060 19224 10088 19255
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12526 19292 12532 19304
rect 12483 19264 12532 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 14332 19264 15209 19292
rect 14332 19252 14338 19264
rect 15197 19261 15209 19264
rect 15243 19292 15255 19295
rect 16298 19292 16304 19304
rect 15243 19264 16304 19292
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16390 19252 16396 19304
rect 16448 19292 16454 19304
rect 16492 19295 16550 19301
rect 16492 19292 16504 19295
rect 16448 19264 16504 19292
rect 16448 19252 16454 19264
rect 16492 19261 16504 19264
rect 16538 19261 16550 19295
rect 16592 19292 16620 19332
rect 16752 19295 16810 19301
rect 16592 19264 16712 19292
rect 16492 19255 16550 19261
rect 10962 19224 10968 19236
rect 10060 19196 10968 19224
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 11698 19224 11704 19236
rect 11659 19196 11704 19224
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 12710 19233 12716 19236
rect 12704 19224 12716 19233
rect 12671 19196 12716 19224
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 14369 19227 14427 19233
rect 14369 19193 14381 19227
rect 14415 19224 14427 19227
rect 16025 19227 16083 19233
rect 14415 19196 14872 19224
rect 14415 19193 14427 19196
rect 14369 19187 14427 19193
rect 11146 19156 11152 19168
rect 9732 19128 9777 19156
rect 9974 19128 11152 19156
rect 9732 19116 9738 19128
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11422 19156 11428 19168
rect 11383 19128 11428 19156
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 13998 19156 14004 19168
rect 13959 19128 14004 19156
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14458 19156 14464 19168
rect 14419 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14844 19165 14872 19196
rect 16025 19193 16037 19227
rect 16071 19224 16083 19227
rect 16574 19224 16580 19236
rect 16071 19196 16580 19224
rect 16071 19193 16083 19196
rect 16025 19187 16083 19193
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 16684 19224 16712 19264
rect 16752 19261 16764 19295
rect 16798 19292 16810 19295
rect 17954 19292 17960 19304
rect 16798 19264 17960 19292
rect 16798 19261 16810 19264
rect 16752 19255 16810 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 18248 19301 18276 19400
rect 22738 19388 22744 19400
rect 22796 19388 22802 19440
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 18966 19292 18972 19304
rect 18279 19264 18972 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 18966 19252 18972 19264
rect 19024 19292 19030 19304
rect 19705 19295 19763 19301
rect 19705 19292 19717 19295
rect 19024 19264 19717 19292
rect 19024 19252 19030 19264
rect 19705 19261 19717 19264
rect 19751 19292 19763 19295
rect 20806 19292 20812 19304
rect 19751 19264 20812 19292
rect 19751 19261 19763 19264
rect 19705 19255 19763 19261
rect 20806 19252 20812 19264
rect 20864 19292 20870 19304
rect 21177 19295 21235 19301
rect 21177 19292 21189 19295
rect 20864 19264 21189 19292
rect 20864 19252 20870 19264
rect 21177 19261 21189 19264
rect 21223 19261 21235 19295
rect 21177 19255 21235 19261
rect 22649 19295 22707 19301
rect 22649 19261 22661 19295
rect 22695 19292 22707 19295
rect 22695 19264 23060 19292
rect 22695 19261 22707 19264
rect 22649 19255 22707 19261
rect 18500 19227 18558 19233
rect 16684 19196 17908 19224
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19125 14887 19159
rect 14829 19119 14887 19125
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 16117 19159 16175 19165
rect 15344 19128 15389 19156
rect 15344 19116 15350 19128
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 17034 19156 17040 19168
rect 16163 19128 17040 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17880 19165 17908 19196
rect 18500 19193 18512 19227
rect 18546 19224 18558 19227
rect 19334 19224 19340 19236
rect 18546 19196 19340 19224
rect 18546 19193 18558 19196
rect 18500 19187 18558 19193
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 19972 19227 20030 19233
rect 19972 19193 19984 19227
rect 20018 19224 20030 19227
rect 20346 19224 20352 19236
rect 20018 19196 20352 19224
rect 20018 19193 20030 19196
rect 19972 19187 20030 19193
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 21444 19227 21502 19233
rect 21444 19193 21456 19227
rect 21490 19224 21502 19227
rect 22278 19224 22284 19236
rect 21490 19196 22284 19224
rect 21490 19193 21502 19196
rect 21444 19187 21502 19193
rect 22278 19184 22284 19196
rect 22336 19184 22342 19236
rect 23032 19168 23060 19264
rect 23382 19252 23388 19304
rect 23440 19292 23446 19304
rect 23569 19295 23627 19301
rect 23569 19292 23581 19295
rect 23440 19264 23581 19292
rect 23440 19252 23446 19264
rect 23569 19261 23581 19264
rect 23615 19261 23627 19295
rect 23569 19255 23627 19261
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19125 17923 19159
rect 17865 19119 17923 19125
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19576 19128 19625 19156
rect 19576 19116 19582 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 21082 19156 21088 19168
rect 21043 19128 21088 19156
rect 19613 19119 19671 19125
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 22557 19159 22615 19165
rect 22557 19156 22569 19159
rect 21692 19128 22569 19156
rect 21692 19116 21698 19128
rect 22557 19125 22569 19128
rect 22603 19125 22615 19159
rect 23014 19156 23020 19168
rect 22975 19128 23020 19156
rect 22557 19119 22615 19125
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 1104 19066 23460 19088
rect 1104 19014 8446 19066
rect 8498 19014 8510 19066
rect 8562 19014 8574 19066
rect 8626 19014 8638 19066
rect 8690 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 23460 19066
rect 1104 18992 23460 19014
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 3053 18955 3111 18961
rect 3053 18952 3065 18955
rect 2924 18924 3065 18952
rect 2924 18912 2930 18924
rect 3053 18921 3065 18924
rect 3099 18921 3111 18955
rect 3053 18915 3111 18921
rect 3145 18955 3203 18961
rect 3145 18921 3157 18955
rect 3191 18952 3203 18955
rect 3510 18952 3516 18964
rect 3191 18924 3516 18952
rect 3191 18921 3203 18924
rect 3145 18915 3203 18921
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 4249 18955 4307 18961
rect 4249 18921 4261 18955
rect 4295 18952 4307 18955
rect 4614 18952 4620 18964
rect 4295 18924 4620 18952
rect 4295 18921 4307 18924
rect 4249 18915 4307 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 4939 18924 5273 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 5261 18915 5319 18921
rect 6549 18955 6607 18961
rect 6549 18921 6561 18955
rect 6595 18952 6607 18955
rect 6730 18952 6736 18964
rect 6595 18924 6736 18952
rect 6595 18921 6607 18924
rect 6549 18915 6607 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7006 18952 7012 18964
rect 6967 18924 7012 18952
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8260 18924 9229 18952
rect 8260 18912 8266 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9950 18912 9956 18964
rect 10008 18952 10014 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 10008 18924 11529 18952
rect 10008 18912 10014 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 12986 18952 12992 18964
rect 12947 18924 12992 18952
rect 11517 18915 11575 18921
rect 12986 18912 12992 18924
rect 13044 18912 13050 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 14516 18924 15301 18952
rect 14516 18912 14522 18924
rect 15289 18921 15301 18924
rect 15335 18921 15347 18955
rect 15289 18915 15347 18921
rect 15562 18912 15568 18964
rect 15620 18952 15626 18964
rect 15657 18955 15715 18961
rect 15657 18952 15669 18955
rect 15620 18924 15669 18952
rect 15620 18912 15626 18924
rect 15657 18921 15669 18924
rect 15703 18921 15715 18955
rect 15657 18915 15715 18921
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 16632 18924 18521 18952
rect 16632 18912 16638 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 19978 18912 19984 18964
rect 20036 18912 20042 18964
rect 20346 18952 20352 18964
rect 20307 18924 20352 18952
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 22278 18952 22284 18964
rect 22239 18924 22284 18952
rect 22278 18912 22284 18924
rect 22336 18952 22342 18964
rect 22741 18955 22799 18961
rect 22741 18952 22753 18955
rect 22336 18924 22753 18952
rect 22336 18912 22342 18924
rect 22741 18921 22753 18924
rect 22787 18921 22799 18955
rect 22741 18915 22799 18921
rect 3418 18844 3424 18896
rect 3476 18884 3482 18896
rect 4801 18887 4859 18893
rect 3476 18856 4108 18884
rect 3476 18844 3482 18856
rect 1578 18776 1584 18828
rect 1636 18816 1642 18828
rect 1673 18819 1731 18825
rect 1673 18816 1685 18819
rect 1636 18788 1685 18816
rect 1636 18776 1642 18788
rect 1673 18785 1685 18788
rect 1719 18785 1731 18819
rect 1673 18779 1731 18785
rect 1940 18819 1998 18825
rect 1940 18785 1952 18819
rect 1986 18816 1998 18819
rect 3050 18816 3056 18828
rect 1986 18788 3056 18816
rect 1986 18785 1998 18788
rect 1940 18779 1998 18785
rect 3050 18776 3056 18788
rect 3108 18776 3114 18828
rect 3510 18816 3516 18828
rect 3471 18788 3516 18816
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 4080 18825 4108 18856
rect 4801 18853 4813 18887
rect 4847 18884 4859 18887
rect 6822 18884 6828 18896
rect 4847 18856 6828 18884
rect 4847 18853 4859 18856
rect 4801 18847 4859 18853
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 9122 18844 9128 18896
rect 9180 18884 9186 18896
rect 9401 18887 9459 18893
rect 9401 18884 9413 18887
rect 9180 18856 9413 18884
rect 9180 18844 9186 18856
rect 9401 18853 9413 18856
rect 9447 18884 9459 18887
rect 9674 18884 9680 18896
rect 9447 18856 9680 18884
rect 9447 18853 9459 18856
rect 9401 18847 9459 18853
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 5626 18816 5632 18828
rect 5587 18788 5632 18816
rect 4065 18779 4123 18785
rect 5626 18776 5632 18788
rect 5684 18776 5690 18828
rect 6086 18816 6092 18828
rect 6047 18788 6092 18816
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8018 18816 8024 18828
rect 6963 18788 8024 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18816 8171 18819
rect 9214 18816 9220 18828
rect 8159 18788 9220 18816
rect 8159 18785 8171 18788
rect 8113 18779 8171 18785
rect 9214 18776 9220 18788
rect 9272 18816 9278 18828
rect 9490 18816 9496 18828
rect 9272 18788 9496 18816
rect 9272 18776 9278 18788
rect 9490 18776 9496 18788
rect 9548 18776 9554 18828
rect 9600 18816 9628 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 12526 18884 12532 18896
rect 11624 18856 12532 18884
rect 10413 18819 10471 18825
rect 9600 18788 10042 18816
rect 10014 18760 10042 18788
rect 10413 18785 10425 18819
rect 10459 18816 10471 18819
rect 11514 18816 11520 18828
rect 10459 18788 11520 18816
rect 10459 18785 10471 18788
rect 10413 18779 10471 18785
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 11624 18825 11652 18856
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 13004 18884 13032 18912
rect 13326 18887 13384 18893
rect 13326 18884 13338 18887
rect 13004 18856 13338 18884
rect 13326 18853 13338 18856
rect 13372 18853 13384 18887
rect 13326 18847 13384 18853
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 19996 18884 20024 18912
rect 14056 18856 16160 18884
rect 14056 18844 14062 18856
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 11876 18819 11934 18825
rect 11876 18785 11888 18819
rect 11922 18816 11934 18819
rect 14274 18816 14280 18828
rect 11922 18788 14280 18816
rect 11922 18785 11934 18788
rect 11876 18779 11934 18785
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14550 18816 14556 18828
rect 14511 18788 14556 18816
rect 14550 18776 14556 18788
rect 14608 18776 14614 18828
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 16132 18825 16160 18856
rect 18156 18856 20024 18884
rect 15749 18819 15807 18825
rect 15749 18816 15761 18819
rect 15528 18788 15761 18816
rect 15528 18776 15534 18788
rect 15749 18785 15761 18788
rect 15795 18785 15807 18819
rect 15749 18779 15807 18785
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18785 16175 18819
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 16117 18779 16175 18785
rect 16224 18788 16589 18816
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18717 3663 18751
rect 3605 18711 3663 18717
rect 3620 18680 3648 18711
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 5077 18751 5135 18757
rect 3752 18720 5028 18748
rect 3752 18708 3758 18720
rect 4246 18680 4252 18692
rect 3620 18652 4252 18680
rect 4246 18640 4252 18652
rect 4304 18640 4310 18692
rect 5000 18680 5028 18720
rect 5077 18717 5089 18751
rect 5123 18748 5135 18751
rect 5534 18748 5540 18760
rect 5123 18720 5540 18748
rect 5123 18717 5135 18720
rect 5077 18711 5135 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5718 18748 5724 18760
rect 5679 18720 5724 18748
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 5813 18751 5871 18757
rect 5813 18717 5825 18751
rect 5859 18717 5871 18751
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 5813 18711 5871 18717
rect 5828 18680 5856 18711
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 5000 18652 5856 18680
rect 6273 18683 6331 18689
rect 6273 18649 6285 18683
rect 6319 18680 6331 18683
rect 7190 18680 7196 18692
rect 6319 18652 7196 18680
rect 6319 18649 6331 18652
rect 6273 18643 6331 18649
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 6178 18612 6184 18624
rect 4479 18584 6184 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 6178 18572 6184 18584
rect 6236 18572 6242 18624
rect 7392 18612 7420 18711
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 7700 18751 7758 18757
rect 7700 18748 7712 18751
rect 7616 18720 7712 18748
rect 7616 18708 7622 18720
rect 7700 18717 7712 18720
rect 7746 18717 7758 18751
rect 7700 18711 7758 18717
rect 7883 18751 7941 18757
rect 7883 18717 7895 18751
rect 7929 18748 7941 18751
rect 9582 18748 9588 18760
rect 7929 18720 9588 18748
rect 7929 18717 7941 18720
rect 7883 18711 7941 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 10014 18757 10048 18760
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 10000 18751 10048 18757
rect 10000 18717 10012 18751
rect 10046 18717 10048 18751
rect 10000 18711 10048 18717
rect 8754 18640 8760 18692
rect 8812 18680 8818 18692
rect 9692 18680 9720 18711
rect 10042 18708 10048 18711
rect 10100 18708 10106 18760
rect 10183 18751 10241 18757
rect 10183 18717 10195 18751
rect 10229 18748 10241 18751
rect 10778 18748 10784 18760
rect 10229 18720 10784 18748
rect 10229 18717 10241 18720
rect 10183 18711 10241 18717
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 13078 18748 13084 18760
rect 13039 18720 13084 18748
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 15930 18748 15936 18760
rect 15891 18720 15936 18748
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 8812 18652 9720 18680
rect 14737 18683 14795 18689
rect 8812 18640 8818 18652
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 15194 18680 15200 18692
rect 14783 18652 15200 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 16224 18680 16252 18788
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 17310 18816 17316 18828
rect 17223 18788 17316 18816
rect 16577 18779 16635 18785
rect 17310 18776 17316 18788
rect 17368 18816 17374 18828
rect 18156 18816 18184 18856
rect 21082 18844 21088 18896
rect 21140 18893 21146 18896
rect 21140 18887 21204 18893
rect 21140 18853 21158 18887
rect 21192 18884 21204 18887
rect 22833 18887 22891 18893
rect 22833 18884 22845 18887
rect 21192 18856 22845 18884
rect 21192 18853 21204 18856
rect 21140 18847 21204 18853
rect 22833 18853 22845 18856
rect 22879 18853 22891 18887
rect 22833 18847 22891 18853
rect 21140 18844 21146 18847
rect 18966 18816 18972 18828
rect 17368 18788 18184 18816
rect 18927 18788 18972 18816
rect 17368 18776 17374 18788
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19236 18819 19294 18825
rect 19236 18785 19248 18819
rect 19282 18816 19294 18819
rect 19978 18816 19984 18828
rect 19282 18788 19984 18816
rect 19282 18785 19294 18788
rect 19236 18779 19294 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20990 18816 20996 18828
rect 20487 18788 20996 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 16298 18708 16304 18760
rect 16356 18708 16362 18760
rect 16850 18708 16856 18760
rect 16908 18757 16914 18760
rect 17126 18757 17132 18760
rect 16908 18751 16958 18757
rect 16908 18717 16912 18751
rect 16946 18717 16958 18751
rect 16908 18711 16958 18717
rect 17083 18751 17132 18757
rect 17083 18717 17095 18751
rect 17129 18717 17132 18751
rect 17083 18711 17132 18717
rect 16908 18708 16914 18711
rect 17126 18708 17132 18711
rect 17184 18708 17190 18760
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22520 18720 22937 18748
rect 22520 18708 22526 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 15620 18652 16252 18680
rect 15620 18640 15626 18652
rect 7650 18612 7656 18624
rect 7392 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18612 7714 18624
rect 8772 18612 8800 18640
rect 7708 18584 8800 18612
rect 7708 18572 7714 18584
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 11790 18612 11796 18624
rect 9456 18584 11796 18612
rect 9456 18572 9462 18584
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 12768 18584 14473 18612
rect 12768 18572 12774 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 15102 18612 15108 18624
rect 15063 18584 15108 18612
rect 14461 18575 14519 18581
rect 15102 18572 15108 18584
rect 15160 18572 15166 18624
rect 16316 18621 16344 18708
rect 22370 18680 22376 18692
rect 22331 18652 22376 18680
rect 22370 18640 22376 18652
rect 22428 18640 22434 18692
rect 16301 18615 16359 18621
rect 16301 18581 16313 18615
rect 16347 18581 16359 18615
rect 18414 18612 18420 18624
rect 18375 18584 18420 18612
rect 16301 18575 16359 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18612 20683 18615
rect 22738 18612 22744 18624
rect 20671 18584 22744 18612
rect 20671 18581 20683 18584
rect 20625 18575 20683 18581
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 1104 18522 23460 18544
rect 1104 18470 4714 18522
rect 4766 18470 4778 18522
rect 4830 18470 4842 18522
rect 4894 18470 4906 18522
rect 4958 18470 12178 18522
rect 12230 18470 12242 18522
rect 12294 18470 12306 18522
rect 12358 18470 12370 18522
rect 12422 18470 19642 18522
rect 19694 18470 19706 18522
rect 19758 18470 19770 18522
rect 19822 18470 19834 18522
rect 19886 18470 23460 18522
rect 1104 18448 23460 18470
rect 3050 18368 3056 18420
rect 3108 18408 3114 18420
rect 3145 18411 3203 18417
rect 3145 18408 3157 18411
rect 3108 18380 3157 18408
rect 3108 18368 3114 18380
rect 3145 18377 3157 18380
rect 3191 18377 3203 18411
rect 3510 18408 3516 18420
rect 3145 18371 3203 18377
rect 3252 18380 3516 18408
rect 3252 18272 3280 18380
rect 3510 18368 3516 18380
rect 3568 18408 3574 18420
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 3568 18380 4629 18408
rect 3568 18368 3574 18380
rect 4617 18377 4629 18380
rect 4663 18377 4675 18411
rect 4617 18371 4675 18377
rect 5166 18368 5172 18420
rect 5224 18408 5230 18420
rect 6457 18411 6515 18417
rect 6457 18408 6469 18411
rect 5224 18380 6469 18408
rect 5224 18368 5230 18380
rect 6457 18377 6469 18380
rect 6503 18377 6515 18411
rect 10778 18408 10784 18420
rect 6457 18371 6515 18377
rect 6840 18380 10272 18408
rect 10739 18380 10784 18408
rect 6840 18340 6868 18380
rect 3160 18244 3280 18272
rect 6104 18312 6868 18340
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2032 18207 2090 18213
rect 2032 18173 2044 18207
rect 2078 18204 2090 18207
rect 3160 18204 3188 18244
rect 2078 18176 3188 18204
rect 3237 18207 3295 18213
rect 2078 18173 2090 18176
rect 2032 18167 2090 18173
rect 3237 18173 3249 18207
rect 3283 18204 3295 18207
rect 3878 18204 3884 18216
rect 3283 18176 3884 18204
rect 3283 18173 3295 18176
rect 3237 18167 3295 18173
rect 3878 18164 3884 18176
rect 3936 18204 3942 18216
rect 4801 18207 4859 18213
rect 4801 18204 4813 18207
rect 3936 18176 4813 18204
rect 3936 18164 3942 18176
rect 4801 18173 4813 18176
rect 4847 18173 4859 18207
rect 4801 18167 4859 18173
rect 5068 18207 5126 18213
rect 5068 18173 5080 18207
rect 5114 18204 5126 18207
rect 6104 18204 6132 18312
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 8076 18244 8309 18272
rect 8076 18232 8082 18244
rect 8297 18241 8309 18244
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8619 18244 9260 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 5114 18176 6132 18204
rect 5114 18173 5126 18176
rect 5068 18167 5126 18173
rect 3504 18139 3562 18145
rect 3504 18105 3516 18139
rect 3550 18136 3562 18139
rect 4246 18136 4252 18148
rect 3550 18108 4252 18136
rect 3550 18105 3562 18108
rect 3504 18099 3562 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 4816 18136 4844 18167
rect 6178 18164 6184 18216
rect 6236 18204 6242 18216
rect 7098 18213 7104 18216
rect 6273 18207 6331 18213
rect 6273 18204 6285 18207
rect 6236 18176 6285 18204
rect 6236 18164 6242 18176
rect 6273 18173 6285 18176
rect 6319 18173 6331 18207
rect 6273 18167 6331 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 7092 18204 7104 18213
rect 7059 18176 7104 18204
rect 6825 18167 6883 18173
rect 7092 18167 7104 18176
rect 6840 18136 6868 18167
rect 7098 18164 7104 18167
rect 7156 18164 7162 18216
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8812 18176 8861 18204
rect 8812 18164 8818 18176
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 9232 18204 9260 18244
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 10042 18272 10048 18284
rect 9364 18244 9409 18272
rect 9508 18244 10048 18272
rect 9364 18232 9370 18244
rect 9508 18204 9536 18244
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 10244 18272 10272 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 11609 18411 11667 18417
rect 11609 18408 11621 18411
rect 11020 18380 11621 18408
rect 11020 18368 11026 18380
rect 11609 18377 11621 18380
rect 11655 18408 11667 18411
rect 12253 18411 12311 18417
rect 12253 18408 12265 18411
rect 11655 18380 12265 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 12253 18377 12265 18380
rect 12299 18377 12311 18411
rect 12253 18371 12311 18377
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 14550 18408 14556 18420
rect 12483 18380 14556 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 16301 18411 16359 18417
rect 16301 18408 16313 18411
rect 15344 18380 16313 18408
rect 15344 18368 15350 18380
rect 16301 18377 16313 18380
rect 16347 18377 16359 18411
rect 16301 18371 16359 18377
rect 10686 18300 10692 18352
rect 10744 18340 10750 18352
rect 10980 18340 11008 18368
rect 11422 18340 11428 18352
rect 10744 18312 11008 18340
rect 11072 18312 11428 18340
rect 10744 18300 10750 18312
rect 11072 18272 11100 18312
rect 11238 18272 11244 18284
rect 10244 18244 11100 18272
rect 11199 18244 11244 18272
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 11348 18281 11376 18312
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 16316 18272 16344 18371
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 17773 18411 17831 18417
rect 17773 18408 17785 18411
rect 16448 18380 17785 18408
rect 16448 18368 16454 18380
rect 17773 18377 17785 18380
rect 17819 18377 17831 18411
rect 18966 18408 18972 18420
rect 17773 18371 17831 18377
rect 18616 18380 18972 18408
rect 13127 18244 13400 18272
rect 16316 18244 16528 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 9232 18176 9536 18204
rect 9585 18207 9643 18213
rect 8849 18167 8907 18173
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 9950 18204 9956 18216
rect 9631 18176 9956 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 11146 18204 11152 18216
rect 11107 18176 11152 18204
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 11790 18204 11796 18216
rect 11751 18176 11796 18204
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 13262 18204 13268 18216
rect 13223 18176 13268 18204
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13372 18204 13400 18244
rect 14366 18204 14372 18216
rect 13372 18176 14372 18204
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15010 18204 15016 18216
rect 14967 18176 15016 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 16390 18204 16396 18216
rect 16351 18176 16396 18204
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16500 18204 16528 18244
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 18616 18281 18644 18380
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19978 18408 19984 18420
rect 19939 18380 19984 18408
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 20128 18380 20173 18408
rect 20128 18368 20134 18380
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 22370 18408 22376 18420
rect 20680 18380 22376 18408
rect 20680 18368 20686 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18104 18244 18613 18272
rect 18104 18232 18110 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 19996 18272 20024 18368
rect 20438 18300 20444 18352
rect 20496 18340 20502 18352
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 20496 18312 20944 18340
rect 20496 18300 20502 18312
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 19996 18244 20545 18272
rect 18601 18235 18659 18241
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 20680 18244 20725 18272
rect 20680 18232 20686 18244
rect 16649 18207 16707 18213
rect 16649 18204 16661 18207
rect 16500 18176 16661 18204
rect 16649 18173 16661 18176
rect 16695 18173 16707 18207
rect 16649 18167 16707 18173
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20916 18213 20944 18312
rect 22388 18312 23029 18340
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 20404 18176 20453 18204
rect 20404 18164 20410 18176
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21361 18207 21419 18213
rect 21361 18173 21373 18207
rect 21407 18204 21419 18207
rect 21450 18204 21456 18216
rect 21407 18176 21456 18204
rect 21407 18173 21419 18176
rect 21361 18167 21419 18173
rect 4816 18108 6868 18136
rect 6288 18080 6316 18108
rect 7558 18096 7564 18148
rect 7616 18136 7622 18148
rect 8018 18136 8024 18148
rect 7616 18108 8024 18136
rect 7616 18096 7622 18108
rect 8018 18096 8024 18108
rect 8076 18136 8082 18148
rect 12805 18139 12863 18145
rect 8076 18108 8340 18136
rect 8076 18096 8082 18108
rect 6178 18068 6184 18080
rect 6139 18040 6184 18068
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6270 18028 6276 18080
rect 6328 18028 6334 18080
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8312 18068 8340 18108
rect 12805 18105 12817 18139
rect 12851 18136 12863 18139
rect 13532 18139 13590 18145
rect 12851 18108 13492 18136
rect 12851 18105 12863 18108
rect 12805 18099 12863 18105
rect 9122 18068 9128 18080
rect 8312 18040 9128 18068
rect 9122 18028 9128 18040
rect 9180 18068 9186 18080
rect 9315 18071 9373 18077
rect 9315 18068 9327 18071
rect 9180 18040 9327 18068
rect 9180 18028 9186 18040
rect 9315 18037 9327 18040
rect 9361 18037 9373 18071
rect 9315 18031 9373 18037
rect 9490 18028 9496 18080
rect 9548 18068 9554 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 9548 18040 10701 18068
rect 9548 18028 9554 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 10689 18031 10747 18037
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 12526 18068 12532 18080
rect 12299 18040 12532 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13464 18068 13492 18108
rect 13532 18105 13544 18139
rect 13578 18136 13590 18139
rect 13998 18136 14004 18148
rect 13578 18108 14004 18136
rect 13578 18105 13590 18108
rect 13532 18099 13590 18105
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 15188 18139 15246 18145
rect 15188 18105 15200 18139
rect 15234 18136 15246 18139
rect 15654 18136 15660 18148
rect 15234 18108 15660 18136
rect 15234 18105 15246 18108
rect 15188 18099 15246 18105
rect 15654 18096 15660 18108
rect 15712 18136 15718 18148
rect 18868 18139 18926 18145
rect 15712 18108 16712 18136
rect 15712 18096 15718 18108
rect 16684 18080 16712 18108
rect 18868 18105 18880 18139
rect 18914 18136 18926 18139
rect 19518 18136 19524 18148
rect 18914 18108 19524 18136
rect 18914 18105 18926 18108
rect 18868 18099 18926 18105
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21376 18136 21404 18167
rect 21450 18164 21456 18176
rect 21508 18164 21514 18216
rect 21634 18213 21640 18216
rect 21628 18204 21640 18213
rect 21595 18176 21640 18204
rect 21628 18167 21640 18176
rect 21634 18164 21640 18167
rect 21692 18164 21698 18216
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22388 18204 22416 18312
rect 23017 18309 23029 18312
rect 23063 18309 23075 18343
rect 23017 18303 23075 18309
rect 21968 18176 22416 18204
rect 22833 18207 22891 18213
rect 21968 18164 21974 18176
rect 22833 18173 22845 18207
rect 22879 18204 22891 18207
rect 23106 18204 23112 18216
rect 22879 18176 23112 18204
rect 22879 18173 22891 18176
rect 22833 18167 22891 18173
rect 23106 18164 23112 18176
rect 23164 18164 23170 18216
rect 22462 18136 22468 18148
rect 20864 18108 21404 18136
rect 21744 18108 22468 18136
rect 20864 18096 20870 18108
rect 14090 18068 14096 18080
rect 12952 18040 12997 18068
rect 13464 18040 14096 18068
rect 12952 18028 12958 18040
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14516 18040 14657 18068
rect 14516 18028 14522 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 14645 18031 14703 18037
rect 16666 18028 16672 18080
rect 16724 18028 16730 18080
rect 21085 18071 21143 18077
rect 21085 18037 21097 18071
rect 21131 18068 21143 18071
rect 21744 18068 21772 18108
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 21131 18040 21772 18068
rect 21131 18037 21143 18040
rect 21085 18031 21143 18037
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 22741 18071 22799 18077
rect 22741 18068 22753 18071
rect 21876 18040 22753 18068
rect 21876 18028 21882 18040
rect 22741 18037 22753 18040
rect 22787 18037 22799 18071
rect 22741 18031 22799 18037
rect 1104 17978 23460 18000
rect 1104 17926 8446 17978
rect 8498 17926 8510 17978
rect 8562 17926 8574 17978
rect 8626 17926 8638 17978
rect 8690 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 23460 17978
rect 1104 17904 23460 17926
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 8941 17867 8999 17873
rect 8941 17864 8953 17867
rect 7800 17836 8953 17864
rect 7800 17824 7806 17836
rect 8941 17833 8953 17836
rect 8987 17833 8999 17867
rect 8941 17827 8999 17833
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 9640 17836 9689 17864
rect 9640 17824 9646 17836
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 10042 17864 10048 17876
rect 10003 17836 10048 17864
rect 9677 17827 9735 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 11793 17867 11851 17873
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 12894 17864 12900 17876
rect 11839 17836 12900 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 13998 17864 14004 17876
rect 13959 17836 14004 17864
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14090 17824 14096 17876
rect 14148 17864 14154 17876
rect 14458 17864 14464 17876
rect 14148 17836 14193 17864
rect 14419 17836 14464 17864
rect 14148 17824 14154 17836
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15010 17864 15016 17876
rect 14967 17836 15016 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 16666 17864 16672 17876
rect 16627 17836 16672 17864
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17497 17867 17555 17873
rect 17497 17864 17509 17867
rect 17184 17836 17509 17864
rect 17184 17824 17190 17836
rect 17497 17833 17509 17836
rect 17543 17833 17555 17867
rect 19426 17864 19432 17876
rect 19387 17836 19432 17864
rect 17497 17827 17555 17833
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 19576 17836 19809 17864
rect 19576 17824 19582 17836
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 21726 17864 21732 17876
rect 19797 17827 19855 17833
rect 21284 17836 21732 17864
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 3234 17796 3240 17808
rect 1820 17768 3240 17796
rect 1820 17756 1826 17768
rect 2148 17737 2176 17768
rect 3234 17756 3240 17768
rect 3292 17796 3298 17808
rect 3878 17796 3884 17808
rect 3292 17768 3884 17796
rect 3292 17756 3298 17768
rect 3878 17756 3884 17768
rect 3936 17796 3942 17808
rect 4614 17796 4620 17808
rect 3936 17768 4620 17796
rect 3936 17756 3942 17768
rect 4614 17756 4620 17768
rect 4672 17796 4678 17808
rect 5068 17799 5126 17805
rect 4672 17768 4844 17796
rect 4672 17756 4678 17768
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17697 2191 17731
rect 2133 17691 2191 17697
rect 2400 17731 2458 17737
rect 2400 17697 2412 17731
rect 2446 17728 2458 17731
rect 3326 17728 3332 17740
rect 2446 17700 3332 17728
rect 2446 17697 2458 17700
rect 2400 17691 2458 17697
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 4816 17737 4844 17768
rect 5068 17765 5080 17799
rect 5114 17796 5126 17799
rect 5718 17796 5724 17808
rect 5114 17768 5724 17796
rect 5114 17765 5126 17768
rect 5068 17759 5126 17765
rect 5718 17756 5724 17768
rect 5776 17796 5782 17808
rect 6178 17796 6184 17808
rect 5776 17768 6184 17796
rect 5776 17756 5782 17768
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 8570 17756 8576 17808
rect 8628 17796 8634 17808
rect 8849 17799 8907 17805
rect 8849 17796 8861 17799
rect 8628 17768 8861 17796
rect 8628 17756 8634 17768
rect 8849 17765 8861 17768
rect 8895 17765 8907 17799
rect 8849 17759 8907 17765
rect 9030 17756 9036 17808
rect 9088 17796 9094 17808
rect 10137 17799 10195 17805
rect 10137 17796 10149 17799
rect 9088 17768 10149 17796
rect 9088 17756 9094 17768
rect 10137 17765 10149 17768
rect 10183 17765 10195 17799
rect 10137 17759 10195 17765
rect 12066 17756 12072 17808
rect 12124 17796 12130 17808
rect 12253 17799 12311 17805
rect 12253 17796 12265 17799
rect 12124 17768 12265 17796
rect 12124 17756 12130 17768
rect 12253 17765 12265 17768
rect 12299 17765 12311 17799
rect 14016 17796 14044 17824
rect 14553 17799 14611 17805
rect 14553 17796 14565 17799
rect 12253 17759 12311 17765
rect 12406 17768 12931 17796
rect 14016 17768 14565 17796
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17697 4859 17731
rect 4801 17691 4859 17697
rect 7276 17731 7334 17737
rect 7276 17697 7288 17731
rect 7322 17728 7334 17731
rect 7322 17700 8248 17728
rect 7322 17697 7334 17700
rect 7276 17691 7334 17697
rect 8220 17672 8248 17700
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9180 17700 9505 17728
rect 9180 17688 9186 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10873 17731 10931 17737
rect 10873 17728 10885 17731
rect 9732 17700 10885 17728
rect 9732 17688 9738 17700
rect 10873 17697 10885 17700
rect 10919 17697 10931 17731
rect 10873 17691 10931 17697
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 12406 17728 12434 17768
rect 12903 17737 12931 17768
rect 14553 17765 14565 17768
rect 14599 17765 14611 17799
rect 15028 17796 15056 17824
rect 15028 17768 15332 17796
rect 14553 17759 14611 17765
rect 15304 17740 15332 17768
rect 15470 17756 15476 17808
rect 15528 17805 15534 17808
rect 15528 17799 15592 17805
rect 15528 17765 15546 17799
rect 15580 17765 15592 17799
rect 15528 17759 15592 17765
rect 17589 17799 17647 17805
rect 17589 17765 17601 17799
rect 17635 17796 17647 17799
rect 18414 17796 18420 17808
rect 17635 17768 18420 17796
rect 17635 17765 17647 17768
rect 17589 17759 17647 17765
rect 15528 17756 15534 17759
rect 18414 17756 18420 17768
rect 18472 17756 18478 17808
rect 20993 17799 21051 17805
rect 20993 17765 21005 17799
rect 21039 17796 21051 17799
rect 21085 17799 21143 17805
rect 21085 17796 21097 17799
rect 21039 17768 21097 17796
rect 21039 17765 21051 17768
rect 20993 17759 21051 17765
rect 21085 17765 21097 17768
rect 21131 17796 21143 17799
rect 21174 17796 21180 17808
rect 21131 17768 21180 17796
rect 21131 17765 21143 17768
rect 21085 17759 21143 17765
rect 21174 17756 21180 17768
rect 21232 17756 21238 17808
rect 21284 17805 21312 17836
rect 21726 17824 21732 17836
rect 21784 17864 21790 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 21784 17836 22937 17864
rect 21784 17824 21790 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 21818 17805 21824 17808
rect 21269 17799 21327 17805
rect 21269 17765 21281 17799
rect 21315 17765 21327 17799
rect 21812 17796 21824 17805
rect 21779 17768 21824 17796
rect 21269 17759 21327 17765
rect 21812 17759 21824 17768
rect 21818 17756 21824 17759
rect 21876 17756 21882 17808
rect 12207 17700 12434 17728
rect 12888 17731 12946 17737
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 12888 17697 12900 17731
rect 12934 17728 12946 17731
rect 13814 17728 13820 17740
rect 12934 17700 13820 17728
rect 12934 17697 12946 17700
rect 12888 17691 12946 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 15102 17728 15108 17740
rect 15063 17700 15108 17728
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15286 17688 15292 17740
rect 15344 17728 15350 17740
rect 15344 17700 15437 17728
rect 15344 17688 15350 17700
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 16448 17700 17969 17728
rect 16448 17688 16454 17700
rect 17957 17697 17969 17700
rect 18003 17728 18015 17731
rect 18046 17728 18052 17740
rect 18003 17700 18052 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 18224 17731 18282 17737
rect 18224 17697 18236 17731
rect 18270 17728 18282 17731
rect 19426 17728 19432 17740
rect 18270 17700 19432 17728
rect 18270 17697 18282 17700
rect 18224 17691 18282 17697
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 20254 17728 20260 17740
rect 20215 17700 20260 17728
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 3142 17620 3148 17672
rect 3200 17660 3206 17672
rect 3602 17660 3608 17672
rect 3200 17632 3608 17660
rect 3200 17620 3206 17632
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 6972 17632 7021 17660
rect 6972 17620 6978 17632
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7009 17623 7067 17629
rect 8202 17620 8208 17672
rect 8260 17660 8266 17672
rect 9033 17663 9091 17669
rect 9033 17660 9045 17663
rect 8260 17632 9045 17660
rect 8260 17620 8266 17632
rect 9033 17629 9045 17632
rect 9079 17629 9091 17663
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 9033 17623 9091 17629
rect 9140 17632 10241 17660
rect 8481 17595 8539 17601
rect 8481 17561 8493 17595
rect 8527 17592 8539 17595
rect 8938 17592 8944 17604
rect 8527 17564 8944 17592
rect 8527 17561 8539 17564
rect 8481 17555 8539 17561
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 3513 17527 3571 17533
rect 3513 17493 3525 17527
rect 3559 17524 3571 17527
rect 3602 17524 3608 17536
rect 3559 17496 3608 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 6178 17524 6184 17536
rect 6139 17496 6184 17524
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8389 17527 8447 17533
rect 8389 17524 8401 17527
rect 8168 17496 8401 17524
rect 8168 17484 8174 17496
rect 8389 17493 8401 17496
rect 8435 17524 8447 17527
rect 9140 17524 9168 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10962 17660 10968 17672
rect 10923 17632 10968 17660
rect 10229 17623 10287 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 11054 17620 11060 17672
rect 11112 17660 11118 17672
rect 11112 17632 11157 17660
rect 11112 17620 11118 17632
rect 12434 17620 12440 17672
rect 12492 17660 12498 17672
rect 12621 17663 12679 17669
rect 12492 17632 12537 17660
rect 12492 17620 12498 17632
rect 12621 17629 12633 17663
rect 12667 17629 12679 17663
rect 14642 17660 14648 17672
rect 14603 17632 14648 17660
rect 12621 17623 12679 17629
rect 8435 17496 9168 17524
rect 9309 17527 9367 17533
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9398 17524 9404 17536
rect 9355 17496 9404 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 10042 17484 10048 17536
rect 10100 17524 10106 17536
rect 10505 17527 10563 17533
rect 10505 17524 10517 17527
rect 10100 17496 10517 17524
rect 10100 17484 10106 17496
rect 10505 17493 10517 17496
rect 10551 17493 10563 17527
rect 12636 17524 12664 17623
rect 14642 17620 14648 17632
rect 14700 17620 14706 17672
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17660 17831 17663
rect 17862 17660 17868 17672
rect 17819 17632 17868 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17660 20131 17663
rect 20162 17660 20168 17672
rect 20119 17632 20168 17660
rect 20119 17629 20131 17632
rect 20073 17623 20131 17629
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17129 17595 17187 17601
rect 17129 17592 17141 17595
rect 17092 17564 17141 17592
rect 17092 17552 17098 17564
rect 17129 17561 17141 17564
rect 17175 17561 17187 17595
rect 19334 17592 19340 17604
rect 19295 17564 19340 17592
rect 17129 17555 17187 17561
rect 19334 17552 19340 17564
rect 19392 17592 19398 17604
rect 19904 17592 19932 17623
rect 20162 17620 20168 17632
rect 20220 17660 20226 17672
rect 20622 17660 20628 17672
rect 20220 17632 20628 17660
rect 20220 17620 20226 17632
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21508 17632 21557 17660
rect 21508 17620 21514 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 23106 17660 23112 17672
rect 23067 17632 23112 17660
rect 21545 17623 21603 17629
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 19392 17564 19932 17592
rect 19392 17552 19398 17564
rect 13262 17524 13268 17536
rect 12636 17496 13268 17524
rect 10505 17487 10563 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 20438 17524 20444 17536
rect 20399 17496 20444 17524
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 21453 17527 21511 17533
rect 21453 17493 21465 17527
rect 21499 17524 21511 17527
rect 22830 17524 22836 17536
rect 21499 17496 22836 17524
rect 21499 17493 21511 17496
rect 21453 17487 21511 17493
rect 22830 17484 22836 17496
rect 22888 17484 22894 17536
rect 1104 17434 23460 17456
rect 1104 17382 4714 17434
rect 4766 17382 4778 17434
rect 4830 17382 4842 17434
rect 4894 17382 4906 17434
rect 4958 17382 12178 17434
rect 12230 17382 12242 17434
rect 12294 17382 12306 17434
rect 12358 17382 12370 17434
rect 12422 17382 19642 17434
rect 19694 17382 19706 17434
rect 19758 17382 19770 17434
rect 19822 17382 19834 17434
rect 19886 17382 23460 17434
rect 1104 17360 23460 17382
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4709 17323 4767 17329
rect 4709 17320 4721 17323
rect 4304 17292 4721 17320
rect 4304 17280 4310 17292
rect 4709 17289 4721 17292
rect 4755 17289 4767 17323
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 4709 17283 4767 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6420 17292 6561 17320
rect 6420 17280 6426 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6822 17320 6828 17332
rect 6783 17292 6828 17320
rect 6549 17283 6607 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 8018 17320 8024 17332
rect 7979 17292 8024 17320
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 9490 17320 9496 17332
rect 8628 17292 9496 17320
rect 8628 17280 8634 17292
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 9585 17323 9643 17329
rect 9585 17289 9597 17323
rect 9631 17320 9643 17323
rect 9766 17320 9772 17332
rect 9631 17292 9772 17320
rect 9631 17289 9643 17292
rect 9585 17283 9643 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 10962 17320 10968 17332
rect 9907 17292 10968 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 12066 17320 12072 17332
rect 12027 17292 12072 17320
rect 12066 17280 12072 17292
rect 12124 17320 12130 17332
rect 12710 17320 12716 17332
rect 12124 17292 12716 17320
rect 12124 17280 12130 17292
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 13814 17320 13820 17332
rect 13775 17292 13820 17320
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 15381 17323 15439 17329
rect 15381 17289 15393 17323
rect 15427 17320 15439 17323
rect 15470 17320 15476 17332
rect 15427 17292 15476 17320
rect 15427 17289 15439 17292
rect 15381 17283 15439 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 19426 17320 19432 17332
rect 19387 17292 19432 17320
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 21545 17323 21603 17329
rect 21545 17320 21557 17323
rect 21416 17292 21557 17320
rect 21416 17280 21422 17292
rect 21545 17289 21557 17292
rect 21591 17289 21603 17323
rect 21545 17283 21603 17289
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 1857 17187 1915 17193
rect 1857 17184 1869 17187
rect 1636 17156 1869 17184
rect 1636 17144 1642 17156
rect 1857 17153 1869 17156
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 3329 17187 3387 17193
rect 3329 17184 3341 17187
rect 3292 17156 3341 17184
rect 3292 17144 3298 17156
rect 3329 17153 3341 17156
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4672 17156 4813 17184
rect 4672 17144 4678 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 3602 17125 3608 17128
rect 3596 17116 3608 17125
rect 3563 17088 3608 17116
rect 3596 17079 3608 17088
rect 3602 17076 3608 17079
rect 3660 17076 3666 17128
rect 2124 17051 2182 17057
rect 2124 17017 2136 17051
rect 2170 17048 2182 17051
rect 3050 17048 3056 17060
rect 2170 17020 3056 17048
rect 2170 17017 2182 17020
rect 2124 17011 2182 17017
rect 3050 17008 3056 17020
rect 3108 17008 3114 17060
rect 4816 17048 4844 17147
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7064 17156 7389 17184
rect 7064 17144 7070 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17184 10563 17187
rect 18046 17184 18052 17196
rect 10551 17156 10824 17184
rect 18007 17156 18052 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 5068 17119 5126 17125
rect 5068 17085 5080 17119
rect 5114 17116 5126 17119
rect 5626 17116 5632 17128
rect 5114 17088 5632 17116
rect 5114 17085 5126 17088
rect 5068 17079 5126 17085
rect 5626 17076 5632 17088
rect 5684 17116 5690 17128
rect 6178 17116 6184 17128
rect 5684 17088 6184 17116
rect 5684 17076 5690 17088
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 6454 17116 6460 17128
rect 6415 17088 6460 17116
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 7650 17116 7656 17128
rect 7611 17088 7656 17116
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 9766 17116 9772 17128
rect 8251 17088 9772 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 10226 17116 10232 17128
rect 9916 17088 10232 17116
rect 9916 17076 9922 17088
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 10686 17116 10692 17128
rect 10647 17088 10692 17116
rect 10686 17076 10692 17088
rect 10744 17076 10750 17128
rect 10796 17116 10824 17156
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 11238 17116 11244 17128
rect 10796 17088 11244 17116
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 12710 17125 12716 17128
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17085 12495 17119
rect 12704 17116 12716 17125
rect 12671 17088 12716 17116
rect 12437 17079 12495 17085
rect 12704 17079 12716 17088
rect 5258 17048 5264 17060
rect 4816 17020 5264 17048
rect 5258 17008 5264 17020
rect 5316 17008 5322 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 6196 17020 7297 17048
rect 6196 16992 6224 17020
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 8294 17048 8300 17060
rect 7285 17011 7343 17017
rect 7852 17020 8300 17048
rect 3237 16983 3295 16989
rect 3237 16949 3249 16983
rect 3283 16980 3295 16983
rect 3418 16980 3424 16992
rect 3283 16952 3424 16980
rect 3283 16949 3295 16952
rect 3237 16943 3295 16949
rect 3418 16940 3424 16952
rect 3476 16940 3482 16992
rect 6178 16980 6184 16992
rect 6091 16952 6184 16980
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 7852 16989 7880 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8472 17051 8530 17057
rect 8472 17017 8484 17051
rect 8518 17048 8530 17051
rect 8938 17048 8944 17060
rect 8518 17020 8944 17048
rect 8518 17017 8530 17020
rect 8472 17011 8530 17017
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 9677 17051 9735 17057
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 10134 17048 10140 17060
rect 9723 17020 10140 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 9876 16992 9904 17020
rect 10134 17008 10140 17020
rect 10192 17048 10198 17060
rect 10956 17051 11014 17057
rect 10192 17020 10548 17048
rect 10192 17008 10198 17020
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6328 16952 7205 16980
rect 6328 16940 6334 16952
rect 7193 16949 7205 16952
rect 7239 16949 7251 16983
rect 7193 16943 7251 16949
rect 7837 16983 7895 16989
rect 7837 16949 7849 16983
rect 7883 16949 7895 16983
rect 7837 16943 7895 16949
rect 9858 16940 9864 16992
rect 9916 16940 9922 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10520 16980 10548 17020
rect 10956 17017 10968 17051
rect 11002 17048 11014 17051
rect 11054 17048 11060 17060
rect 11002 17020 11060 17048
rect 11002 17017 11014 17020
rect 10956 17011 11014 17017
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 12452 17048 12480 17079
rect 12710 17076 12716 17079
rect 12768 17076 12774 17128
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13538 17116 13544 17128
rect 13320 17088 13544 17116
rect 13320 17076 13326 17088
rect 13538 17076 13544 17088
rect 13596 17116 13602 17128
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13596 17088 14013 17116
rect 13596 17076 13602 17088
rect 14001 17085 14013 17088
rect 14047 17116 14059 17119
rect 15286 17116 15292 17128
rect 14047 17088 15292 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 19444 17116 19472 17280
rect 22186 17252 22192 17264
rect 21192 17224 22192 17252
rect 20162 17184 20168 17196
rect 20123 17156 20168 17184
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 21192 17193 21220 17224
rect 22186 17212 22192 17224
rect 22244 17252 22250 17264
rect 22244 17224 22968 17252
rect 22244 17212 22250 17224
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 22097 17187 22155 17193
rect 22097 17153 22109 17187
rect 22143 17184 22155 17187
rect 22370 17184 22376 17196
rect 22143 17156 22376 17184
rect 22143 17153 22155 17156
rect 22097 17147 22155 17153
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 22462 17144 22468 17196
rect 22520 17184 22526 17196
rect 22940 17193 22968 17224
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22520 17156 22845 17184
rect 22520 17144 22526 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19444 17088 19901 17116
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 20438 17076 20444 17128
rect 20496 17116 20502 17128
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20496 17088 20913 17116
rect 20496 17076 20502 17088
rect 20901 17085 20913 17088
rect 20947 17085 20959 17119
rect 20901 17079 20959 17085
rect 21818 17076 21824 17128
rect 21876 17116 21882 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21876 17088 21925 17116
rect 21876 17076 21882 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 22738 17116 22744 17128
rect 22699 17088 22744 17116
rect 21913 17079 21971 17085
rect 22738 17076 22744 17088
rect 22796 17076 22802 17128
rect 12526 17048 12532 17060
rect 12452 17020 12532 17048
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 14268 17051 14326 17057
rect 14268 17017 14280 17051
rect 14314 17048 14326 17051
rect 14458 17048 14464 17060
rect 14314 17020 14464 17048
rect 14314 17017 14326 17020
rect 14268 17011 14326 17017
rect 14458 17008 14464 17020
rect 14516 17008 14522 17060
rect 18316 17051 18374 17057
rect 18316 17017 18328 17051
rect 18362 17048 18374 17051
rect 19058 17048 19064 17060
rect 18362 17020 19064 17048
rect 18362 17017 18374 17020
rect 18316 17011 18374 17017
rect 19058 17008 19064 17020
rect 19116 17048 19122 17060
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 19116 17020 19993 17048
rect 19116 17008 19122 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 21542 17048 21548 17060
rect 19981 17011 20039 17017
rect 20548 17020 21548 17048
rect 12710 16980 12716 16992
rect 10376 16952 10421 16980
rect 10520 16952 12716 16980
rect 10376 16940 10382 16952
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 19521 16983 19579 16989
rect 19521 16949 19533 16983
rect 19567 16980 19579 16983
rect 19702 16980 19708 16992
rect 19567 16952 19708 16980
rect 19567 16949 19579 16952
rect 19521 16943 19579 16949
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 20548 16989 20576 17020
rect 21542 17008 21548 17020
rect 21600 17008 21606 17060
rect 21634 17008 21640 17060
rect 21692 17048 21698 17060
rect 22005 17051 22063 17057
rect 22005 17048 22017 17051
rect 21692 17020 22017 17048
rect 21692 17008 21698 17020
rect 22005 17017 22017 17020
rect 22051 17017 22063 17051
rect 22005 17011 22063 17017
rect 20533 16983 20591 16989
rect 20533 16949 20545 16983
rect 20579 16949 20591 16983
rect 20990 16980 20996 16992
rect 20951 16952 20996 16980
rect 20533 16943 20591 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 22370 16980 22376 16992
rect 22331 16952 22376 16980
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 1104 16890 23460 16912
rect 1104 16838 8446 16890
rect 8498 16838 8510 16890
rect 8562 16838 8574 16890
rect 8626 16838 8638 16890
rect 8690 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 23460 16890
rect 1104 16816 23460 16838
rect 3050 16776 3056 16788
rect 3011 16748 3056 16776
rect 3050 16736 3056 16748
rect 3108 16776 3114 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 3108 16748 3617 16776
rect 3108 16736 3114 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 3605 16739 3663 16745
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4120 16748 4445 16776
rect 4120 16736 4126 16748
rect 4433 16745 4445 16748
rect 4479 16776 4491 16779
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4479 16748 4537 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 6454 16776 6460 16788
rect 4764 16748 6460 16776
rect 4764 16736 4770 16748
rect 6454 16736 6460 16748
rect 6512 16736 6518 16788
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 8260 16748 9413 16776
rect 8260 16736 8266 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 9401 16739 9459 16745
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11149 16779 11207 16785
rect 11149 16776 11161 16779
rect 11112 16748 11161 16776
rect 11112 16736 11118 16748
rect 11149 16745 11161 16748
rect 11195 16745 11207 16779
rect 11149 16739 11207 16745
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 14921 16779 14979 16785
rect 14921 16776 14933 16779
rect 11296 16748 14933 16776
rect 11296 16736 11302 16748
rect 14921 16745 14933 16748
rect 14967 16745 14979 16779
rect 14921 16739 14979 16745
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16745 15347 16779
rect 15289 16739 15347 16745
rect 17405 16779 17463 16785
rect 17405 16745 17417 16779
rect 17451 16776 17463 16779
rect 19058 16776 19064 16788
rect 17451 16748 17724 16776
rect 19019 16748 19064 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 1940 16711 1998 16717
rect 1940 16677 1952 16711
rect 1986 16708 1998 16711
rect 2682 16708 2688 16720
rect 1986 16680 2688 16708
rect 1986 16677 1998 16680
rect 1940 16671 1998 16677
rect 2682 16668 2688 16680
rect 2740 16668 2746 16720
rect 5068 16711 5126 16717
rect 5068 16677 5080 16711
rect 5114 16708 5126 16711
rect 6178 16708 6184 16720
rect 5114 16680 6184 16708
rect 5114 16677 5126 16680
rect 5068 16671 5126 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 8846 16708 8852 16720
rect 8404 16680 8852 16708
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1636 16612 1685 16640
rect 1636 16600 1642 16612
rect 1673 16609 1685 16612
rect 1719 16609 1731 16643
rect 1673 16603 1731 16609
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 3510 16640 3516 16652
rect 3471 16612 3516 16640
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4479 16612 4660 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 3160 16513 3188 16600
rect 3694 16532 3700 16584
rect 3752 16572 3758 16584
rect 4632 16572 4660 16612
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 6273 16643 6331 16649
rect 4764 16612 4809 16640
rect 4764 16600 4770 16612
rect 6273 16609 6285 16643
rect 6319 16640 6331 16643
rect 6362 16640 6368 16652
rect 6319 16612 6368 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 7190 16649 7196 16652
rect 7184 16603 7196 16649
rect 7248 16640 7254 16652
rect 7248 16612 7284 16640
rect 7190 16600 7196 16603
rect 7248 16600 7254 16612
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 3752 16544 3797 16572
rect 4632 16544 4813 16572
rect 3752 16532 3758 16544
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 6914 16572 6920 16584
rect 6875 16544 6920 16572
rect 4801 16535 4859 16541
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 3145 16507 3203 16513
rect 3145 16473 3157 16507
rect 3191 16473 3203 16507
rect 6178 16504 6184 16516
rect 6139 16476 6184 16504
rect 3145 16467 3203 16473
rect 6178 16464 6184 16476
rect 6236 16464 6242 16516
rect 8404 16513 8432 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 10036 16711 10094 16717
rect 10036 16677 10048 16711
rect 10082 16708 10094 16711
rect 11256 16708 11284 16736
rect 10082 16680 11284 16708
rect 10082 16677 10094 16680
rect 10036 16671 10094 16677
rect 14090 16668 14096 16720
rect 14148 16708 14154 16720
rect 15102 16708 15108 16720
rect 14148 16680 15108 16708
rect 14148 16668 14154 16680
rect 15102 16668 15108 16680
rect 15160 16708 15166 16720
rect 15304 16708 15332 16739
rect 15160 16680 15332 16708
rect 15924 16711 15982 16717
rect 15160 16668 15166 16680
rect 15924 16677 15936 16711
rect 15970 16708 15982 16711
rect 16206 16708 16212 16720
rect 15970 16680 16212 16708
rect 15970 16677 15982 16680
rect 15924 16671 15982 16677
rect 16206 16668 16212 16680
rect 16264 16668 16270 16720
rect 17696 16708 17724 16748
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19153 16779 19211 16785
rect 19153 16745 19165 16779
rect 19199 16776 19211 16779
rect 20441 16779 20499 16785
rect 20441 16776 20453 16779
rect 19199 16748 20453 16776
rect 19199 16745 19211 16748
rect 19153 16739 19211 16745
rect 20441 16745 20453 16748
rect 20487 16745 20499 16779
rect 20441 16739 20499 16745
rect 21361 16779 21419 16785
rect 21361 16745 21373 16779
rect 21407 16776 21419 16779
rect 22462 16776 22468 16788
rect 21407 16748 22468 16776
rect 21407 16745 21419 16748
rect 21361 16739 21419 16745
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 23106 16776 23112 16788
rect 23067 16748 23112 16776
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 18046 16708 18052 16720
rect 17696 16680 18052 16708
rect 8757 16643 8815 16649
rect 8757 16609 8769 16643
rect 8803 16640 8815 16643
rect 9030 16640 9036 16652
rect 8803 16612 9036 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9214 16640 9220 16652
rect 9175 16612 9220 16640
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16640 11759 16643
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 11747 16612 12173 16640
rect 11747 16609 11759 16612
rect 11701 16603 11759 16609
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 13538 16640 13544 16652
rect 13499 16612 13544 16640
rect 12161 16603 12219 16609
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 13808 16643 13866 16649
rect 13808 16609 13820 16643
rect 13854 16640 13866 16643
rect 14182 16640 14188 16652
rect 13854 16612 14188 16640
rect 13854 16609 13866 16612
rect 13808 16603 13866 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16640 15531 16643
rect 17218 16640 17224 16652
rect 15519 16612 17224 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 17586 16640 17592 16652
rect 17547 16612 17592 16640
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 17696 16649 17724 16680
rect 18046 16668 18052 16680
rect 18104 16708 18110 16720
rect 18690 16708 18696 16720
rect 18104 16680 18696 16708
rect 18104 16668 18110 16680
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 19702 16668 19708 16720
rect 19760 16708 19766 16720
rect 20349 16711 20407 16717
rect 20349 16708 20361 16711
rect 19760 16680 20361 16708
rect 19760 16668 19766 16680
rect 20349 16677 20361 16680
rect 20395 16677 20407 16711
rect 20349 16671 20407 16677
rect 21726 16668 21732 16720
rect 21784 16717 21790 16720
rect 21784 16711 21848 16717
rect 21784 16677 21802 16711
rect 21836 16677 21848 16711
rect 21784 16671 21848 16677
rect 21784 16668 21790 16671
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17948 16643 18006 16649
rect 17948 16609 17960 16643
rect 17994 16640 18006 16643
rect 19426 16640 19432 16652
rect 17994 16612 19432 16640
rect 17994 16609 18006 16612
rect 17948 16603 18006 16609
rect 19426 16600 19432 16612
rect 19484 16640 19490 16652
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 19484 16612 19533 16640
rect 19484 16600 19490 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 21174 16640 21180 16652
rect 21135 16612 21180 16640
rect 19521 16603 19579 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21450 16600 21456 16652
rect 21508 16640 21514 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21508 16612 21557 16640
rect 21508 16600 21514 16612
rect 21545 16609 21557 16612
rect 21591 16609 21603 16643
rect 21545 16603 21603 16609
rect 8846 16572 8852 16584
rect 8807 16544 8852 16572
rect 8846 16532 8852 16544
rect 8904 16532 8910 16584
rect 8938 16532 8944 16584
rect 8996 16572 9002 16584
rect 9766 16572 9772 16584
rect 8996 16544 9041 16572
rect 9727 16544 9772 16572
rect 8996 16532 9002 16544
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 11974 16572 11980 16584
rect 11935 16544 11980 16572
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15344 16544 15669 16572
rect 15344 16532 15350 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 19392 16544 19625 16572
rect 19392 16532 19398 16544
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20162 16572 20168 16584
rect 19843 16544 20168 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16572 20683 16575
rect 20671 16544 21036 16572
rect 20671 16541 20683 16544
rect 20625 16535 20683 16541
rect 8389 16507 8447 16513
rect 8389 16473 8401 16507
rect 8435 16473 8447 16507
rect 8389 16467 8447 16473
rect 12529 16507 12587 16513
rect 12529 16473 12541 16507
rect 12575 16504 12587 16507
rect 12710 16504 12716 16516
rect 12575 16476 12716 16504
rect 12575 16473 12587 16476
rect 12529 16467 12587 16473
rect 12710 16464 12716 16476
rect 12768 16504 12774 16516
rect 19981 16507 20039 16513
rect 12768 16476 13308 16504
rect 12768 16464 12774 16476
rect 5810 16396 5816 16448
rect 5868 16436 5874 16448
rect 6457 16439 6515 16445
rect 6457 16436 6469 16439
rect 5868 16408 6469 16436
rect 5868 16396 5874 16408
rect 6457 16405 6469 16408
rect 6503 16405 6515 16439
rect 8294 16436 8300 16448
rect 8255 16408 8300 16436
rect 6457 16399 6515 16405
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 11333 16439 11391 16445
rect 11333 16405 11345 16439
rect 11379 16436 11391 16439
rect 11882 16436 11888 16448
rect 11379 16408 11888 16436
rect 11379 16405 11391 16408
rect 11333 16399 11391 16405
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 13280 16436 13308 16476
rect 19981 16473 19993 16507
rect 20027 16504 20039 16507
rect 20254 16504 20260 16516
rect 20027 16476 20260 16504
rect 20027 16473 20039 16476
rect 19981 16467 20039 16473
rect 20254 16464 20260 16476
rect 20312 16464 20318 16516
rect 15194 16436 15200 16448
rect 13280 16408 15200 16436
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 17034 16436 17040 16448
rect 16995 16408 17040 16436
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 20898 16396 20904 16448
rect 20956 16436 20962 16448
rect 21008 16436 21036 16544
rect 21910 16436 21916 16448
rect 20956 16408 21916 16436
rect 20956 16396 20962 16408
rect 21910 16396 21916 16408
rect 21968 16396 21974 16448
rect 22922 16436 22928 16448
rect 22883 16408 22928 16436
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 1104 16346 23460 16368
rect 1104 16294 4714 16346
rect 4766 16294 4778 16346
rect 4830 16294 4842 16346
rect 4894 16294 4906 16346
rect 4958 16294 12178 16346
rect 12230 16294 12242 16346
rect 12294 16294 12306 16346
rect 12358 16294 12370 16346
rect 12422 16294 19642 16346
rect 19694 16294 19706 16346
rect 19758 16294 19770 16346
rect 19822 16294 19834 16346
rect 19886 16294 23460 16346
rect 1104 16272 23460 16294
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3384 16204 3433 16232
rect 3384 16192 3390 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 3421 16195 3479 16201
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 3786 16232 3792 16244
rect 3559 16204 3792 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 3436 16096 3464 16195
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 5537 16235 5595 16241
rect 5537 16201 5549 16235
rect 5583 16232 5595 16235
rect 8018 16232 8024 16244
rect 5583 16204 8024 16232
rect 5583 16201 5595 16204
rect 5537 16195 5595 16201
rect 8018 16192 8024 16204
rect 8076 16192 8082 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8846 16232 8852 16244
rect 8343 16204 8852 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 9306 16232 9312 16244
rect 9267 16204 9312 16232
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 11425 16235 11483 16241
rect 11425 16201 11437 16235
rect 11471 16232 11483 16235
rect 11790 16232 11796 16244
rect 11471 16204 11796 16232
rect 11471 16201 11483 16204
rect 11425 16195 11483 16201
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 13909 16235 13967 16241
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 14918 16232 14924 16244
rect 13955 16204 14924 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17310 16232 17316 16244
rect 17083 16204 17316 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 19426 16232 19432 16244
rect 19387 16204 19432 16232
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 21174 16232 21180 16244
rect 21135 16204 21180 16232
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 22370 16232 22376 16244
rect 21560 16204 22376 16232
rect 3694 16124 3700 16176
rect 3752 16164 3758 16176
rect 4525 16167 4583 16173
rect 3752 16136 4108 16164
rect 3752 16124 3758 16136
rect 4080 16105 4108 16136
rect 4525 16133 4537 16167
rect 4571 16164 4583 16167
rect 8036 16164 8064 16192
rect 11333 16167 11391 16173
rect 4571 16136 5948 16164
rect 8036 16136 9168 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3436 16068 3985 16096
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 5261 16099 5319 16105
rect 5261 16096 5273 16099
rect 4672 16068 5273 16096
rect 4672 16056 4678 16068
rect 5261 16065 5273 16068
rect 5307 16096 5319 16099
rect 5810 16096 5816 16108
rect 5307 16068 5816 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 1670 15988 1676 16040
rect 1728 16028 1734 16040
rect 2038 16028 2044 16040
rect 1728 16000 2044 16028
rect 1728 15988 1734 16000
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2308 16031 2366 16037
rect 2308 15997 2320 16031
rect 2354 16028 2366 16031
rect 3510 16028 3516 16040
rect 2354 16000 3516 16028
rect 2354 15997 2366 16000
rect 2308 15991 2366 15997
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3660 16000 3893 16028
rect 3660 15988 3666 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 16028 4399 16031
rect 4387 16000 4752 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 4724 15901 4752 16000
rect 5074 15988 5080 16040
rect 5132 16028 5138 16040
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 5132 16000 5181 16028
rect 5132 15988 5138 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 5350 15988 5356 16040
rect 5408 16028 5414 16040
rect 5920 16037 5948 16136
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6546 16096 6552 16108
rect 6227 16068 6552 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 6546 16056 6552 16068
rect 6604 16096 6610 16108
rect 6604 16068 6960 16096
rect 6604 16056 6610 16068
rect 5905 16031 5963 16037
rect 5408 16000 5847 16028
rect 5408 15988 5414 16000
rect 5718 15960 5724 15972
rect 5092 15932 5724 15960
rect 5092 15901 5120 15932
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 5819 15960 5847 16000
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 6365 16031 6423 16037
rect 6365 15997 6377 16031
rect 6411 16028 6423 16031
rect 6638 16028 6644 16040
rect 6411 16000 6644 16028
rect 6411 15997 6423 16000
rect 6365 15991 6423 15997
rect 6638 15988 6644 16000
rect 6696 15988 6702 16040
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6932 16028 6960 16068
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 8352 16068 8861 16096
rect 8352 16056 8358 16068
rect 8849 16065 8861 16068
rect 8895 16065 8907 16099
rect 8849 16059 8907 16065
rect 7374 16028 7380 16040
rect 6932 16000 7380 16028
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 8754 16028 8760 16040
rect 8711 16000 8760 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 8754 15988 8760 16000
rect 8812 15988 8818 16040
rect 9140 16037 9168 16136
rect 11333 16133 11345 16167
rect 11379 16164 11391 16167
rect 11379 16136 11928 16164
rect 11379 16133 11391 16136
rect 11333 16127 11391 16133
rect 11900 16108 11928 16136
rect 9858 16105 9864 16108
rect 9816 16099 9864 16105
rect 9816 16065 9828 16099
rect 9862 16065 9864 16099
rect 9816 16059 9864 16065
rect 9858 16056 9864 16059
rect 9916 16056 9922 16108
rect 10042 16105 10048 16108
rect 9999 16099 10048 16105
rect 9999 16065 10011 16099
rect 10045 16065 10048 16099
rect 9999 16059 10048 16065
rect 10042 16056 10048 16059
rect 10100 16056 10106 16108
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 11882 16096 11888 16108
rect 11795 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 12299 16068 12572 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9539 16000 10916 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 5997 15963 6055 15969
rect 5997 15960 6009 15963
rect 5819 15932 6009 15960
rect 5997 15929 6009 15932
rect 6043 15929 6055 15963
rect 5997 15923 6055 15929
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 7070 15963 7128 15969
rect 7070 15960 7082 15963
rect 6972 15932 7082 15960
rect 6972 15920 6978 15932
rect 7070 15929 7082 15932
rect 7116 15929 7128 15963
rect 7070 15923 7128 15929
rect 8386 15920 8392 15972
rect 8444 15960 8450 15972
rect 8444 15932 8800 15960
rect 8444 15920 8450 15932
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15861 4767 15895
rect 4709 15855 4767 15861
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15861 5135 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 5077 15855 5135 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 8772 15901 8800 15932
rect 8846 15920 8852 15972
rect 8904 15960 8910 15972
rect 9508 15960 9536 15991
rect 8904 15932 9536 15960
rect 10888 15960 10916 16000
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11992 16028 12020 16059
rect 12544 16040 12572 16068
rect 14182 16056 14188 16108
rect 14240 16096 14246 16108
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 14240 16068 14473 16096
rect 14240 16056 14246 16068
rect 14461 16065 14473 16068
rect 14507 16096 14519 16099
rect 14550 16096 14556 16108
rect 14507 16068 14556 16096
rect 14507 16065 14519 16068
rect 14461 16059 14519 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 15712 16068 15757 16096
rect 15712 16056 15718 16068
rect 17034 16056 17040 16108
rect 17092 16096 17098 16108
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 17092 16068 17693 16096
rect 17092 16056 17098 16068
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 20162 16096 20168 16108
rect 20123 16068 20168 16096
rect 17681 16059 17739 16065
rect 20162 16056 20168 16068
rect 20220 16056 20226 16108
rect 20898 16096 20904 16108
rect 20859 16068 20904 16096
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 11112 16000 12020 16028
rect 11112 15988 11118 16000
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 12124 16000 12449 16028
rect 12124 15988 12130 16000
rect 12437 15997 12449 16000
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 15197 16031 15255 16037
rect 15197 16028 15209 16031
rect 12584 16000 15209 16028
rect 12584 15988 12590 16000
rect 15197 15997 15209 16000
rect 15243 15997 15255 16031
rect 15197 15991 15255 15997
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15344 16000 15945 16028
rect 15344 15988 15350 16000
rect 15933 15997 15945 16000
rect 15979 16028 15991 16031
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 15979 16000 17509 16028
rect 15979 15997 15991 16000
rect 15933 15991 15991 15997
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 17497 15991 17555 15997
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 20346 16028 20352 16040
rect 18156 16000 20352 16028
rect 10888 15932 11928 15960
rect 8904 15920 8910 15932
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7248 15864 8217 15892
rect 7248 15852 7254 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8757 15895 8815 15901
rect 8757 15861 8769 15895
rect 8803 15861 8815 15895
rect 8757 15855 8815 15861
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 11793 15895 11851 15901
rect 11793 15892 11805 15895
rect 10376 15864 11805 15892
rect 10376 15852 10382 15864
rect 11793 15861 11805 15864
rect 11839 15861 11851 15895
rect 11900 15892 11928 15932
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 12682 15963 12740 15969
rect 12682 15960 12694 15963
rect 12032 15932 12694 15960
rect 12032 15920 12038 15932
rect 12682 15929 12694 15932
rect 12728 15929 12740 15963
rect 12682 15923 12740 15929
rect 14277 15963 14335 15969
rect 14277 15929 14289 15963
rect 14323 15960 14335 15963
rect 14737 15963 14795 15969
rect 14737 15960 14749 15963
rect 14323 15932 14749 15960
rect 14323 15929 14335 15932
rect 14277 15923 14335 15929
rect 14737 15929 14749 15932
rect 14783 15929 14795 15963
rect 17589 15963 17647 15969
rect 14737 15923 14795 15929
rect 16583 15932 17356 15960
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 11900 15864 12265 15892
rect 11793 15855 11851 15861
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 13814 15892 13820 15904
rect 13775 15864 13820 15892
rect 12253 15855 12311 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 14240 15864 14381 15892
rect 14240 15852 14246 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 14369 15855 14427 15861
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15194 15892 15200 15904
rect 15151 15864 15200 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 15663 15895 15721 15901
rect 15663 15892 15675 15895
rect 15252 15864 15675 15892
rect 15252 15852 15258 15864
rect 15663 15861 15675 15864
rect 15709 15892 15721 15895
rect 16583 15892 16611 15932
rect 15709 15864 16611 15892
rect 15709 15861 15721 15864
rect 15663 15855 15721 15861
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 17328 15892 17356 15932
rect 17589 15929 17601 15963
rect 17635 15960 17647 15963
rect 17678 15960 17684 15972
rect 17635 15932 17684 15960
rect 17635 15929 17647 15932
rect 17589 15923 17647 15929
rect 17678 15920 17684 15932
rect 17736 15920 17742 15972
rect 18156 15892 18184 16000
rect 20346 15988 20352 16000
rect 20404 15988 20410 16040
rect 18316 15963 18374 15969
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 19334 15960 19340 15972
rect 18362 15932 19340 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19536 15932 20729 15960
rect 19536 15901 19564 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 21560 15904 21588 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 21634 16056 21640 16108
rect 21692 16096 21698 16108
rect 21821 16099 21879 16105
rect 21692 16068 21737 16096
rect 21692 16056 21698 16068
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 22278 16096 22284 16108
rect 21867 16068 22284 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 22278 16056 22284 16068
rect 22336 16056 22342 16108
rect 22462 16096 22468 16108
rect 22423 16068 22468 16096
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16096 22707 16099
rect 22922 16096 22928 16108
rect 22695 16068 22928 16096
rect 22695 16065 22707 16068
rect 22649 16059 22707 16065
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 21652 16028 21680 16056
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 21652 16000 22845 16028
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 22373 15963 22431 15969
rect 22373 15929 22385 15963
rect 22419 15960 22431 15963
rect 22419 15932 23060 15960
rect 22419 15929 22431 15932
rect 22373 15923 22431 15929
rect 17184 15864 17229 15892
rect 17328 15864 18184 15892
rect 19521 15895 19579 15901
rect 17184 15852 17190 15864
rect 19521 15861 19533 15895
rect 19567 15861 19579 15895
rect 19886 15892 19892 15904
rect 19847 15864 19892 15892
rect 19521 15855 19579 15861
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20349 15895 20407 15901
rect 20036 15864 20081 15892
rect 20036 15852 20042 15864
rect 20349 15861 20361 15895
rect 20395 15892 20407 15895
rect 20438 15892 20444 15904
rect 20395 15864 20444 15892
rect 20395 15861 20407 15864
rect 20349 15855 20407 15861
rect 20438 15852 20444 15864
rect 20496 15852 20502 15904
rect 20806 15892 20812 15904
rect 20767 15864 20812 15892
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 21542 15892 21548 15904
rect 21503 15864 21548 15892
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22186 15892 22192 15904
rect 22051 15864 22192 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23032 15901 23060 15932
rect 23017 15895 23075 15901
rect 23017 15861 23029 15895
rect 23063 15861 23075 15895
rect 23017 15855 23075 15861
rect 1104 15802 23460 15824
rect 1104 15750 8446 15802
rect 8498 15750 8510 15802
rect 8562 15750 8574 15802
rect 8626 15750 8638 15802
rect 8690 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 23460 15802
rect 1104 15728 23460 15750
rect 7466 15688 7472 15700
rect 7116 15660 7472 15688
rect 4522 15620 4528 15632
rect 3896 15592 4528 15620
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 1670 15552 1676 15564
rect 1627 15524 1676 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 1670 15512 1676 15524
rect 1728 15512 1734 15564
rect 1848 15555 1906 15561
rect 1848 15521 1860 15555
rect 1894 15552 1906 15555
rect 3050 15552 3056 15564
rect 1894 15524 3056 15552
rect 1894 15521 1906 15524
rect 1848 15515 1906 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 3418 15552 3424 15564
rect 3379 15524 3424 15552
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3513 15487 3571 15493
rect 3513 15484 3525 15487
rect 3016 15456 3525 15484
rect 3016 15444 3022 15456
rect 3513 15453 3525 15456
rect 3559 15453 3571 15487
rect 3513 15447 3571 15453
rect 3697 15487 3755 15493
rect 3697 15453 3709 15487
rect 3743 15484 3755 15487
rect 3896 15484 3924 15592
rect 4522 15580 4528 15592
rect 4580 15580 4586 15632
rect 7116 15629 7144 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 9030 15688 9036 15700
rect 8991 15660 9036 15688
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9953 15691 10011 15697
rect 9953 15657 9965 15691
rect 9999 15688 10011 15691
rect 10318 15688 10324 15700
rect 9999 15660 10324 15688
rect 9999 15657 10011 15660
rect 9953 15651 10011 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12161 15691 12219 15697
rect 12161 15688 12173 15691
rect 12032 15660 12173 15688
rect 12032 15648 12038 15660
rect 12161 15657 12173 15660
rect 12207 15657 12219 15691
rect 12161 15651 12219 15657
rect 12710 15648 12716 15700
rect 12768 15697 12774 15700
rect 12768 15688 12777 15697
rect 14182 15688 14188 15700
rect 12768 15660 12813 15688
rect 14143 15660 14188 15688
rect 12768 15651 12777 15660
rect 12768 15648 12774 15651
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 14645 15691 14703 15697
rect 14645 15657 14657 15691
rect 14691 15688 14703 15691
rect 15286 15688 15292 15700
rect 14691 15660 15292 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 7101 15623 7159 15629
rect 7101 15589 7113 15623
rect 7147 15589 7159 15623
rect 7101 15583 7159 15589
rect 7190 15580 7196 15632
rect 7248 15620 7254 15632
rect 7285 15623 7343 15629
rect 7285 15620 7297 15623
rect 7248 15592 7297 15620
rect 7248 15580 7254 15592
rect 7285 15589 7297 15592
rect 7331 15589 7343 15623
rect 7285 15583 7343 15589
rect 7828 15623 7886 15629
rect 7828 15589 7840 15623
rect 7874 15620 7886 15623
rect 8294 15620 8300 15632
rect 7874 15592 8300 15620
rect 7874 15589 7886 15592
rect 7828 15583 7886 15589
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 10413 15623 10471 15629
rect 10413 15589 10425 15623
rect 10459 15620 10471 15623
rect 10459 15592 11836 15620
rect 10459 15589 10471 15592
rect 10413 15583 10471 15589
rect 4332 15555 4390 15561
rect 4332 15521 4344 15555
rect 4378 15552 4390 15555
rect 4614 15552 4620 15564
rect 4378 15524 4620 15552
rect 4378 15521 4390 15524
rect 4332 15515 4390 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 5316 15524 5549 15552
rect 5316 15512 5322 15524
rect 5537 15521 5549 15524
rect 5583 15521 5595 15555
rect 5537 15515 5595 15521
rect 5804 15555 5862 15561
rect 5804 15521 5816 15555
rect 5850 15552 5862 15555
rect 6362 15552 6368 15564
rect 5850 15524 6368 15552
rect 5850 15521 5862 15524
rect 5804 15515 5862 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 9214 15552 9220 15564
rect 7515 15524 9220 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9456 15524 9505 15552
rect 9456 15512 9462 15524
rect 9493 15521 9505 15524
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 11054 15561 11060 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10100 15524 10333 15552
rect 10100 15512 10106 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 11048 15552 11060 15561
rect 11015 15524 11060 15552
rect 10321 15515 10379 15521
rect 11048 15515 11060 15524
rect 11054 15512 11060 15515
rect 11112 15512 11118 15564
rect 4062 15484 4068 15496
rect 3743 15456 3924 15484
rect 4023 15456 4068 15484
rect 3743 15453 3755 15456
rect 3697 15447 3755 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7064 15456 7573 15484
rect 7064 15444 7070 15456
rect 7561 15453 7573 15456
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2832 15320 2973 15348
rect 2832 15308 2838 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 2961 15311 3019 15317
rect 3053 15351 3111 15357
rect 3053 15317 3065 15351
rect 3099 15348 3111 15351
rect 3510 15348 3516 15360
rect 3099 15320 3516 15348
rect 3099 15317 3111 15320
rect 3053 15311 3111 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 5258 15308 5264 15360
rect 5316 15348 5322 15360
rect 5445 15351 5503 15357
rect 5445 15348 5457 15351
rect 5316 15320 5457 15348
rect 5316 15308 5322 15320
rect 5445 15317 5457 15320
rect 5491 15317 5503 15351
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 5445 15311 5503 15317
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 7576 15348 7604 15447
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 10781 15487 10839 15493
rect 10560 15456 10605 15484
rect 10560 15444 10566 15456
rect 10781 15453 10793 15487
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 8938 15416 8944 15428
rect 8899 15388 8944 15416
rect 8938 15376 8944 15388
rect 8996 15376 9002 15428
rect 9309 15419 9367 15425
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 9766 15416 9772 15428
rect 9355 15388 9772 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 9324 15348 9352 15379
rect 9766 15376 9772 15388
rect 9824 15416 9830 15428
rect 10796 15416 10824 15447
rect 9824 15388 10824 15416
rect 11808 15416 11836 15592
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 11940 15524 13001 15552
rect 11940 15512 11946 15524
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12434 15484 12440 15496
rect 12299 15456 12440 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12434 15444 12440 15456
rect 12492 15444 12498 15496
rect 12759 15487 12817 15493
rect 12759 15453 12771 15487
rect 12805 15484 12817 15487
rect 13446 15484 13452 15496
rect 12805 15456 13452 15484
rect 12805 15453 12817 15456
rect 12759 15447 12817 15453
rect 13446 15444 13452 15456
rect 13504 15484 13510 15496
rect 14568 15484 14596 15515
rect 13504 15456 14596 15484
rect 14737 15487 14795 15493
rect 13504 15444 13510 15456
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 11808 15388 12296 15416
rect 9824 15376 9830 15388
rect 7576 15320 9352 15348
rect 10796 15348 10824 15388
rect 11422 15348 11428 15360
rect 10796 15320 11428 15348
rect 11422 15308 11428 15320
rect 11480 15348 11486 15360
rect 12066 15348 12072 15360
rect 11480 15320 12072 15348
rect 11480 15308 11486 15320
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 12268 15348 12296 15388
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 14752 15416 14780 15447
rect 13872 15388 14780 15416
rect 13872 15376 13878 15388
rect 13906 15348 13912 15360
rect 12268 15320 13912 15348
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15348 14151 15351
rect 14844 15348 14872 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 19334 15688 19340 15700
rect 18739 15660 19340 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15657 20407 15691
rect 20349 15651 20407 15657
rect 20625 15691 20683 15697
rect 20625 15657 20637 15691
rect 20671 15688 20683 15691
rect 20990 15688 20996 15700
rect 20671 15660 20996 15688
rect 20671 15657 20683 15660
rect 20625 15651 20683 15657
rect 15556 15623 15614 15629
rect 15556 15589 15568 15623
rect 15602 15620 15614 15623
rect 17034 15620 17040 15632
rect 15602 15592 17040 15620
rect 15602 15589 15614 15592
rect 15556 15583 15614 15589
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 17580 15623 17638 15629
rect 17580 15589 17592 15623
rect 17626 15620 17638 15623
rect 19886 15620 19892 15632
rect 17626 15592 19892 15620
rect 17626 15589 17638 15592
rect 17580 15583 17638 15589
rect 19886 15580 19892 15592
rect 19944 15620 19950 15632
rect 20364 15620 20392 15651
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 23017 15691 23075 15697
rect 23017 15688 23029 15691
rect 22612 15660 23029 15688
rect 22612 15648 22618 15660
rect 23017 15657 23029 15660
rect 23063 15657 23075 15691
rect 23017 15651 23075 15657
rect 19944 15592 20392 15620
rect 21628 15623 21686 15629
rect 19944 15580 19950 15592
rect 21628 15589 21640 15623
rect 21674 15620 21686 15623
rect 22922 15620 22928 15632
rect 21674 15592 22928 15620
rect 21674 15589 21686 15592
rect 21628 15583 21686 15589
rect 22922 15580 22928 15592
rect 22980 15580 22986 15632
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 16390 15552 16396 15564
rect 15335 15524 16396 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 16390 15512 16396 15524
rect 16448 15552 16454 15564
rect 17218 15552 17224 15564
rect 16448 15524 16896 15552
rect 17179 15524 17224 15552
rect 16448 15512 16454 15524
rect 16758 15484 16764 15496
rect 16719 15456 16764 15484
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 16868 15484 16896 15524
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 18506 15552 18512 15564
rect 18104 15524 18512 15552
rect 18104 15512 18110 15524
rect 18506 15512 18512 15524
rect 18564 15552 18570 15564
rect 18969 15555 19027 15561
rect 18969 15552 18981 15555
rect 18564 15524 18981 15552
rect 18564 15512 18570 15524
rect 18969 15521 18981 15524
rect 19015 15521 19027 15555
rect 18969 15515 19027 15521
rect 19236 15555 19294 15561
rect 19236 15521 19248 15555
rect 19282 15552 19294 15555
rect 19978 15552 19984 15564
rect 19282 15524 19984 15552
rect 19282 15521 19294 15524
rect 19236 15515 19294 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20438 15552 20444 15564
rect 20399 15524 20444 15552
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15552 22891 15555
rect 23106 15552 23112 15564
rect 22879 15524 23112 15552
rect 22879 15521 22891 15524
rect 22833 15515 22891 15521
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 17313 15487 17371 15493
rect 17313 15484 17325 15487
rect 16868 15456 17325 15484
rect 17313 15453 17325 15456
rect 17359 15453 17371 15487
rect 21358 15484 21364 15496
rect 21319 15456 21364 15484
rect 17313 15447 17371 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 16666 15348 16672 15360
rect 14139 15320 14872 15348
rect 16627 15320 16672 15348
rect 14139 15317 14151 15320
rect 14093 15311 14151 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 17034 15348 17040 15360
rect 16995 15320 17040 15348
rect 17034 15308 17040 15320
rect 17092 15348 17098 15360
rect 17586 15348 17592 15360
rect 17092 15320 17592 15348
rect 17092 15308 17098 15320
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 17678 15308 17684 15360
rect 17736 15348 17742 15360
rect 19334 15348 19340 15360
rect 17736 15320 19340 15348
rect 17736 15308 17742 15320
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 22370 15308 22376 15360
rect 22428 15348 22434 15360
rect 22741 15351 22799 15357
rect 22741 15348 22753 15351
rect 22428 15320 22753 15348
rect 22428 15308 22434 15320
rect 22741 15317 22753 15320
rect 22787 15317 22799 15351
rect 22741 15311 22799 15317
rect 1104 15258 23460 15280
rect 1104 15206 4714 15258
rect 4766 15206 4778 15258
rect 4830 15206 4842 15258
rect 4894 15206 4906 15258
rect 4958 15206 12178 15258
rect 12230 15206 12242 15258
rect 12294 15206 12306 15258
rect 12358 15206 12370 15258
rect 12422 15206 19642 15258
rect 19694 15206 19706 15258
rect 19758 15206 19770 15258
rect 19822 15206 19834 15258
rect 19886 15206 23460 15258
rect 1104 15184 23460 15206
rect 6362 15144 6368 15156
rect 6323 15116 6368 15144
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 7650 15144 7656 15156
rect 6512 15116 6557 15144
rect 7611 15116 7656 15144
rect 6512 15104 6518 15116
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8754 15144 8760 15156
rect 8711 15116 8760 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 8849 15147 8907 15153
rect 8849 15113 8861 15147
rect 8895 15144 8907 15147
rect 9122 15144 9128 15156
rect 8895 15116 9128 15144
rect 8895 15113 8907 15116
rect 8849 15107 8907 15113
rect 4614 15036 4620 15088
rect 4672 15076 4678 15088
rect 4893 15079 4951 15085
rect 4893 15076 4905 15079
rect 4672 15048 4905 15076
rect 4672 15036 4678 15048
rect 4893 15045 4905 15048
rect 4939 15045 4951 15079
rect 4893 15039 4951 15045
rect 6825 15079 6883 15085
rect 6825 15045 6837 15079
rect 6871 15076 6883 15079
rect 6871 15048 8156 15076
rect 6871 15045 6883 15048
rect 6825 15039 6883 15045
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 8128 15017 8156 15048
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2038 14940 2044 14952
rect 1820 14912 2044 14940
rect 1820 14900 1826 14912
rect 2038 14900 2044 14912
rect 2096 14940 2102 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 2096 14912 3525 14940
rect 2096 14900 2102 14912
rect 3513 14909 3525 14912
rect 3559 14940 3571 14943
rect 4062 14940 4068 14952
rect 3559 14912 4068 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 4062 14900 4068 14912
rect 4120 14940 4126 14952
rect 5258 14949 5264 14952
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 4120 14912 4997 14940
rect 4120 14900 4126 14912
rect 4985 14909 4997 14912
rect 5031 14909 5043 14943
rect 5252 14940 5264 14949
rect 5219 14912 5264 14940
rect 4985 14903 5043 14909
rect 5252 14903 5264 14912
rect 5258 14900 5264 14903
rect 5316 14900 5322 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 8018 14940 8024 14952
rect 6687 14912 7880 14940
rect 7979 14912 8024 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 2308 14875 2366 14881
rect 2308 14841 2320 14875
rect 2354 14872 2366 14875
rect 3142 14872 3148 14884
rect 2354 14844 3148 14872
rect 2354 14841 2366 14844
rect 2308 14835 2366 14841
rect 3142 14832 3148 14844
rect 3200 14832 3206 14884
rect 3758 14875 3816 14881
rect 3758 14872 3770 14875
rect 3436 14844 3770 14872
rect 3436 14813 3464 14844
rect 3758 14841 3770 14844
rect 3804 14872 3816 14875
rect 4430 14872 4436 14884
rect 3804 14844 4436 14872
rect 3804 14841 3816 14844
rect 3758 14835 3816 14841
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 5166 14832 5172 14884
rect 5224 14872 5230 14884
rect 7285 14875 7343 14881
rect 7285 14872 7297 14875
rect 5224 14844 7297 14872
rect 5224 14832 5230 14844
rect 7285 14841 7297 14844
rect 7331 14841 7343 14875
rect 7852 14872 7880 14912
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8128 14940 8156 14971
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8260 14980 8305 15008
rect 8260 14968 8266 14980
rect 8481 14943 8539 14949
rect 8481 14940 8493 14943
rect 8128 14912 8493 14940
rect 8481 14909 8493 14912
rect 8527 14909 8539 14943
rect 8481 14903 8539 14909
rect 8864 14872 8892 15107
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9309 15147 9367 15153
rect 9309 15113 9321 15147
rect 9355 15144 9367 15147
rect 10502 15144 10508 15156
rect 9355 15116 10508 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11112 15116 11529 15144
rect 11112 15104 11118 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12584 15116 12817 15144
rect 12584 15104 12590 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 14550 15144 14556 15156
rect 14511 15116 14556 15144
rect 12805 15107 12863 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15654 15144 15660 15156
rect 15615 15116 15660 15144
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 17773 15147 17831 15153
rect 17773 15113 17785 15147
rect 17819 15144 17831 15147
rect 19334 15144 19340 15156
rect 17819 15116 19340 15144
rect 17819 15113 17831 15116
rect 17773 15107 17831 15113
rect 11701 15079 11759 15085
rect 11701 15045 11713 15079
rect 11747 15076 11759 15079
rect 12618 15076 12624 15088
rect 11747 15048 12624 15076
rect 11747 15045 11759 15048
rect 11701 15039 11759 15045
rect 9953 15011 10011 15017
rect 9953 14977 9965 15011
rect 9999 15008 10011 15011
rect 9999 14980 10272 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 9030 14940 9036 14952
rect 8991 14912 9036 14940
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 10137 14943 10195 14949
rect 10137 14940 10149 14943
rect 9732 14912 10149 14940
rect 9732 14900 9738 14912
rect 10137 14909 10149 14912
rect 10183 14909 10195 14943
rect 10244 14940 10272 14980
rect 11330 14940 11336 14952
rect 10244 14912 11336 14940
rect 10137 14903 10195 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11808 14949 11836 15048
rect 12618 15036 12624 15048
rect 12676 15036 12682 15088
rect 16206 15036 16212 15088
rect 16264 15076 16270 15088
rect 17497 15079 17555 15085
rect 17497 15076 17509 15079
rect 16264 15048 17509 15076
rect 16264 15036 16270 15048
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15378 15008 15384 15020
rect 15335 14980 15384 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 16298 15008 16304 15020
rect 16259 14980 16304 15008
rect 16298 14968 16304 14980
rect 16356 15008 16362 15020
rect 16666 15008 16672 15020
rect 16356 14980 16672 15008
rect 16356 14968 16362 14980
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 17052 15017 17080 15048
rect 17497 15045 17509 15048
rect 17543 15045 17555 15079
rect 17497 15039 17555 15045
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12207 14912 12449 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13262 14940 13268 14952
rect 13219 14912 13268 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 10410 14881 10416 14884
rect 10404 14872 10416 14881
rect 7852 14844 8892 14872
rect 10371 14844 10416 14872
rect 7285 14835 7343 14841
rect 10404 14835 10416 14844
rect 10410 14832 10416 14835
rect 10468 14832 10474 14884
rect 11974 14872 11980 14884
rect 11935 14844 11980 14872
rect 11974 14832 11980 14844
rect 12032 14832 12038 14884
rect 13004 14872 13032 14903
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13440 14943 13498 14949
rect 13440 14909 13452 14943
rect 13486 14940 13498 14943
rect 13814 14940 13820 14952
rect 13486 14912 13820 14940
rect 13486 14909 13498 14912
rect 13440 14903 13498 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14940 16083 14943
rect 16758 14940 16764 14952
rect 16071 14912 16764 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17788 14940 17816 15107
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 20036 15116 20085 15144
rect 20036 15104 20042 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 20806 15144 20812 15156
rect 20211 15116 20812 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 22278 15104 22284 15156
rect 22336 15144 22342 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22336 15116 23029 15144
rect 22336 15104 22342 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18598 15076 18604 15088
rect 18012 15048 18604 15076
rect 18012 15036 18018 15048
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 18690 15008 18696 15020
rect 18651 14980 18696 15008
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 20162 14968 20168 15020
rect 20220 15008 20226 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20220 14980 20729 15008
rect 20220 14968 20226 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 18046 14940 18052 14952
rect 17359 14912 17816 14940
rect 18007 14912 18052 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 21358 14940 21364 14952
rect 21319 14912 21364 14940
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 21628 14943 21686 14949
rect 21628 14909 21640 14943
rect 21674 14940 21686 14943
rect 22370 14940 22376 14952
rect 21674 14912 22376 14940
rect 21674 14909 21686 14912
rect 21628 14903 21686 14909
rect 22370 14900 22376 14912
rect 22428 14900 22434 14952
rect 22830 14940 22836 14952
rect 22791 14912 22836 14940
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 14458 14872 14464 14884
rect 13004 14844 14464 14872
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 15654 14872 15660 14884
rect 14660 14844 15660 14872
rect 3421 14807 3479 14813
rect 3421 14773 3433 14807
rect 3467 14773 3479 14807
rect 3421 14767 3479 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 7524 14776 9137 14804
rect 7524 14764 7530 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 9125 14767 9183 14773
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9456 14776 9689 14804
rect 9456 14764 9462 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9677 14767 9735 14773
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 9858 14804 9864 14816
rect 9815 14776 9864 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 12618 14804 12624 14816
rect 12579 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 14660 14813 14688 14844
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 16117 14875 16175 14881
rect 16117 14841 16129 14875
rect 16163 14872 16175 14875
rect 17126 14872 17132 14884
rect 16163 14844 17132 14872
rect 16163 14841 16175 14844
rect 16117 14835 16175 14841
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 18782 14872 18788 14884
rect 18248 14844 18788 14872
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15013 14807 15071 14813
rect 15013 14804 15025 14807
rect 14792 14776 15025 14804
rect 14792 14764 14798 14776
rect 15013 14773 15025 14776
rect 15059 14773 15071 14807
rect 15013 14767 15071 14773
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 16482 14804 16488 14816
rect 15160 14776 15205 14804
rect 16443 14776 16488 14804
rect 15160 14764 15166 14776
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16850 14804 16856 14816
rect 16811 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 16945 14807 17003 14813
rect 16945 14773 16957 14807
rect 16991 14804 17003 14807
rect 17218 14804 17224 14816
rect 16991 14776 17224 14804
rect 16991 14773 17003 14776
rect 16945 14767 17003 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 18248 14813 18276 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 18960 14875 19018 14881
rect 18960 14841 18972 14875
rect 19006 14872 19018 14875
rect 19794 14872 19800 14884
rect 19006 14844 19800 14872
rect 19006 14841 19018 14844
rect 18960 14835 19018 14841
rect 19794 14832 19800 14844
rect 19852 14872 19858 14884
rect 20533 14875 20591 14881
rect 20533 14872 20545 14875
rect 19852 14844 20545 14872
rect 19852 14832 19858 14844
rect 20533 14841 20545 14844
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14773 18291 14807
rect 18233 14767 18291 14773
rect 18509 14807 18567 14813
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 19334 14804 19340 14816
rect 18555 14776 19340 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 19484 14776 20637 14804
rect 19484 14764 19490 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20625 14767 20683 14773
rect 21085 14807 21143 14813
rect 21085 14773 21097 14807
rect 21131 14804 21143 14807
rect 22278 14804 22284 14816
rect 21131 14776 22284 14804
rect 21131 14773 21143 14776
rect 21085 14767 21143 14773
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 22741 14807 22799 14813
rect 22741 14773 22753 14807
rect 22787 14804 22799 14807
rect 22922 14804 22928 14816
rect 22787 14776 22928 14804
rect 22787 14773 22799 14776
rect 22741 14767 22799 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 1104 14714 23460 14736
rect 1104 14662 8446 14714
rect 8498 14662 8510 14714
rect 8562 14662 8574 14714
rect 8626 14662 8638 14714
rect 8690 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 23460 14714
rect 1104 14640 23460 14662
rect 3142 14600 3148 14612
rect 3103 14572 3148 14600
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3476 14572 4077 14600
rect 3476 14560 3482 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4430 14600 4436 14612
rect 4391 14572 4436 14600
rect 4065 14563 4123 14569
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14600 4951 14603
rect 5074 14600 5080 14612
rect 4939 14572 5080 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5258 14600 5264 14612
rect 5219 14572 5264 14600
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5718 14600 5724 14612
rect 5679 14572 5724 14600
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6362 14600 6368 14612
rect 6227 14572 6368 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10410 14560 10416 14612
rect 10468 14600 10474 14612
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 10468 14572 11069 14600
rect 10468 14560 10474 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 12710 14600 12716 14612
rect 11057 14563 11115 14569
rect 11164 14572 12716 14600
rect 2032 14535 2090 14541
rect 2032 14501 2044 14535
rect 2078 14532 2090 14535
rect 2774 14532 2780 14544
rect 2078 14504 2780 14532
rect 2078 14501 2090 14504
rect 2032 14495 2090 14501
rect 2774 14492 2780 14504
rect 2832 14492 2838 14544
rect 3160 14532 3188 14560
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 3160 14504 4537 14532
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 5353 14535 5411 14541
rect 5353 14532 5365 14535
rect 4672 14504 5365 14532
rect 4672 14492 4678 14504
rect 5353 14501 5365 14504
rect 5399 14501 5411 14535
rect 5353 14495 5411 14501
rect 6089 14535 6147 14541
rect 6089 14501 6101 14535
rect 6135 14532 6147 14535
rect 6914 14532 6920 14544
rect 6135 14504 6920 14532
rect 6135 14501 6147 14504
rect 6089 14495 6147 14501
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 7552 14535 7610 14541
rect 7552 14501 7564 14535
rect 7598 14532 7610 14535
rect 8110 14532 8116 14544
rect 7598 14504 8116 14532
rect 7598 14501 7610 14504
rect 7552 14495 7610 14501
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 9944 14535 10002 14541
rect 8864 14504 9904 14532
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 3510 14464 3516 14476
rect 3471 14436 3516 14464
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 7374 14464 7380 14476
rect 7331 14436 7380 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 8864 14473 8892 14504
rect 8849 14467 8907 14473
rect 8849 14433 8861 14467
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 9217 14467 9275 14473
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 9766 14464 9772 14476
rect 9263 14436 9772 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9876 14464 9904 14504
rect 9944 14501 9956 14535
rect 9990 14532 10002 14535
rect 11164 14532 11192 14572
rect 12710 14560 12716 14572
rect 12768 14560 12774 14612
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14569 15347 14603
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15289 14563 15347 14569
rect 13004 14532 13032 14563
rect 9990 14504 11192 14532
rect 11256 14504 13032 14532
rect 13624 14535 13682 14541
rect 9990 14501 10002 14504
rect 9944 14495 10002 14501
rect 10318 14464 10324 14476
rect 9876 14436 10324 14464
rect 10318 14424 10324 14436
rect 10376 14464 10382 14476
rect 10376 14436 10732 14464
rect 10376 14424 10382 14436
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4755 14368 5549 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5537 14365 5549 14368
rect 5583 14396 5595 14399
rect 6365 14399 6423 14405
rect 6365 14396 6377 14399
rect 5583 14368 6377 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 6365 14365 6377 14368
rect 6411 14396 6423 14399
rect 6546 14396 6552 14408
rect 6411 14368 6552 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10704 14396 10732 14436
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11256 14464 11284 14504
rect 13624 14501 13636 14535
rect 13670 14532 13682 14535
rect 14550 14532 14556 14544
rect 13670 14504 14556 14532
rect 13670 14501 13682 14504
rect 13624 14495 13682 14501
rect 14550 14492 14556 14504
rect 14608 14532 14614 14544
rect 15102 14532 15108 14544
rect 14608 14504 15108 14532
rect 14608 14492 14614 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 10928 14436 11284 14464
rect 11333 14467 11391 14473
rect 10928 14424 10934 14436
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11422 14464 11428 14476
rect 11379 14436 11428 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 11600 14467 11658 14473
rect 11600 14433 11612 14467
rect 11646 14464 11658 14467
rect 11974 14464 11980 14476
rect 11646 14436 11980 14464
rect 11646 14433 11658 14436
rect 11600 14427 11658 14433
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 12802 14464 12808 14476
rect 12763 14436 12808 14464
rect 12802 14424 12808 14436
rect 12860 14464 12866 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 12860 14436 13185 14464
rect 12860 14424 12866 14436
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14464 14887 14467
rect 15304 14464 15332 14563
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 19794 14600 19800 14612
rect 17092 14572 19472 14600
rect 19755 14572 19800 14600
rect 17092 14560 17098 14572
rect 19334 14532 19340 14544
rect 17788 14504 19340 14532
rect 14875 14436 15332 14464
rect 16301 14467 16359 14473
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 16301 14433 16313 14467
rect 16347 14464 16359 14467
rect 16390 14464 16396 14476
rect 16347 14436 16396 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16574 14473 16580 14476
rect 16568 14427 16580 14473
rect 16632 14464 16638 14476
rect 17788 14473 17816 14504
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 19444 14532 19472 14572
rect 19794 14560 19800 14572
rect 19852 14560 19858 14612
rect 20254 14600 20260 14612
rect 20215 14572 20260 14600
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 19444 14504 20116 14532
rect 17773 14467 17831 14473
rect 16632 14436 16668 14464
rect 16574 14424 16580 14427
rect 16632 14424 16638 14436
rect 17773 14433 17785 14467
rect 17819 14433 17831 14467
rect 17773 14427 17831 14433
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18288 14436 18337 14464
rect 18288 14424 18294 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14464 18475 14467
rect 18506 14464 18512 14476
rect 18463 14436 18512 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 18684 14467 18742 14473
rect 18684 14433 18696 14467
rect 18730 14464 18742 14467
rect 19426 14464 19432 14476
rect 18730 14436 19432 14464
rect 18730 14433 18742 14436
rect 18684 14427 18742 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 20088 14473 20116 14504
rect 20073 14467 20131 14473
rect 20073 14433 20085 14467
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21542 14464 21548 14476
rect 20947 14436 21548 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21542 14424 21548 14436
rect 21600 14424 21606 14476
rect 21904 14467 21962 14473
rect 21904 14433 21916 14467
rect 21950 14464 21962 14467
rect 22922 14464 22928 14476
rect 21950 14436 22928 14464
rect 21950 14433 21962 14436
rect 21904 14427 21962 14433
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10704 14368 11161 14396
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 11149 14359 11207 14365
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16206 14396 16212 14408
rect 15887 14368 16212 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 3697 14331 3755 14337
rect 3697 14297 3709 14331
rect 3743 14328 3755 14331
rect 5350 14328 5356 14340
rect 3743 14300 5356 14328
rect 3743 14297 3755 14300
rect 3697 14291 3755 14297
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15856 14328 15884 14359
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 21358 14396 21364 14408
rect 19904 14368 21364 14396
rect 15712 14300 15884 14328
rect 15712 14288 15718 14300
rect 17310 14288 17316 14340
rect 17368 14328 17374 14340
rect 18141 14331 18199 14337
rect 18141 14328 18153 14331
rect 17368 14300 18153 14328
rect 17368 14288 17374 14300
rect 18141 14297 18153 14300
rect 18187 14297 18199 14331
rect 18141 14291 18199 14297
rect 8662 14260 8668 14272
rect 8623 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9033 14263 9091 14269
rect 9033 14229 9045 14263
rect 9079 14260 9091 14263
rect 9398 14260 9404 14272
rect 9079 14232 9404 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 12710 14260 12716 14272
rect 12623 14232 12716 14260
rect 12710 14220 12716 14232
rect 12768 14260 12774 14272
rect 13998 14260 14004 14272
rect 12768 14232 14004 14260
rect 12768 14220 12774 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 15013 14263 15071 14269
rect 15013 14229 15025 14263
rect 15059 14260 15071 14263
rect 17034 14260 17040 14272
rect 15059 14232 17040 14260
rect 15059 14229 15071 14232
rect 15013 14223 15071 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 17678 14260 17684 14272
rect 17639 14232 17684 14260
rect 17678 14220 17684 14232
rect 17736 14220 17742 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 17957 14263 18015 14269
rect 17957 14260 17969 14263
rect 17920 14232 17969 14260
rect 17920 14220 17926 14232
rect 17957 14229 17969 14232
rect 18003 14229 18015 14263
rect 17957 14223 18015 14229
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19904 14269 19932 14368
rect 21358 14356 21364 14368
rect 21416 14396 21422 14408
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21416 14368 21649 14396
rect 21416 14356 21422 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 18656 14232 19901 14260
rect 18656 14220 18662 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 20346 14260 20352 14272
rect 20307 14232 20352 14260
rect 19889 14223 19947 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20588 14232 21097 14260
rect 20588 14220 20594 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 21085 14223 21143 14229
rect 22646 14220 22652 14272
rect 22704 14260 22710 14272
rect 23017 14263 23075 14269
rect 23017 14260 23029 14263
rect 22704 14232 23029 14260
rect 22704 14220 22710 14232
rect 23017 14229 23029 14232
rect 23063 14229 23075 14263
rect 23017 14223 23075 14229
rect 1104 14170 23460 14192
rect 1104 14118 4714 14170
rect 4766 14118 4778 14170
rect 4830 14118 4842 14170
rect 4894 14118 4906 14170
rect 4958 14118 12178 14170
rect 12230 14118 12242 14170
rect 12294 14118 12306 14170
rect 12358 14118 12370 14170
rect 12422 14118 19642 14170
rect 19694 14118 19706 14170
rect 19758 14118 19770 14170
rect 19822 14118 19834 14170
rect 19886 14118 23460 14170
rect 1104 14096 23460 14118
rect 1762 14056 1768 14068
rect 1504 14028 1768 14056
rect 1504 13929 1532 14028
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2958 14056 2964 14068
rect 2919 14028 2964 14056
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 5166 14056 5172 14068
rect 4847 14028 5172 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 11790 14056 11796 14068
rect 10551 14028 11796 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 13446 14056 13452 14068
rect 12268 14028 12480 14056
rect 13407 14028 13452 14056
rect 2869 13991 2927 13997
rect 2869 13957 2881 13991
rect 2915 13988 2927 13991
rect 3050 13988 3056 14000
rect 2915 13960 3056 13988
rect 2915 13957 2927 13960
rect 2869 13951 2927 13957
rect 3050 13948 3056 13960
rect 3108 13988 3114 14000
rect 3789 13991 3847 13997
rect 3108 13960 3464 13988
rect 3108 13948 3114 13960
rect 3436 13929 3464 13960
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 5077 13991 5135 13997
rect 3835 13960 4660 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 1489 13923 1547 13929
rect 1489 13889 1501 13923
rect 1535 13889 1547 13923
rect 1489 13883 1547 13889
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3602 13920 3608 13932
rect 3563 13892 3608 13920
rect 3421 13883 3479 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4522 13920 4528 13932
rect 4479 13892 4528 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4632 13861 4660 13960
rect 5077 13957 5089 13991
rect 5123 13988 5135 13991
rect 6730 13988 6736 14000
rect 5123 13960 6736 13988
rect 5123 13957 5135 13960
rect 5077 13951 5135 13957
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 8849 13991 8907 13997
rect 8849 13957 8861 13991
rect 8895 13988 8907 13991
rect 10134 13988 10140 14000
rect 8895 13960 10140 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 11333 13991 11391 13997
rect 10376 13960 11192 13988
rect 10376 13948 10382 13960
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5592 13892 5733 13920
rect 5592 13880 5598 13892
rect 5721 13889 5733 13892
rect 5767 13920 5779 13923
rect 6546 13920 6552 13932
rect 5767 13892 6552 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 9398 13920 9404 13932
rect 9359 13892 9404 13920
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 10226 13920 10232 13932
rect 10139 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10870 13920 10876 13932
rect 10284 13892 10876 13920
rect 10284 13880 10290 13892
rect 10870 13880 10876 13892
rect 10928 13920 10934 13932
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 10928 13892 11069 13920
rect 10928 13880 10934 13892
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 11164 13920 11192 13960
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 12268 13988 12296 14028
rect 11379 13960 12296 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11164 13892 11805 13920
rect 11057 13883 11115 13889
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13821 4675 13855
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 4617 13815 4675 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7374 13852 7380 13864
rect 7335 13824 7380 13852
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 7644 13855 7702 13861
rect 7644 13821 7656 13855
rect 7690 13852 7702 13855
rect 8662 13852 8668 13864
rect 7690 13824 8668 13852
rect 7690 13821 7702 13824
rect 7644 13815 7702 13821
rect 8662 13812 8668 13824
rect 8720 13852 8726 13864
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 8720 13824 9321 13852
rect 8720 13812 8726 13824
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 9674 13812 9680 13864
rect 9732 13812 9738 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 10008 13824 10149 13852
rect 10008 13812 10014 13824
rect 10137 13821 10149 13824
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11330 13852 11336 13864
rect 11011 13824 11336 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11900 13852 11928 13883
rect 11480 13824 11928 13852
rect 12452 13852 12480 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 15010 14056 15016 14068
rect 14516 14028 15016 14056
rect 14516 14016 14522 14028
rect 15010 14016 15016 14028
rect 15068 14056 15074 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 15068 14028 15117 14056
rect 15068 14016 15074 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 17954 14056 17960 14068
rect 15105 14019 15163 14025
rect 15212 14028 17960 14056
rect 15212 13988 15240 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 19426 14056 19432 14068
rect 18104 14028 19012 14056
rect 19387 14028 19432 14056
rect 18104 14016 18110 14028
rect 14660 13960 15240 13988
rect 17681 13991 17739 13997
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12676 13892 13001 13920
rect 12676 13880 12682 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12452 13824 12817 13852
rect 11480 13812 11486 13824
rect 12805 13821 12817 13824
rect 12851 13852 12863 13855
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12851 13824 13277 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13852 13875 13855
rect 14660 13852 14688 13960
rect 17681 13957 17693 13991
rect 17727 13988 17739 13991
rect 17770 13988 17776 14000
rect 17727 13960 17776 13988
rect 17727 13957 17739 13960
rect 17681 13951 17739 13957
rect 17770 13948 17776 13960
rect 17828 13948 17834 14000
rect 18984 13988 19012 14028
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 20438 14016 20444 14068
rect 20496 14056 20502 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 20496 14028 21833 14056
rect 20496 14016 20502 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 21821 14019 21879 14025
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 18984 13960 19901 13988
rect 19889 13957 19901 13960
rect 19935 13957 19947 13991
rect 19889 13951 19947 13957
rect 21913 13991 21971 13997
rect 21913 13957 21925 13991
rect 21959 13988 21971 13991
rect 23106 13988 23112 14000
rect 21959 13960 23112 13988
rect 21959 13957 21971 13960
rect 21913 13951 21971 13957
rect 23106 13948 23112 13960
rect 23164 13948 23170 14000
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 20254 13920 20260 13932
rect 14792 13892 15792 13920
rect 14792 13880 14798 13892
rect 13863 13824 14688 13852
rect 15657 13855 15715 13861
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 15657 13821 15669 13855
rect 15703 13821 15715 13855
rect 15764 13852 15792 13892
rect 19536 13892 20260 13920
rect 15913 13855 15971 13861
rect 15913 13852 15925 13855
rect 15764 13824 15925 13852
rect 15657 13815 15715 13821
rect 15913 13821 15925 13824
rect 15959 13821 15971 13855
rect 15913 13815 15971 13821
rect 1756 13787 1814 13793
rect 1756 13753 1768 13787
rect 1802 13784 1814 13787
rect 2682 13784 2688 13796
rect 1802 13756 2688 13784
rect 1802 13753 1814 13756
rect 1756 13747 1814 13753
rect 2682 13744 2688 13756
rect 2740 13744 2746 13796
rect 2774 13744 2780 13796
rect 2832 13784 2838 13796
rect 3329 13787 3387 13793
rect 3329 13784 3341 13787
rect 2832 13756 3341 13784
rect 2832 13744 2838 13756
rect 3329 13753 3341 13756
rect 3375 13753 3387 13787
rect 3329 13747 3387 13753
rect 3510 13744 3516 13796
rect 3568 13784 3574 13796
rect 4249 13787 4307 13793
rect 4249 13784 4261 13787
rect 3568 13756 4261 13784
rect 3568 13744 3574 13756
rect 4249 13753 4261 13756
rect 4295 13753 4307 13787
rect 4249 13747 4307 13753
rect 5445 13787 5503 13793
rect 5445 13753 5457 13787
rect 5491 13784 5503 13787
rect 6086 13784 6092 13796
rect 5491 13756 6092 13784
rect 5491 13753 5503 13756
rect 5445 13747 5503 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 6270 13784 6276 13796
rect 6231 13756 6276 13784
rect 6270 13744 6276 13756
rect 6328 13744 6334 13796
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 8772 13756 9229 13784
rect 8772 13728 8800 13756
rect 9217 13753 9229 13756
rect 9263 13753 9275 13787
rect 9692 13784 9720 13812
rect 10686 13784 10692 13796
rect 9692 13756 10692 13784
rect 9217 13747 9275 13753
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 11701 13787 11759 13793
rect 11701 13753 11713 13787
rect 11747 13784 11759 13787
rect 12618 13784 12624 13796
rect 11747 13756 12624 13784
rect 11747 13753 11759 13756
rect 11701 13747 11759 13753
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 12894 13784 12900 13796
rect 12855 13756 12900 13784
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 15672 13784 15700 13815
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 16540 13824 17141 13852
rect 16540 13812 16546 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 17497 13855 17555 13861
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 17586 13852 17592 13864
rect 17543 13824 17592 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 18322 13861 18328 13864
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18316 13852 18328 13861
rect 18283 13824 18328 13852
rect 18049 13815 18107 13821
rect 18316 13815 18328 13824
rect 16390 13784 16396 13796
rect 15344 13756 16396 13784
rect 15344 13744 15350 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 18064 13784 18092 13815
rect 18322 13812 18328 13815
rect 18380 13812 18386 13864
rect 19536 13861 19564 13892
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 20530 13929 20536 13932
rect 20487 13923 20536 13929
rect 20487 13889 20499 13923
rect 20533 13889 20536 13923
rect 20487 13883 20536 13889
rect 20530 13880 20536 13883
rect 20588 13880 20594 13932
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22244 13892 22385 13920
rect 22244 13880 22250 13892
rect 22373 13889 22385 13892
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13821 19579 13855
rect 19521 13815 19579 13821
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13852 20039 13855
rect 20070 13852 20076 13864
rect 20027 13824 20076 13852
rect 20027 13821 20039 13824
rect 19981 13815 20039 13821
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 20714 13852 20720 13864
rect 20675 13824 20720 13852
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 22278 13852 22284 13864
rect 22239 13824 22284 13852
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 22572 13852 22600 13883
rect 22520 13824 22600 13852
rect 22520 13812 22526 13824
rect 18506 13784 18512 13796
rect 18064 13756 18512 13784
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 19610 13744 19616 13796
rect 19668 13784 19674 13796
rect 19705 13787 19763 13793
rect 19705 13784 19717 13787
rect 19668 13756 19717 13784
rect 19668 13744 19674 13756
rect 19705 13753 19717 13756
rect 19751 13753 19763 13787
rect 19705 13747 19763 13753
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 4120 13688 4169 13716
rect 4120 13676 4126 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4157 13679 4215 13685
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5316 13688 5549 13716
rect 5316 13676 5322 13688
rect 5537 13685 5549 13688
rect 5583 13685 5595 13719
rect 5537 13679 5595 13685
rect 5905 13719 5963 13725
rect 5905 13685 5917 13719
rect 5951 13716 5963 13719
rect 6178 13716 6184 13728
rect 5951 13688 6184 13716
rect 5951 13685 5963 13688
rect 5905 13679 5963 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 8754 13716 8760 13728
rect 6420 13688 6465 13716
rect 8715 13688 8760 13716
rect 6420 13676 6426 13688
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 9674 13716 9680 13728
rect 9635 13688 9680 13716
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 10410 13716 10416 13728
rect 10091 13688 10416 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10870 13716 10876 13728
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12492 13688 12537 13716
rect 12492 13676 12498 13688
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 15304 13716 15332 13744
rect 17034 13716 17040 13728
rect 13412 13688 15332 13716
rect 16995 13688 17040 13716
rect 13412 13676 13418 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17310 13716 17316 13728
rect 17271 13688 17316 13716
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 20254 13676 20260 13728
rect 20312 13716 20318 13728
rect 20447 13719 20505 13725
rect 20447 13716 20459 13719
rect 20312 13688 20459 13716
rect 20312 13676 20318 13688
rect 20447 13685 20459 13688
rect 20493 13685 20505 13719
rect 22738 13716 22744 13728
rect 22699 13688 22744 13716
rect 20447 13679 20505 13685
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 1104 13626 23460 13648
rect 1104 13574 8446 13626
rect 8498 13574 8510 13626
rect 8562 13574 8574 13626
rect 8626 13574 8638 13626
rect 8690 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 23460 13626
rect 1104 13552 23460 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 3510 13512 3516 13524
rect 2915 13484 3516 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4062 13512 4068 13524
rect 4023 13484 4068 13512
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 6822 13512 6828 13524
rect 6503 13484 6828 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13481 9735 13515
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 9677 13475 9735 13481
rect 3237 13447 3295 13453
rect 3237 13413 3249 13447
rect 3283 13444 3295 13447
rect 3418 13444 3424 13456
rect 3283 13416 3424 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 5442 13444 5448 13456
rect 4908 13416 5448 13444
rect 4430 13376 4436 13388
rect 4391 13348 4436 13376
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 3326 13308 3332 13320
rect 3287 13280 3332 13308
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 3528 13240 3556 13271
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4028 13280 4537 13308
rect 4028 13268 4034 13280
rect 4525 13277 4537 13280
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 4908 13308 4936 13416
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 6917 13447 6975 13453
rect 6917 13444 6929 13447
rect 6788 13416 6929 13444
rect 6788 13404 6794 13416
rect 6917 13413 6929 13416
rect 6963 13413 6975 13447
rect 6917 13407 6975 13413
rect 7644 13447 7702 13453
rect 7644 13413 7656 13447
rect 7690 13444 7702 13447
rect 8754 13444 8760 13456
rect 7690 13416 8760 13444
rect 7690 13413 7702 13416
rect 7644 13407 7702 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 9692 13444 9720 13475
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 10928 13484 12357 13512
rect 10928 13472 10934 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 12345 13475 12403 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 16942 13472 16948 13524
rect 17000 13472 17006 13524
rect 18506 13472 18512 13524
rect 18564 13472 18570 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 19242 13512 19248 13524
rect 18932 13484 19248 13512
rect 18932 13472 18938 13484
rect 19242 13472 19248 13484
rect 19300 13512 19306 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19300 13484 19809 13512
rect 19300 13472 19306 13484
rect 19797 13481 19809 13484
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 20349 13515 20407 13521
rect 20349 13481 20361 13515
rect 20395 13512 20407 13515
rect 20530 13512 20536 13524
rect 20395 13484 20536 13512
rect 20395 13481 20407 13484
rect 20349 13475 20407 13481
rect 12434 13444 12440 13456
rect 8864 13416 9720 13444
rect 9968 13416 12440 13444
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5074 13376 5080 13388
rect 5031 13348 5080 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5252 13379 5310 13385
rect 5252 13345 5264 13379
rect 5298 13376 5310 13379
rect 6086 13376 6092 13388
rect 5298 13348 6092 13376
rect 5298 13345 5310 13348
rect 5252 13339 5310 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6178 13336 6184 13388
rect 6236 13376 6242 13388
rect 8864 13385 8892 13416
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6236 13348 6837 13376
rect 6236 13336 6242 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 8849 13379 8907 13385
rect 8849 13345 8861 13379
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9968 13376 9996 13416
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 13354 13404 13360 13456
rect 13412 13404 13418 13456
rect 15556 13447 15614 13453
rect 15556 13413 15568 13447
rect 15602 13444 15614 13447
rect 16960 13444 16988 13472
rect 15602 13416 16988 13444
rect 17028 13447 17086 13453
rect 15602 13413 15614 13416
rect 15556 13407 15614 13413
rect 17028 13413 17040 13447
rect 17074 13444 17086 13447
rect 17678 13444 17684 13456
rect 17074 13416 17684 13444
rect 17074 13413 17086 13416
rect 17028 13407 17086 13413
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 18524 13444 18552 13472
rect 18064 13416 18552 13444
rect 19812 13444 19840 13475
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 22554 13512 22560 13524
rect 20640 13484 22560 13512
rect 20438 13444 20444 13456
rect 19812 13416 20444 13444
rect 9263 13348 9996 13376
rect 10045 13379 10103 13385
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 10045 13345 10057 13379
rect 10091 13345 10103 13379
rect 10502 13376 10508 13388
rect 10463 13348 10508 13376
rect 10045 13339 10103 13345
rect 4755 13280 4936 13308
rect 7009 13311 7067 13317
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7374 13308 7380 13320
rect 7335 13280 7380 13308
rect 7009 13271 7067 13277
rect 3602 13240 3608 13252
rect 3515 13212 3608 13240
rect 3602 13200 3608 13212
rect 3660 13240 3666 13252
rect 4724 13240 4752 13271
rect 7024 13240 7052 13271
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 10060 13308 10088 13339
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 11140 13379 11198 13385
rect 11140 13345 11152 13379
rect 11186 13376 11198 13379
rect 11882 13376 11888 13388
rect 11186 13348 11888 13376
rect 11186 13345 11198 13348
rect 11140 13339 11198 13345
rect 11882 13336 11888 13348
rect 11940 13376 11946 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 11940 13348 12725 13376
rect 11940 13336 11946 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13173 13379 13231 13385
rect 13173 13376 13185 13379
rect 13044 13348 13185 13376
rect 13044 13336 13050 13348
rect 13173 13345 13185 13348
rect 13219 13376 13231 13379
rect 13372 13376 13400 13404
rect 13219 13348 13400 13376
rect 13440 13379 13498 13385
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 13440 13345 13452 13379
rect 13486 13376 13498 13379
rect 14366 13376 14372 13388
rect 13486 13348 14372 13376
rect 13486 13345 13498 13348
rect 13440 13339 13498 13345
rect 14366 13336 14372 13348
rect 14424 13336 14430 13388
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 14829 13379 14887 13385
rect 14829 13376 14841 13379
rect 14516 13348 14841 13376
rect 14516 13336 14522 13348
rect 14829 13345 14841 13348
rect 14875 13345 14887 13379
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 14829 13339 14887 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15838 13376 15844 13388
rect 15436 13348 15844 13376
rect 15436 13336 15442 13348
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18064 13376 18092 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 18489 13379 18547 13385
rect 18489 13376 18501 13379
rect 16807 13348 18092 13376
rect 18156 13348 18501 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 10226 13308 10232 13320
rect 8996 13280 10088 13308
rect 10187 13280 10232 13308
rect 8996 13268 9002 13280
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10686 13268 10692 13320
rect 10744 13308 10750 13320
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10744 13280 10885 13308
rect 10744 13268 10750 13280
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12805 13311 12863 13317
rect 12805 13308 12817 13311
rect 12400 13280 12817 13308
rect 12400 13268 12406 13280
rect 12805 13277 12817 13280
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 3660 13212 4752 13240
rect 5920 13212 7052 13240
rect 9033 13243 9091 13249
rect 3660 13200 3666 13212
rect 4522 13132 4528 13184
rect 4580 13172 4586 13184
rect 5920 13172 5948 13212
rect 9033 13209 9045 13243
rect 9079 13240 9091 13243
rect 9858 13240 9864 13252
rect 9079 13212 9864 13240
rect 9079 13209 9091 13212
rect 9033 13203 9091 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12253 13243 12311 13249
rect 12253 13240 12265 13243
rect 12032 13212 12265 13240
rect 12032 13200 12038 13212
rect 12253 13209 12265 13212
rect 12299 13209 12311 13243
rect 12253 13203 12311 13209
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 12912 13240 12940 13271
rect 14826 13240 14832 13252
rect 12584 13212 12940 13240
rect 14108 13212 14832 13240
rect 12584 13200 12590 13212
rect 6362 13172 6368 13184
rect 4580 13144 5948 13172
rect 6323 13144 6368 13172
rect 4580 13132 4586 13144
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 8754 13172 8760 13184
rect 8715 13144 8760 13172
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 10594 13172 10600 13184
rect 9447 13144 10600 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 14108 13172 14136 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 10735 13144 14136 13172
rect 15013 13175 15071 13181
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 16206 13172 16212 13184
rect 15059 13144 16212 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 18156 13181 18184 13348
rect 18489 13345 18501 13348
rect 18535 13345 18547 13379
rect 18489 13339 18547 13345
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20640 13376 20668 13484
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 21168 13447 21226 13453
rect 21168 13413 21180 13447
rect 21214 13444 21226 13447
rect 22646 13444 22652 13456
rect 21214 13416 22652 13444
rect 21214 13413 21226 13416
rect 21168 13407 21226 13413
rect 22646 13404 22652 13416
rect 22704 13404 22710 13456
rect 22741 13447 22799 13453
rect 22741 13413 22753 13447
rect 22787 13444 22799 13447
rect 23106 13444 23112 13456
rect 22787 13416 23112 13444
rect 22787 13413 22799 13416
rect 22741 13407 22799 13413
rect 23106 13404 23112 13416
rect 23164 13404 23170 13456
rect 20404 13348 20668 13376
rect 20404 13336 20410 13348
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 22002 13376 22008 13388
rect 20772 13348 22008 13376
rect 20772 13336 20778 13348
rect 22002 13336 22008 13348
rect 22060 13376 22066 13388
rect 22833 13379 22891 13385
rect 22833 13376 22845 13379
rect 22060 13348 22845 13376
rect 22060 13336 22066 13348
rect 22833 13345 22845 13348
rect 22879 13345 22891 13379
rect 22833 13339 22891 13345
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 20625 13271 20683 13277
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 18012 13144 18153 13172
rect 18012 13132 18018 13144
rect 18141 13141 18153 13144
rect 18187 13141 18199 13175
rect 18248 13172 18276 13271
rect 18506 13172 18512 13184
rect 18248 13144 18512 13172
rect 18141 13135 18199 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19576 13144 19625 13172
rect 19576 13132 19582 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20162 13172 20168 13184
rect 20027 13144 20168 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 20640 13172 20668 13271
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 22922 13268 22928 13320
rect 22980 13308 22986 13320
rect 22980 13280 23025 13308
rect 22980 13268 22986 13280
rect 20806 13172 20812 13184
rect 20640 13144 20812 13172
rect 20806 13132 20812 13144
rect 20864 13172 20870 13184
rect 22281 13175 22339 13181
rect 22281 13172 22293 13175
rect 20864 13144 22293 13172
rect 20864 13132 20870 13144
rect 22281 13141 22293 13144
rect 22327 13141 22339 13175
rect 22281 13135 22339 13141
rect 22373 13175 22431 13181
rect 22373 13141 22385 13175
rect 22419 13172 22431 13175
rect 22462 13172 22468 13184
rect 22419 13144 22468 13172
rect 22419 13141 22431 13144
rect 22373 13135 22431 13141
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 1104 13082 23460 13104
rect 1104 13030 4714 13082
rect 4766 13030 4778 13082
rect 4830 13030 4842 13082
rect 4894 13030 4906 13082
rect 4958 13030 12178 13082
rect 12230 13030 12242 13082
rect 12294 13030 12306 13082
rect 12358 13030 12370 13082
rect 12422 13030 19642 13082
rect 19694 13030 19706 13082
rect 19758 13030 19770 13082
rect 19822 13030 19834 13082
rect 19886 13030 23460 13082
rect 1104 13008 23460 13030
rect 3970 12968 3976 12980
rect 3931 12940 3976 12968
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 5074 12968 5080 12980
rect 4724 12940 5080 12968
rect 4062 12900 4068 12912
rect 3975 12872 4068 12900
rect 4062 12860 4068 12872
rect 4120 12900 4126 12912
rect 4724 12900 4752 12940
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 6086 12968 6092 12980
rect 6047 12940 6092 12968
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 9122 12968 9128 12980
rect 6656 12940 9128 12968
rect 4120 12872 4752 12900
rect 4120 12860 4126 12872
rect 4724 12841 4752 12872
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 2038 12724 2044 12776
rect 2096 12764 2102 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2096 12736 2605 12764
rect 2096 12724 2102 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4249 12727 4307 12733
rect 4976 12767 5034 12773
rect 4976 12733 4988 12767
rect 5022 12764 5034 12767
rect 5258 12764 5264 12776
rect 5022 12736 5264 12764
rect 5022 12733 5034 12736
rect 4976 12727 5034 12733
rect 2608 12628 2636 12727
rect 2860 12699 2918 12705
rect 2860 12665 2872 12699
rect 2906 12696 2918 12699
rect 3418 12696 3424 12708
rect 2906 12668 3424 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 4062 12628 4068 12640
rect 2608 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4264 12628 4292 12727
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 6656 12773 6684 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 9766 12968 9772 12980
rect 9723 12940 9772 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10962 12968 10968 12980
rect 9876 12940 10968 12968
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 8938 12900 8944 12912
rect 8803 12872 8944 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9398 12900 9404 12912
rect 9324 12872 9404 12900
rect 9324 12841 9352 12872
rect 9398 12860 9404 12872
rect 9456 12900 9462 12912
rect 9876 12900 9904 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11940 12940 11989 12968
rect 11940 12928 11946 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 11977 12931 12035 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 14366 12968 14372 12980
rect 14327 12940 14372 12968
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 15289 12971 15347 12977
rect 15289 12937 15301 12971
rect 15335 12968 15347 12971
rect 15746 12968 15752 12980
rect 15335 12940 15752 12968
rect 15335 12937 15347 12940
rect 15289 12931 15347 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 16908 12940 16957 12968
rect 16908 12928 16914 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17644 12940 17785 12968
rect 17644 12928 17650 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 20346 12968 20352 12980
rect 19751 12940 20352 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 20898 12968 20904 12980
rect 20548 12940 20904 12968
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 9456 12872 9904 12900
rect 11624 12872 12081 12900
rect 9456 12860 9462 12872
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12801 9367 12835
rect 10226 12832 10232 12844
rect 10187 12804 10232 12832
rect 9309 12795 9367 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7374 12764 7380 12776
rect 7331 12736 7380 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7208 12696 7236 12727
rect 6472 12668 7236 12696
rect 6472 12637 6500 12668
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 4264 12600 6469 12628
rect 6457 12597 6469 12600
rect 6503 12597 6515 12631
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 6457 12591 6515 12597
rect 7006 12588 7012 12600
rect 7064 12628 7070 12640
rect 7300 12628 7328 12727
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7552 12767 7610 12773
rect 7552 12733 7564 12767
rect 7598 12764 7610 12767
rect 8754 12764 8760 12776
rect 7598 12736 8760 12764
rect 7598 12733 7610 12736
rect 7552 12727 7610 12733
rect 8754 12724 8760 12736
rect 8812 12764 8818 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8812 12736 9229 12764
rect 8812 12724 8818 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10686 12764 10692 12776
rect 10643 12736 10692 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10686 12724 10692 12736
rect 10744 12764 10750 12776
rect 11624 12764 11652 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 14384 12900 14412 12928
rect 16117 12903 16175 12909
rect 14384 12872 15700 12900
rect 12069 12863 12127 12869
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12986 12832 12992 12844
rect 11848 12804 12480 12832
rect 12947 12804 12992 12832
rect 11848 12792 11854 12804
rect 10744 12736 11652 12764
rect 10744 12724 10750 12736
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 12452 12773 12480 12804
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14056 12804 15025 12832
rect 14056 12792 14062 12804
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 15672 12773 15700 12872
rect 16117 12869 16129 12903
rect 16163 12900 16175 12903
rect 17218 12900 17224 12912
rect 16163 12872 17224 12900
rect 16163 12869 16175 12872
rect 16117 12863 16175 12869
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 17862 12900 17868 12912
rect 17328 12872 17868 12900
rect 15838 12832 15844 12844
rect 15799 12804 15844 12832
rect 15838 12792 15844 12804
rect 15896 12832 15902 12844
rect 16390 12832 16396 12844
rect 15896 12804 16396 12832
rect 15896 12792 15902 12804
rect 16390 12792 16396 12804
rect 16448 12832 16454 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16448 12804 16681 12832
rect 16448 12792 16454 12804
rect 16669 12801 16681 12804
rect 16715 12832 16727 12835
rect 17328 12832 17356 12872
rect 17512 12841 17540 12872
rect 17862 12860 17868 12872
rect 17920 12860 17926 12912
rect 16715 12804 17356 12832
rect 17497 12835 17555 12841
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 20162 12832 20168 12844
rect 20123 12804 20168 12832
rect 17497 12795 17555 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 20438 12832 20444 12844
rect 20395 12804 20444 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 11756 12736 12265 12764
rect 11756 12724 11762 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 12437 12727 12495 12733
rect 13188 12736 14933 12764
rect 9125 12699 9183 12705
rect 9125 12696 9137 12699
rect 8680 12668 9137 12696
rect 7064 12600 7328 12628
rect 7064 12588 7070 12600
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8680 12637 8708 12668
rect 9125 12665 9137 12668
rect 9171 12665 9183 12699
rect 9125 12659 9183 12665
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 9824 12668 10149 12696
rect 9824 12656 9830 12668
rect 10137 12665 10149 12668
rect 10183 12665 10195 12699
rect 10137 12659 10195 12665
rect 10864 12699 10922 12705
rect 10864 12665 10876 12699
rect 10910 12696 10922 12699
rect 12066 12696 12072 12708
rect 10910 12668 12072 12696
rect 10910 12665 10922 12668
rect 10864 12659 10922 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8352 12600 8677 12628
rect 8352 12588 8358 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8665 12591 8723 12597
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9916 12600 10057 12628
rect 9916 12588 9922 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 10045 12591 10103 12597
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 13188 12628 13216 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 15657 12767 15715 12773
rect 15657 12733 15669 12767
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 16485 12767 16543 12773
rect 16485 12733 16497 12767
rect 16531 12764 16543 12767
rect 16574 12764 16580 12776
rect 16531 12736 16580 12764
rect 16531 12733 16543 12736
rect 16485 12727 16543 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12764 17371 12767
rect 17954 12764 17960 12776
rect 17359 12736 17960 12764
rect 17359 12733 17371 12736
rect 17313 12727 17371 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18316 12767 18374 12773
rect 18316 12733 18328 12767
rect 18362 12764 18374 12767
rect 19518 12764 19524 12776
rect 18362 12736 19524 12764
rect 18362 12733 18374 12736
rect 18316 12727 18374 12733
rect 13256 12699 13314 12705
rect 13256 12665 13268 12699
rect 13302 12696 13314 12699
rect 14642 12696 14648 12708
rect 13302 12668 14648 12696
rect 13302 12665 13314 12668
rect 13256 12659 13314 12665
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 14826 12696 14832 12708
rect 14787 12668 14832 12696
rect 14826 12656 14832 12668
rect 14884 12656 14890 12708
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 17678 12696 17684 12708
rect 17451 12668 17684 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 18064 12696 18092 12727
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 20548 12773 20576 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 21232 12940 22017 12968
rect 21232 12928 21238 12940
rect 22005 12937 22017 12940
rect 22051 12968 22063 12971
rect 23290 12968 23296 12980
rect 22051 12940 23296 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 22462 12832 22468 12844
rect 22423 12804 22468 12832
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 22646 12832 22652 12844
rect 22607 12804 22652 12832
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 20806 12773 20812 12776
rect 20533 12767 20591 12773
rect 20533 12764 20545 12767
rect 20272 12736 20545 12764
rect 18506 12696 18512 12708
rect 18064 12668 18512 12696
rect 18506 12656 18512 12668
rect 18564 12696 18570 12708
rect 20272 12696 20300 12736
rect 20533 12733 20545 12736
rect 20579 12733 20591 12767
rect 20800 12764 20812 12773
rect 20767 12736 20812 12764
rect 20533 12727 20591 12733
rect 20800 12727 20812 12736
rect 20806 12724 20812 12727
rect 20864 12724 20870 12776
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12764 22431 12767
rect 22738 12764 22744 12776
rect 22419 12736 22744 12764
rect 22419 12733 22431 12736
rect 22373 12727 22431 12733
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 18564 12668 20300 12696
rect 18564 12656 18570 12668
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20990 12696 20996 12708
rect 20496 12668 20996 12696
rect 20496 12656 20502 12668
rect 20990 12656 20996 12668
rect 21048 12656 21054 12708
rect 22833 12699 22891 12705
rect 22833 12696 22845 12699
rect 21100 12668 22845 12696
rect 10652 12600 13216 12628
rect 10652 12588 10658 12600
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 13964 12600 14473 12628
rect 13964 12588 13970 12600
rect 14461 12597 14473 12600
rect 14507 12597 14519 12631
rect 14461 12591 14519 12597
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15160 12600 15761 12628
rect 15160 12588 15166 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 16577 12631 16635 12637
rect 16577 12597 16589 12631
rect 16623 12628 16635 12631
rect 17034 12628 17040 12640
rect 16623 12600 17040 12628
rect 16623 12597 16635 12600
rect 16577 12591 16635 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12628 19487 12631
rect 19610 12628 19616 12640
rect 19475 12600 19616 12628
rect 19475 12597 19487 12600
rect 19429 12591 19487 12597
rect 19610 12588 19616 12600
rect 19668 12588 19674 12640
rect 20073 12631 20131 12637
rect 20073 12597 20085 12631
rect 20119 12628 20131 12631
rect 21100 12628 21128 12668
rect 22833 12665 22845 12668
rect 22879 12665 22891 12699
rect 22833 12659 22891 12665
rect 20119 12600 21128 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 21913 12631 21971 12637
rect 21913 12628 21925 12631
rect 21876 12600 21925 12628
rect 21876 12588 21882 12600
rect 21913 12597 21925 12600
rect 21959 12597 21971 12631
rect 21913 12591 21971 12597
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 23106 12628 23112 12640
rect 22796 12600 23112 12628
rect 22796 12588 22802 12600
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 1104 12538 23460 12560
rect 1104 12486 8446 12538
rect 8498 12486 8510 12538
rect 8562 12486 8574 12538
rect 8626 12486 8638 12538
rect 8690 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 23460 12538
rect 1104 12464 23460 12486
rect 3418 12424 3424 12436
rect 3379 12396 3424 12424
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5316 12396 5457 12424
rect 5316 12384 5322 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5445 12387 5503 12393
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6328 12396 6929 12424
rect 6328 12384 6334 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 9088 12396 9321 12424
rect 9088 12384 9094 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 10042 12424 10048 12436
rect 9723 12396 10048 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10686 12424 10692 12436
rect 10192 12396 10692 12424
rect 10192 12384 10198 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11517 12427 11575 12433
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 12066 12424 12072 12436
rect 11563 12396 12072 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 14829 12427 14887 12433
rect 14829 12424 14841 12427
rect 14700 12396 14841 12424
rect 14700 12384 14706 12396
rect 14829 12393 14841 12396
rect 14875 12424 14887 12427
rect 15102 12424 15108 12436
rect 14875 12396 15108 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15562 12424 15568 12436
rect 15335 12396 15568 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16264 12396 16773 12424
rect 16264 12384 16270 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 16761 12387 16819 12393
rect 17052 12396 17233 12424
rect 2308 12359 2366 12365
rect 2308 12325 2320 12359
rect 2354 12356 2366 12359
rect 2774 12356 2780 12368
rect 2354 12328 2780 12356
rect 2354 12325 2366 12328
rect 2308 12319 2366 12325
rect 2774 12316 2780 12328
rect 2832 12356 2838 12368
rect 3326 12356 3332 12368
rect 2832 12328 3332 12356
rect 2832 12316 2838 12328
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 4332 12359 4390 12365
rect 4332 12325 4344 12359
rect 4378 12356 4390 12359
rect 4430 12356 4436 12368
rect 4378 12328 4436 12356
rect 4378 12325 4390 12328
rect 4332 12319 4390 12325
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 5804 12359 5862 12365
rect 5804 12325 5816 12359
rect 5850 12356 5862 12359
rect 6362 12356 6368 12368
rect 5850 12328 6368 12356
rect 5850 12325 5862 12328
rect 5804 12319 5862 12325
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 7276 12359 7334 12365
rect 7276 12325 7288 12359
rect 7322 12356 7334 12359
rect 8294 12356 8300 12368
rect 7322 12328 8300 12356
rect 7322 12325 7334 12328
rect 7276 12319 7334 12325
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 13357 12359 13415 12365
rect 13357 12356 13369 12359
rect 9508 12328 13369 12356
rect 4062 12288 4068 12300
rect 3975 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12288 4126 12300
rect 5537 12291 5595 12297
rect 5537 12288 5549 12291
rect 4120 12260 5549 12288
rect 4120 12248 4126 12260
rect 5537 12257 5549 12260
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 9508 12297 9536 12328
rect 13357 12325 13369 12328
rect 13403 12356 13415 12359
rect 13403 12328 14412 12356
rect 13403 12325 13415 12328
rect 13357 12319 13415 12325
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8260 12260 8861 12288
rect 8260 12248 8266 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 9493 12251 9551 12257
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10404 12291 10462 12297
rect 10404 12257 10416 12291
rect 10450 12288 10462 12291
rect 11514 12288 11520 12300
rect 10450 12260 11520 12288
rect 10450 12257 10462 12260
rect 10404 12251 10462 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 13716 12291 13774 12297
rect 13716 12257 13728 12291
rect 13762 12288 13774 12291
rect 14274 12288 14280 12300
rect 13762 12260 14280 12288
rect 13762 12257 13774 12260
rect 13716 12251 13774 12257
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6972 12192 7021 12220
rect 6972 12180 6978 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 7009 12183 7067 12189
rect 8404 12192 8953 12220
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 8404 12161 8432 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9398 12220 9404 12232
rect 9171 12192 9404 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 11624 12220 11652 12251
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 14384 12288 14412 12328
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 15580 12356 15608 12384
rect 16666 12356 16672 12368
rect 15068 12328 15516 12356
rect 15580 12328 16672 12356
rect 15068 12316 15074 12328
rect 15488 12297 15516 12328
rect 16666 12316 16672 12328
rect 16724 12316 16730 12368
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14384 12260 15117 12288
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16482 12288 16488 12300
rect 15979 12260 16488 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 17052 12288 17080 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 17221 12387 17279 12393
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 17368 12396 17601 12424
rect 17368 12384 17374 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 17589 12387 17647 12393
rect 23014 12384 23020 12436
rect 23072 12424 23078 12436
rect 23072 12396 23244 12424
rect 23072 12384 23078 12396
rect 23216 12368 23244 12396
rect 17126 12316 17132 12368
rect 17184 12356 17190 12368
rect 17681 12359 17739 12365
rect 17681 12356 17693 12359
rect 17184 12328 17693 12356
rect 17184 12316 17190 12328
rect 17681 12325 17693 12328
rect 17727 12325 17739 12359
rect 20438 12356 20444 12368
rect 20399 12328 20444 12356
rect 17681 12319 17739 12325
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 20990 12316 20996 12368
rect 21048 12356 21054 12368
rect 21422 12359 21480 12365
rect 21422 12356 21434 12359
rect 21048 12328 21434 12356
rect 21048 12316 21054 12328
rect 21422 12325 21434 12328
rect 21468 12356 21480 12359
rect 21818 12356 21824 12368
rect 21468 12328 21824 12356
rect 21468 12325 21480 12328
rect 21422 12319 21480 12325
rect 21818 12316 21824 12328
rect 21876 12316 21882 12368
rect 23198 12316 23204 12368
rect 23256 12316 23262 12368
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 17052 12260 18613 12288
rect 18601 12257 18613 12260
rect 18647 12288 18659 12291
rect 19242 12288 19248 12300
rect 18647 12260 19248 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19426 12288 19432 12300
rect 19387 12260 19432 12288
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 22922 12288 22928 12300
rect 20395 12260 22928 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 11532 12192 11652 12220
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 8352 12124 8401 12152
rect 8352 12112 8358 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 8389 12115 8447 12121
rect 8481 12155 8539 12161
rect 8481 12121 8493 12155
rect 8527 12152 8539 12155
rect 9766 12152 9772 12164
rect 8527 12124 9772 12152
rect 8527 12121 8539 12124
rect 8481 12115 8539 12121
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 11532 12084 11560 12192
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 12986 12220 12992 12232
rect 12676 12192 12992 12220
rect 12676 12180 12682 12192
rect 12986 12180 12992 12192
rect 13044 12220 13050 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13044 12192 13461 12220
rect 13044 12180 13050 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 15654 12180 15660 12232
rect 15712 12220 15718 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15712 12192 16037 12220
rect 15712 12180 15718 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 16853 12223 16911 12229
rect 16172 12192 16217 12220
rect 16172 12180 16178 12192
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17770 12220 17776 12232
rect 17083 12192 17776 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 14921 12155 14979 12161
rect 14921 12121 14933 12155
rect 14967 12152 14979 12155
rect 15378 12152 15384 12164
rect 14967 12124 15384 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 16868 12152 16896 12183
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18230 12220 18236 12232
rect 18012 12192 18236 12220
rect 18012 12180 18018 12192
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18708 12152 18736 12183
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 19518 12220 19524 12232
rect 18840 12192 18885 12220
rect 19479 12192 19524 12220
rect 18840 12180 18846 12192
rect 19518 12180 19524 12192
rect 19576 12180 19582 12232
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 20530 12220 20536 12232
rect 19668 12192 19713 12220
rect 20491 12192 20536 12220
rect 19668 12180 19674 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 20898 12180 20904 12232
rect 20956 12220 20962 12232
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 20956 12192 21189 12220
rect 20956 12180 20962 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 15528 12124 16896 12152
rect 17144 12124 18736 12152
rect 15528 12112 15534 12124
rect 17144 12096 17172 12124
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 19628 12152 19656 12180
rect 19392 12124 19656 12152
rect 19392 12112 19398 12124
rect 15562 12084 15568 12096
rect 3200 12056 11560 12084
rect 15523 12056 15568 12084
rect 3200 12044 3206 12056
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 17126 12084 17132 12096
rect 16439 12056 17132 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 18104 12056 18245 12084
rect 18104 12044 18110 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19061 12087 19119 12093
rect 19061 12084 19073 12087
rect 19024 12056 19073 12084
rect 19024 12044 19030 12056
rect 19061 12053 19073 12056
rect 19107 12053 19119 12087
rect 19978 12084 19984 12096
rect 19939 12056 19984 12084
rect 19061 12047 19119 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 22557 12087 22615 12093
rect 22557 12053 22569 12087
rect 22603 12084 22615 12087
rect 22646 12084 22652 12096
rect 22603 12056 22652 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 1104 11994 23460 12016
rect 1104 11942 4714 11994
rect 4766 11942 4778 11994
rect 4830 11942 4842 11994
rect 4894 11942 4906 11994
rect 4958 11942 12178 11994
rect 12230 11942 12242 11994
rect 12294 11942 12306 11994
rect 12358 11942 12370 11994
rect 12422 11942 19642 11994
rect 19694 11942 19706 11994
rect 19758 11942 19770 11994
rect 19822 11942 19834 11994
rect 19886 11942 23460 11994
rect 1104 11920 23460 11942
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4488 11852 4537 11880
rect 4488 11840 4494 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 4525 11843 4583 11849
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 8754 11880 8760 11892
rect 8435 11852 8760 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 10229 11883 10287 11889
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10318 11880 10324 11892
rect 10275 11852 10324 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 12618 11880 12624 11892
rect 12579 11852 12624 11880
rect 11793 11843 11851 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 14090 11880 14096 11892
rect 12820 11852 14096 11880
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 2096 11716 3157 11744
rect 2096 11704 2102 11716
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 10134 11744 10140 11756
rect 3145 11707 3203 11713
rect 9600 11716 10140 11744
rect 3412 11679 3470 11685
rect 3412 11645 3424 11679
rect 3458 11676 3470 11679
rect 3970 11676 3976 11688
rect 3458 11648 3976 11676
rect 3458 11645 3470 11648
rect 3412 11639 3470 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6972 11648 7021 11676
rect 6972 11636 6978 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9600 11676 9628 11716
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10192 11716 10425 11744
rect 10192 11704 10198 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 8619 11648 9628 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 12820 11685 12848 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14274 11880 14280 11892
rect 14235 11852 14280 11880
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15470 11880 15476 11892
rect 15431 11852 15476 11880
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 16482 11880 16488 11892
rect 16443 11852 16488 11880
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17773 11883 17831 11889
rect 17773 11849 17785 11883
rect 17819 11880 17831 11883
rect 19426 11880 19432 11892
rect 17819 11852 19432 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 22097 11883 22155 11889
rect 22097 11880 22109 11883
rect 20496 11852 22109 11880
rect 20496 11840 20502 11852
rect 22097 11849 22109 11852
rect 22143 11849 22155 11883
rect 22097 11843 22155 11849
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9732 11648 10057 11676
rect 9732 11636 9738 11648
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 14292 11676 14320 11840
rect 15378 11772 15384 11824
rect 15436 11812 15442 11824
rect 17954 11812 17960 11824
rect 15436 11784 17960 11812
rect 15436 11772 15442 11784
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 22002 11812 22008 11824
rect 21963 11784 22008 11812
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15194 11744 15200 11756
rect 15059 11716 15200 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15194 11704 15200 11716
rect 15252 11744 15258 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 15252 11716 16221 11744
rect 15252 11704 15258 11716
rect 16209 11713 16221 11716
rect 16255 11744 16267 11747
rect 16390 11744 16396 11756
rect 16255 11716 16396 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16390 11704 16396 11716
rect 16448 11744 16454 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16448 11716 17049 11744
rect 16448 11704 16454 11716
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19300 11716 19564 11744
rect 19300 11704 19306 11716
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 12952 11648 12997 11676
rect 14292 11648 14749 11676
rect 12952 11636 12958 11648
rect 14737 11645 14749 11648
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 15562 11676 15568 11688
rect 15335 11648 15568 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 16114 11676 16120 11688
rect 15948 11648 16120 11676
rect 7276 11611 7334 11617
rect 7276 11577 7288 11611
rect 7322 11608 7334 11611
rect 8202 11608 8208 11620
rect 7322 11580 8208 11608
rect 7322 11577 7334 11580
rect 7276 11571 7334 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8840 11611 8898 11617
rect 8840 11577 8852 11611
rect 8886 11608 8898 11611
rect 9306 11608 9312 11620
rect 8886 11580 9312 11608
rect 8886 11577 8898 11580
rect 8840 11571 8898 11577
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 10680 11611 10738 11617
rect 10680 11577 10692 11611
rect 10726 11608 10738 11611
rect 11790 11608 11796 11620
rect 10726 11580 11796 11608
rect 10726 11577 10738 11580
rect 10680 11571 10738 11577
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 13164 11611 13222 11617
rect 13164 11577 13176 11611
rect 13210 11608 13222 11611
rect 14182 11608 14188 11620
rect 13210 11580 14188 11608
rect 13210 11577 13222 11580
rect 13164 11571 13222 11577
rect 14182 11568 14188 11580
rect 14240 11608 14246 11620
rect 14829 11611 14887 11617
rect 14829 11608 14841 11611
rect 14240 11580 14841 11608
rect 14240 11568 14246 11580
rect 14829 11577 14841 11580
rect 14875 11577 14887 11611
rect 14829 11571 14887 11577
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 15746 11608 15752 11620
rect 14976 11580 15752 11608
rect 14976 11568 14982 11580
rect 15746 11568 15752 11580
rect 15804 11608 15810 11620
rect 15948 11608 15976 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 17184 11648 17601 11676
rect 17184 11636 17190 11648
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 18012 11648 18061 11676
rect 18012 11636 18018 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 18316 11679 18374 11685
rect 18316 11645 18328 11679
rect 18362 11676 18374 11679
rect 19334 11676 19340 11688
rect 18362 11648 19340 11676
rect 18362 11645 18374 11648
rect 18316 11639 18374 11645
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 19536 11685 19564 11716
rect 19978 11704 19984 11756
rect 20036 11744 20042 11756
rect 20628 11747 20686 11753
rect 20628 11744 20640 11747
rect 20036 11716 20640 11744
rect 20036 11704 20042 11716
rect 20628 11713 20640 11716
rect 20674 11713 20686 11747
rect 20628 11707 20686 11713
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 22370 11744 22376 11756
rect 20772 11716 22376 11744
rect 20772 11704 20778 11716
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 22646 11744 22652 11756
rect 22607 11716 22652 11744
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 22922 11744 22928 11756
rect 22883 11716 22928 11744
rect 22922 11704 22928 11716
rect 22980 11704 22986 11756
rect 19521 11679 19579 11685
rect 19521 11645 19533 11679
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 20128 11648 20177 11676
rect 20128 11636 20134 11648
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 20488 11679 20546 11685
rect 20488 11676 20500 11679
rect 20312 11648 20500 11676
rect 20312 11636 20318 11648
rect 20488 11645 20500 11648
rect 20534 11645 20546 11679
rect 20488 11639 20546 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 22557 11679 22615 11685
rect 20947 11648 21680 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 15804 11580 15976 11608
rect 16025 11611 16083 11617
rect 15804 11568 15810 11580
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16390 11608 16396 11620
rect 16071 11580 16396 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 19981 11611 20039 11617
rect 19981 11608 19993 11611
rect 18748 11580 19993 11608
rect 18748 11568 18754 11580
rect 19981 11577 19993 11580
rect 20027 11608 20039 11611
rect 20272 11608 20300 11636
rect 21652 11620 21680 11648
rect 22557 11645 22569 11679
rect 22603 11676 22615 11679
rect 22738 11676 22744 11688
rect 22603 11648 22744 11676
rect 22603 11645 22615 11648
rect 22557 11639 22615 11645
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 20027 11580 20300 11608
rect 20027 11577 20039 11580
rect 19981 11571 20039 11577
rect 21634 11568 21640 11620
rect 21692 11608 21698 11620
rect 22465 11611 22523 11617
rect 22465 11608 22477 11611
rect 21692 11580 22477 11608
rect 21692 11568 21698 11580
rect 22465 11577 22477 11580
rect 22511 11577 22523 11611
rect 22465 11571 22523 11577
rect 9950 11540 9956 11552
rect 9911 11512 9956 11540
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 14550 11540 14556 11552
rect 14415 11512 14556 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16206 11540 16212 11552
rect 16163 11512 16212 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17000 11512 17045 11540
rect 17000 11500 17006 11512
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19116 11512 19441 11540
rect 19116 11500 19122 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 19705 11543 19763 11549
rect 19705 11509 19717 11543
rect 19751 11540 19763 11543
rect 19886 11540 19892 11552
rect 19751 11512 19892 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 23460 11472
rect 1104 11398 8446 11450
rect 8498 11398 8510 11450
rect 8562 11398 8574 11450
rect 8626 11398 8638 11450
rect 8690 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 23460 11450
rect 1104 11376 23460 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 8202 11336 8208 11348
rect 2832 11308 2877 11336
rect 8163 11308 8208 11336
rect 2832 11296 2838 11308
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 10042 11336 10048 11348
rect 8855 11308 10048 11336
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 1642 11271 1700 11277
rect 1642 11268 1654 11271
rect 1452 11240 1654 11268
rect 1452 11228 1458 11240
rect 1642 11237 1654 11240
rect 1688 11237 1700 11271
rect 1642 11231 1700 11237
rect 7092 11271 7150 11277
rect 7092 11237 7104 11271
rect 7138 11268 7150 11271
rect 8294 11268 8300 11280
rect 7138 11240 8300 11268
rect 7138 11237 7150 11240
rect 7092 11231 7150 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 2038 11200 2044 11212
rect 1412 11172 2044 11200
rect 1412 11141 1440 11172
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11200 6883 11203
rect 6914 11200 6920 11212
rect 6871 11172 6920 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 8662 11200 8668 11212
rect 8623 11172 8668 11200
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 8754 11132 8760 11144
rect 8715 11104 8760 11132
rect 1397 11095 1455 11101
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 8855 11141 8883 11308
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10134 11296 10140 11348
rect 10192 11296 10198 11348
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 11701 11339 11759 11345
rect 11701 11336 11713 11339
rect 11572 11308 11713 11336
rect 11572 11296 11578 11308
rect 11701 11305 11713 11308
rect 11747 11305 11759 11339
rect 11701 11299 11759 11305
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 16761 11339 16819 11345
rect 11848 11308 11893 11336
rect 11848 11296 11854 11308
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 20714 11336 20720 11348
rect 18892 11308 20720 11336
rect 10152 11268 10180 11296
rect 13998 11268 14004 11280
rect 9876 11240 10180 11268
rect 12820 11240 14004 11268
rect 9030 11160 9036 11212
rect 9088 11200 9094 11212
rect 9876 11209 9904 11240
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9088 11172 9321 11200
rect 9088 11160 9094 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 10128 11203 10186 11209
rect 10128 11169 10140 11203
rect 10174 11200 10186 11203
rect 10686 11200 10692 11212
rect 10174 11172 10692 11200
rect 10174 11169 10186 11172
rect 10128 11163 10186 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 12820 11209 12848 11240
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 17396 11271 17454 11277
rect 17396 11237 17408 11271
rect 17442 11268 17454 11271
rect 18892 11268 18920 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 20901 11339 20959 11345
rect 20901 11305 20913 11339
rect 20947 11336 20959 11339
rect 22462 11336 22468 11348
rect 20947 11308 22468 11336
rect 20947 11305 20959 11308
rect 20901 11299 20959 11305
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 19058 11277 19064 11280
rect 19052 11268 19064 11277
rect 17442 11240 18920 11268
rect 19019 11240 19064 11268
rect 17442 11237 17454 11240
rect 17396 11231 17454 11237
rect 19052 11231 19064 11240
rect 19058 11228 19064 11231
rect 19116 11228 19122 11280
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 20257 11271 20315 11277
rect 20257 11268 20269 11271
rect 19392 11240 20269 11268
rect 19392 11228 19398 11240
rect 20257 11237 20269 11240
rect 20303 11237 20315 11271
rect 21358 11268 21364 11280
rect 21271 11240 21364 11268
rect 20257 11231 20315 11237
rect 21358 11228 21364 11240
rect 21416 11268 21422 11280
rect 21634 11268 21640 11280
rect 21416 11240 21640 11268
rect 21416 11228 21422 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 21996 11271 22054 11277
rect 21996 11237 22008 11271
rect 22042 11268 22054 11271
rect 22646 11268 22652 11280
rect 22042 11240 22652 11268
rect 22042 11237 22054 11240
rect 21996 11231 22054 11237
rect 22646 11228 22652 11240
rect 22704 11228 22710 11280
rect 12805 11203 12863 11209
rect 12805 11169 12817 11203
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 13164 11203 13222 11209
rect 13164 11169 13176 11203
rect 13210 11200 13222 11203
rect 14090 11200 14096 11212
rect 13210 11172 14096 11200
rect 13210 11169 13222 11172
rect 13164 11163 13222 11169
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14332 11172 14749 11200
rect 14332 11160 14338 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 15160 11172 15393 11200
rect 15160 11160 15166 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15648 11203 15706 11209
rect 15648 11169 15660 11203
rect 15694 11200 15706 11203
rect 16390 11200 16396 11212
rect 15694 11172 16396 11200
rect 15694 11169 15706 11172
rect 15648 11163 15706 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17954 11200 17960 11212
rect 17175 11172 17960 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17954 11160 17960 11172
rect 18012 11200 18018 11212
rect 18785 11203 18843 11209
rect 18785 11200 18797 11203
rect 18012 11172 18797 11200
rect 18012 11160 18018 11172
rect 18785 11169 18797 11172
rect 18831 11169 18843 11203
rect 18785 11163 18843 11169
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 19944 11172 21281 11200
rect 19944 11160 19950 11172
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 21450 11160 21456 11212
rect 21508 11200 21514 11212
rect 21729 11203 21787 11209
rect 21729 11200 21741 11203
rect 21508 11172 21741 11200
rect 21508 11160 21514 11172
rect 21729 11169 21741 11172
rect 21775 11169 21787 11203
rect 21729 11163 21787 11169
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 9766 11132 9772 11144
rect 8849 11095 8907 11101
rect 8956 11104 9772 11132
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 8956 11064 8984 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10962 11132 10968 11144
rect 10875 11104 10968 11132
rect 9122 11064 9128 11076
rect 8343 11036 8984 11064
rect 9035 11036 9128 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 9122 11024 9128 11036
rect 9180 11064 9186 11076
rect 9674 11064 9680 11076
rect 9180 11036 9680 11064
rect 9180 11024 9186 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 10888 10996 10916 11104
rect 10962 11092 10968 11104
rect 11020 11132 11026 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11020 11104 11897 11132
rect 11020 11092 11026 11104
rect 11885 11101 11897 11104
rect 11931 11132 11943 11135
rect 12526 11132 12532 11144
rect 11931 11104 12532 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12894 11132 12900 11144
rect 12855 11104 12900 11132
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 14108 11132 14136 11160
rect 14829 11135 14887 11141
rect 14829 11132 14841 11135
rect 14108 11104 14841 11132
rect 14829 11101 14841 11104
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11132 15071 11135
rect 15194 11132 15200 11144
rect 15059 11104 15200 11132
rect 15059 11101 15071 11104
rect 15013 11095 15071 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 21634 11132 21640 11144
rect 21591 11104 21640 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 12621 11067 12679 11073
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 12912 11064 12940 11092
rect 14274 11064 14280 11076
rect 12667 11036 12940 11064
rect 14235 11036 14280 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 14274 11024 14280 11036
rect 14332 11024 14338 11076
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 18380 11036 18521 11064
rect 18380 11024 18386 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 18690 11064 18696 11076
rect 18651 11036 18696 11064
rect 18509 11027 18567 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 20530 11064 20536 11076
rect 20312 11036 20536 11064
rect 20312 11024 20318 11036
rect 20530 11024 20536 11036
rect 20588 11064 20594 11076
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 20588 11036 21772 11064
rect 20588 11024 20594 11036
rect 10100 10968 10916 10996
rect 10100 10956 10106 10968
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11241 10999 11299 11005
rect 11241 10996 11253 10999
rect 11112 10968 11253 10996
rect 11112 10956 11118 10968
rect 11241 10965 11253 10968
rect 11287 10965 11299 10999
rect 11241 10959 11299 10965
rect 14366 10956 14372 11008
rect 14424 10996 14430 11008
rect 14424 10968 14469 10996
rect 14424 10956 14430 10968
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 19426 10996 19432 11008
rect 14700 10968 19432 10996
rect 14700 10956 14706 10968
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 20162 10996 20168 11008
rect 20123 10968 20168 10996
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 21744 10996 21772 11036
rect 22664 11036 23121 11064
rect 22664 10996 22692 11036
rect 23109 11033 23121 11036
rect 23155 11033 23167 11067
rect 23109 11027 23167 11033
rect 21744 10968 22692 10996
rect 1104 10906 23460 10928
rect 1104 10854 4714 10906
rect 4766 10854 4778 10906
rect 4830 10854 4842 10906
rect 4894 10854 4906 10906
rect 4958 10854 12178 10906
rect 12230 10854 12242 10906
rect 12294 10854 12306 10906
rect 12358 10854 12370 10906
rect 12422 10854 19642 10906
rect 19694 10854 19706 10906
rect 19758 10854 19770 10906
rect 19822 10854 19834 10906
rect 19886 10854 23460 10906
rect 1104 10832 23460 10854
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8662 10792 8668 10804
rect 8352 10764 8668 10792
rect 8352 10752 8358 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 10686 10792 10692 10804
rect 10647 10764 10692 10792
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11848 10764 12173 10792
rect 11848 10752 11854 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 14090 10792 14096 10804
rect 14051 10764 14096 10792
rect 12161 10755 12219 10761
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 14458 10792 14464 10804
rect 14231 10764 14464 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 16390 10792 16396 10804
rect 16351 10764 16396 10792
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 20070 10792 20076 10804
rect 18279 10764 19288 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6972 10628 7297 10656
rect 6972 10616 6978 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14424 10628 14657 10656
rect 14424 10616 14430 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 14918 10656 14924 10668
rect 14875 10628 14924 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 19058 10656 19064 10668
rect 19019 10628 19064 10656
rect 19058 10616 19064 10628
rect 19116 10616 19122 10668
rect 7552 10591 7610 10597
rect 7552 10557 7564 10591
rect 7598 10588 7610 10591
rect 8754 10588 8760 10600
rect 7598 10560 8760 10588
rect 7598 10557 7610 10560
rect 7552 10551 7610 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9576 10591 9634 10597
rect 9576 10557 9588 10591
rect 9622 10588 9634 10591
rect 9950 10588 9956 10600
rect 9622 10560 9956 10588
rect 9622 10557 9634 10560
rect 9576 10551 9634 10557
rect 9324 10520 9352 10551
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 11054 10597 11060 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10192 10560 10793 10588
rect 10192 10548 10198 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 11048 10588 11060 10597
rect 11015 10560 11060 10588
rect 10781 10551 10839 10557
rect 11048 10551 11060 10560
rect 11054 10548 11060 10551
rect 11112 10548 11118 10600
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 12802 10588 12808 10600
rect 12759 10560 12808 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 14550 10588 14556 10600
rect 14511 10560 14556 10588
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15102 10588 15108 10600
rect 15059 10560 15108 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 16482 10588 16488 10600
rect 16443 10560 16488 10588
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18966 10588 18972 10600
rect 18927 10560 18972 10588
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 19260 10588 19288 10764
rect 19444 10764 20076 10792
rect 19444 10668 19472 10764
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 21269 10795 21327 10801
rect 21269 10761 21281 10795
rect 21315 10792 21327 10795
rect 21358 10792 21364 10804
rect 21315 10764 21364 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22428 10764 22753 10792
rect 22428 10752 22434 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 19426 10656 19432 10668
rect 19339 10628 19432 10656
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19978 10665 19984 10668
rect 19935 10659 19984 10665
rect 19935 10625 19947 10659
rect 19981 10625 19984 10659
rect 19935 10619 19984 10625
rect 19978 10616 19984 10619
rect 20036 10616 20042 10668
rect 19518 10588 19524 10600
rect 19260 10560 19524 10588
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 20128 10560 20177 10588
rect 20128 10548 20134 10560
rect 20165 10557 20177 10560
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 20898 10548 20904 10600
rect 20956 10588 20962 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 20956 10560 21373 10588
rect 20956 10548 20962 10560
rect 21361 10557 21373 10560
rect 21407 10588 21419 10591
rect 21450 10588 21456 10600
rect 21407 10560 21456 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 21450 10548 21456 10560
rect 21508 10548 21514 10600
rect 10152 10520 10180 10548
rect 9324 10492 10180 10520
rect 12980 10523 13038 10529
rect 12980 10489 12992 10523
rect 13026 10520 13038 10523
rect 15280 10523 15338 10529
rect 13026 10492 15240 10520
rect 13026 10489 13038 10492
rect 12980 10483 13038 10489
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 15212 10452 15240 10492
rect 15280 10489 15292 10523
rect 15326 10520 15338 10523
rect 16206 10520 16212 10532
rect 15326 10492 16212 10520
rect 15326 10489 15338 10492
rect 15280 10483 15338 10489
rect 16206 10480 16212 10492
rect 16264 10520 16270 10532
rect 16390 10520 16396 10532
rect 16264 10492 16396 10520
rect 16264 10480 16270 10492
rect 16390 10480 16396 10492
rect 16448 10480 16454 10532
rect 16752 10523 16810 10529
rect 16752 10489 16764 10523
rect 16798 10520 16810 10523
rect 16942 10520 16948 10532
rect 16798 10492 16948 10520
rect 16798 10489 16810 10492
rect 16752 10483 16810 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 17034 10480 17040 10532
rect 17092 10520 17098 10532
rect 18877 10523 18935 10529
rect 17092 10492 18552 10520
rect 17092 10480 17098 10492
rect 16850 10452 16856 10464
rect 15212 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10452 16914 10464
rect 18524 10461 18552 10492
rect 18877 10489 18889 10523
rect 18923 10520 18935 10523
rect 19334 10520 19340 10532
rect 18923 10492 19340 10520
rect 18923 10489 18935 10492
rect 18877 10483 18935 10489
rect 19334 10480 19340 10492
rect 19392 10480 19398 10532
rect 21634 10529 21640 10532
rect 21628 10520 21640 10529
rect 21595 10492 21640 10520
rect 21628 10483 21640 10492
rect 21634 10480 21640 10483
rect 21692 10480 21698 10532
rect 17865 10455 17923 10461
rect 17865 10452 17877 10455
rect 16908 10424 17877 10452
rect 16908 10412 16914 10424
rect 17865 10421 17877 10424
rect 17911 10421 17923 10455
rect 17865 10415 17923 10421
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 18598 10452 18604 10464
rect 18555 10424 18604 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19895 10455 19953 10461
rect 19895 10452 19907 10455
rect 18748 10424 19907 10452
rect 18748 10412 18754 10424
rect 19895 10421 19907 10424
rect 19941 10421 19953 10455
rect 19895 10415 19953 10421
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 22888 10424 22933 10452
rect 22888 10412 22894 10424
rect 1104 10362 23460 10384
rect 1104 10310 8446 10362
rect 8498 10310 8510 10362
rect 8562 10310 8574 10362
rect 8626 10310 8638 10362
rect 8690 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 23460 10362
rect 1104 10288 23460 10310
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 9858 10248 9864 10260
rect 9723 10220 9864 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 10008 10220 10057 10248
rect 10008 10208 10014 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 10505 10251 10563 10257
rect 10505 10248 10517 10251
rect 10468 10220 10517 10248
rect 10468 10208 10474 10220
rect 10505 10217 10517 10220
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11054 10248 11060 10260
rect 10919 10220 11060 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 14369 10251 14427 10257
rect 14369 10217 14381 10251
rect 14415 10248 14427 10251
rect 19337 10251 19395 10257
rect 14415 10220 17632 10248
rect 14415 10217 14427 10220
rect 14369 10211 14427 10217
rect 8196 10183 8254 10189
rect 8196 10149 8208 10183
rect 8242 10180 8254 10183
rect 8294 10180 8300 10192
rect 8242 10152 8300 10180
rect 8242 10149 8254 10152
rect 8196 10143 8254 10149
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 9324 10180 9352 10208
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 9324 10152 10149 10180
rect 10137 10149 10149 10152
rect 10183 10149 10195 10183
rect 10137 10143 10195 10149
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 10965 10183 11023 10189
rect 10965 10180 10977 10183
rect 10744 10152 10977 10180
rect 10744 10140 10750 10152
rect 10965 10149 10977 10152
rect 11011 10149 11023 10183
rect 10965 10143 11023 10149
rect 13164 10183 13222 10189
rect 13164 10149 13176 10183
rect 13210 10180 13222 10183
rect 14274 10180 14280 10192
rect 13210 10152 14280 10180
rect 13210 10149 13222 10152
rect 13164 10143 13222 10149
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 14737 10183 14795 10189
rect 14737 10149 14749 10183
rect 14783 10180 14795 10183
rect 17221 10183 17279 10189
rect 17221 10180 17233 10183
rect 14783 10152 17233 10180
rect 14783 10149 14795 10152
rect 14737 10143 14795 10149
rect 17221 10149 17233 10152
rect 17267 10149 17279 10183
rect 17221 10143 17279 10149
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 9582 10112 9588 10124
rect 7975 10084 9588 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12483 10084 12541 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12529 10081 12541 10084
rect 12575 10112 12587 10115
rect 14642 10112 14648 10124
rect 12575 10084 14648 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 14829 10115 14887 10121
rect 14829 10081 14841 10115
rect 14875 10112 14887 10115
rect 15378 10112 15384 10124
rect 14875 10084 15384 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15562 10121 15568 10124
rect 15556 10112 15568 10121
rect 15523 10084 15568 10112
rect 15556 10075 15568 10084
rect 15562 10072 15568 10075
rect 15620 10072 15626 10124
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 16724 10084 17509 10112
rect 16724 10072 16730 10084
rect 17420 10056 17448 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 17604 10112 17632 10220
rect 19337 10217 19349 10251
rect 19383 10248 19395 10251
rect 19981 10251 20039 10257
rect 19981 10248 19993 10251
rect 19383 10220 19993 10248
rect 19383 10217 19395 10220
rect 19337 10211 19395 10217
rect 19981 10217 19993 10220
rect 20027 10248 20039 10251
rect 20070 10248 20076 10260
rect 20027 10220 20076 10248
rect 20027 10217 20039 10220
rect 19981 10211 20039 10217
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 21692 10220 22293 10248
rect 21692 10208 21698 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 22741 10251 22799 10257
rect 22741 10217 22753 10251
rect 22787 10248 22799 10251
rect 22830 10248 22836 10260
rect 22787 10220 22836 10248
rect 22787 10217 22799 10220
rect 22741 10211 22799 10217
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 18966 10140 18972 10192
rect 19024 10180 19030 10192
rect 19426 10180 19432 10192
rect 19024 10152 19432 10180
rect 19024 10140 19030 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 17604 10084 18003 10112
rect 17497 10075 17555 10081
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 10100 10016 10241 10044
rect 10100 10004 10106 10016
rect 10229 10013 10241 10016
rect 10275 10044 10287 10047
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 10275 10016 11069 10044
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 11057 10013 11069 10016
rect 11103 10013 11115 10047
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 11057 10007 11115 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 15010 10044 15016 10056
rect 14971 10016 15016 10044
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15160 10016 15301 10044
rect 15160 10004 15166 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 17092 10016 17141 10044
rect 17092 10004 17098 10016
rect 17129 10013 17141 10016
rect 17175 10044 17187 10047
rect 17175 10016 17356 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 14240 9948 14289 9976
rect 14240 9936 14246 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14277 9939 14335 9945
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16448 9948 16681 9976
rect 16448 9936 16454 9948
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16669 9939 16727 9945
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17328 9976 17356 10016
rect 17402 10004 17408 10056
rect 17460 10004 17466 10056
rect 17975 10053 18003 10084
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 19889 10115 19947 10121
rect 19889 10112 19901 10115
rect 18656 10084 19901 10112
rect 18656 10072 18662 10084
rect 19889 10081 19901 10084
rect 19935 10081 19947 10115
rect 19889 10075 19947 10081
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 20898 10112 20904 10124
rect 20772 10084 20904 10112
rect 20772 10072 20778 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21174 10121 21180 10124
rect 21168 10075 21180 10121
rect 21232 10112 21238 10124
rect 21232 10084 21268 10112
rect 21174 10072 21180 10075
rect 21232 10072 21238 10084
rect 22462 10072 22468 10124
rect 22520 10112 22526 10124
rect 22833 10115 22891 10121
rect 22833 10112 22845 10115
rect 22520 10084 22845 10112
rect 22520 10072 22526 10084
rect 22833 10081 22845 10084
rect 22879 10081 22891 10115
rect 22833 10075 22891 10081
rect 17820 10047 17878 10053
rect 17820 10044 17832 10047
rect 17512 10016 17832 10044
rect 17512 9976 17540 10016
rect 17820 10013 17832 10016
rect 17866 10013 17878 10047
rect 17820 10007 17878 10013
rect 17960 10047 18018 10053
rect 17960 10013 17972 10047
rect 18006 10013 18018 10047
rect 18230 10044 18236 10056
rect 18191 10016 18236 10044
rect 17960 10007 18018 10013
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 20162 10044 20168 10056
rect 20123 10016 20168 10044
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20806 10044 20812 10056
rect 20579 10016 20812 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 22925 10047 22983 10053
rect 22925 10044 22937 10047
rect 22428 10016 22937 10044
rect 22428 10004 22434 10016
rect 22925 10013 22937 10016
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 16908 9948 17172 9976
rect 17328 9948 17540 9976
rect 16908 9936 16914 9948
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 12124 9880 12725 9908
rect 12124 9868 12130 9880
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 17144 9908 17172 9948
rect 20070 9936 20076 9988
rect 20128 9976 20134 9988
rect 20622 9976 20628 9988
rect 20128 9948 20628 9976
rect 20128 9936 20134 9948
rect 20622 9936 20628 9948
rect 20680 9936 20686 9988
rect 18230 9908 18236 9920
rect 17144 9880 18236 9908
rect 12713 9871 12771 9877
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 19521 9911 19579 9917
rect 19521 9877 19533 9911
rect 19567 9908 19579 9911
rect 21542 9908 21548 9920
rect 19567 9880 21548 9908
rect 19567 9877 19579 9880
rect 19521 9871 19579 9877
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 22373 9911 22431 9917
rect 22373 9877 22385 9911
rect 22419 9908 22431 9911
rect 23106 9908 23112 9920
rect 22419 9880 23112 9908
rect 22419 9877 22431 9880
rect 22373 9871 22431 9877
rect 23106 9868 23112 9880
rect 23164 9868 23170 9920
rect 1104 9818 23460 9840
rect 1104 9766 4714 9818
rect 4766 9766 4778 9818
rect 4830 9766 4842 9818
rect 4894 9766 4906 9818
rect 4958 9766 12178 9818
rect 12230 9766 12242 9818
rect 12294 9766 12306 9818
rect 12358 9766 12370 9818
rect 12422 9766 19642 9818
rect 19694 9766 19706 9818
rect 19758 9766 19770 9818
rect 19822 9766 19834 9818
rect 19886 9766 23460 9818
rect 1104 9744 23460 9766
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18230 9704 18236 9716
rect 18012 9676 18236 9704
rect 18012 9664 18018 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 21174 9704 21180 9716
rect 21135 9676 21180 9704
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 23569 9707 23627 9713
rect 23569 9704 23581 9707
rect 22756 9676 23060 9704
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 9766 9636 9772 9648
rect 9723 9608 9772 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 9766 9596 9772 9608
rect 9824 9636 9830 9648
rect 11698 9636 11704 9648
rect 9824 9608 11704 9636
rect 9824 9596 9830 9608
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 15378 9596 15384 9648
rect 15436 9636 15442 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 15436 9608 16313 9636
rect 15436 9596 15442 9608
rect 16301 9605 16313 9608
rect 16347 9605 16359 9639
rect 18046 9636 18052 9648
rect 16301 9599 16359 9605
rect 16868 9608 18052 9636
rect 12066 9568 12072 9580
rect 12027 9540 12072 9568
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 16868 9568 16896 9608
rect 17696 9577 17724 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 19426 9636 19432 9648
rect 19387 9608 19432 9636
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 15764 9540 16896 9568
rect 16945 9571 17003 9577
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9732 9472 9873 9500
rect 9732 9460 9738 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12986 9500 12992 9512
rect 12483 9472 12992 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13872 9472 14197 9500
rect 13872 9460 13878 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14452 9503 14510 9509
rect 14452 9469 14464 9503
rect 14498 9500 14510 9503
rect 15764 9500 15792 9540
rect 16945 9537 16957 9571
rect 16991 9568 17003 9571
rect 17681 9571 17739 9577
rect 16991 9540 17172 9568
rect 16991 9537 17003 9540
rect 16945 9531 17003 9537
rect 14498 9472 15792 9500
rect 15841 9503 15899 9509
rect 14498 9469 14510 9472
rect 14452 9463 14510 9469
rect 15841 9469 15853 9503
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9500 16727 9503
rect 16850 9500 16856 9512
rect 16715 9472 16856 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 11885 9435 11943 9441
rect 11885 9432 11897 9435
rect 10928 9404 11897 9432
rect 10928 9392 10934 9404
rect 11885 9401 11897 9404
rect 11931 9401 11943 9435
rect 11885 9395 11943 9401
rect 12704 9435 12762 9441
rect 12704 9401 12716 9435
rect 12750 9432 12762 9435
rect 13170 9432 13176 9444
rect 12750 9404 13176 9432
rect 12750 9401 12762 9404
rect 12704 9395 12762 9401
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 15856 9432 15884 9463
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 17144 9500 17172 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 21192 9568 21220 9664
rect 21269 9639 21327 9645
rect 21269 9605 21281 9639
rect 21315 9636 21327 9639
rect 22646 9636 22652 9648
rect 21315 9608 22652 9636
rect 21315 9605 21327 9608
rect 21269 9599 21327 9605
rect 22646 9596 22652 9608
rect 22704 9636 22710 9648
rect 22756 9636 22784 9676
rect 22922 9636 22928 9648
rect 22704 9608 22784 9636
rect 22883 9608 22928 9636
rect 22704 9596 22710 9608
rect 22922 9596 22928 9608
rect 22980 9596 22986 9648
rect 23032 9636 23060 9676
rect 23492 9676 23581 9704
rect 23032 9608 23152 9636
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 17681 9531 17739 9537
rect 17788 9540 18184 9568
rect 21192 9540 21833 9568
rect 17788 9500 17816 9540
rect 17144 9472 17816 9500
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 18012 9472 18061 9500
rect 18012 9460 18018 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18156 9500 18184 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 22741 9571 22799 9577
rect 22741 9568 22753 9571
rect 21821 9531 21879 9537
rect 22296 9540 22753 9568
rect 18322 9509 18328 9512
rect 18316 9500 18328 9509
rect 18156 9472 18328 9500
rect 18049 9463 18107 9469
rect 18316 9463 18328 9472
rect 18322 9460 18328 9463
rect 18380 9460 18386 9512
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 18656 9472 19717 9500
rect 18656 9460 18662 9472
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 19843 9472 20760 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 15528 9404 15884 9432
rect 16761 9435 16819 9441
rect 15528 9392 15534 9404
rect 16761 9401 16773 9435
rect 16807 9432 16819 9435
rect 16942 9432 16948 9444
rect 16807 9404 16948 9432
rect 16807 9401 16819 9404
rect 16761 9395 16819 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 17144 9404 18276 9432
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 11606 9364 11612 9376
rect 11563 9336 11612 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 13538 9364 13544 9376
rect 12023 9336 13544 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 13538 9324 13544 9336
rect 13596 9364 13602 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13596 9336 13829 9364
rect 13596 9324 13602 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15436 9336 15577 9364
rect 15436 9324 15442 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16390 9364 16396 9376
rect 15712 9336 16396 9364
rect 15712 9324 15718 9336
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 17144 9373 17172 9404
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9333 17187 9367
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 17129 9327 17187 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 18248 9364 18276 9404
rect 18414 9392 18420 9444
rect 18472 9432 18478 9444
rect 19812 9432 19840 9463
rect 20732 9444 20760 9472
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 22296 9509 22324 9540
rect 22741 9537 22753 9540
rect 22787 9568 22799 9571
rect 23014 9568 23020 9580
rect 22787 9540 23020 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 21637 9503 21695 9509
rect 21637 9500 21649 9503
rect 20864 9472 21649 9500
rect 20864 9460 20870 9472
rect 21637 9469 21649 9472
rect 21683 9469 21695 9503
rect 21637 9463 21695 9469
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9469 22339 9503
rect 22281 9463 22339 9469
rect 18472 9404 19840 9432
rect 20064 9435 20122 9441
rect 18472 9392 18478 9404
rect 19444 9376 19472 9404
rect 20064 9401 20076 9435
rect 20110 9432 20122 9435
rect 20162 9432 20168 9444
rect 20110 9404 20168 9432
rect 20110 9401 20122 9404
rect 20064 9395 20122 9401
rect 20162 9392 20168 9404
rect 20220 9392 20226 9444
rect 20714 9392 20720 9444
rect 20772 9392 20778 9444
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 21729 9435 21787 9441
rect 21729 9432 21741 9435
rect 21600 9404 21741 9432
rect 21600 9392 21606 9404
rect 21729 9401 21741 9404
rect 21775 9401 21787 9435
rect 21729 9395 21787 9401
rect 19334 9364 19340 9376
rect 17644 9336 17689 9364
rect 18248 9336 19340 9364
rect 17644 9324 17650 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 19521 9367 19579 9373
rect 19521 9364 19533 9367
rect 19484 9336 19533 9364
rect 19484 9324 19490 9336
rect 19521 9333 19533 9336
rect 19567 9333 19579 9367
rect 19521 9327 19579 9333
rect 19794 9324 19800 9376
rect 19852 9364 19858 9376
rect 22465 9367 22523 9373
rect 22465 9364 22477 9367
rect 19852 9336 22477 9364
rect 19852 9324 19858 9336
rect 22465 9333 22477 9336
rect 22511 9333 22523 9367
rect 23014 9364 23020 9376
rect 22975 9336 23020 9364
rect 22465 9327 22523 9333
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 23124 9364 23152 9608
rect 23492 9432 23520 9676
rect 23569 9673 23581 9676
rect 23615 9673 23627 9707
rect 23569 9667 23627 9673
rect 23569 9571 23627 9577
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 23658 9568 23664 9580
rect 23615 9540 23664 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 23658 9432 23664 9444
rect 23492 9404 23664 9432
rect 23658 9392 23664 9404
rect 23716 9392 23722 9444
rect 23569 9367 23627 9373
rect 23569 9364 23581 9367
rect 23124 9336 23581 9364
rect 23569 9333 23581 9336
rect 23615 9333 23627 9367
rect 23569 9327 23627 9333
rect 1104 9274 23460 9296
rect 1104 9222 8446 9274
rect 8498 9222 8510 9274
rect 8562 9222 8574 9274
rect 8626 9222 8638 9274
rect 8690 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 23460 9274
rect 1104 9200 23460 9222
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 10928 9132 14657 9160
rect 10928 9120 10934 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 19794 9160 19800 9172
rect 15804 9132 19800 9160
rect 15804 9120 15810 9132
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 21545 9163 21603 9169
rect 21545 9129 21557 9163
rect 21591 9160 21603 9163
rect 21910 9160 21916 9172
rect 21591 9132 21916 9160
rect 21591 9129 21603 9132
rect 21545 9123 21603 9129
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 13538 9101 13544 9104
rect 13532 9092 13544 9101
rect 11808 9064 12940 9092
rect 13499 9064 13544 9092
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9640 8996 9689 9024
rect 9640 8984 9646 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9944 9027 10002 9033
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 10502 9024 10508 9036
rect 9990 8996 10508 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11514 9024 11520 9036
rect 11471 8996 11520 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11808 9033 11836 9064
rect 12912 9036 12940 9064
rect 13532 9055 13544 9064
rect 13538 9052 13544 9055
rect 13596 9052 13602 9104
rect 14016 9064 15148 9092
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 12060 9027 12118 9033
rect 12060 8993 12072 9027
rect 12106 9024 12118 9027
rect 12618 9024 12624 9036
rect 12106 8996 12624 9024
rect 12106 8993 12118 8996
rect 12060 8987 12118 8993
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 13265 9027 13323 9033
rect 13265 9024 13277 9027
rect 12952 8996 13277 9024
rect 12952 8984 12958 8996
rect 13265 8993 13277 8996
rect 13311 9024 13323 9027
rect 14016 9024 14044 9064
rect 15120 9036 15148 9064
rect 16758 9052 16764 9104
rect 16816 9092 16822 9104
rect 17304 9095 17362 9101
rect 16816 9064 17264 9092
rect 16816 9052 16822 9064
rect 14918 9024 14924 9036
rect 13311 8996 14044 9024
rect 14879 8996 14924 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 15102 8984 15108 9036
rect 15160 9024 15166 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15160 8996 15301 9024
rect 15160 8984 15166 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15545 9027 15603 9033
rect 15545 9024 15557 9027
rect 15289 8987 15347 8993
rect 15396 8996 15557 9024
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15396 8956 15424 8996
rect 15545 8993 15557 8996
rect 15591 8993 15603 9027
rect 15545 8987 15603 8993
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16448 8996 16957 9024
rect 16448 8984 16454 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 17236 9024 17264 9064
rect 17304 9061 17316 9095
rect 17350 9092 17362 9095
rect 17954 9092 17960 9104
rect 17350 9064 17960 9092
rect 17350 9061 17362 9064
rect 17304 9055 17362 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 19334 9052 19340 9104
rect 19392 9092 19398 9104
rect 23658 9092 23664 9104
rect 19392 9064 23664 9092
rect 19392 9052 19398 9064
rect 23658 9052 23664 9064
rect 23716 9052 23722 9104
rect 17862 9024 17868 9036
rect 17236 8996 17868 9024
rect 16945 8987 17003 8993
rect 17862 8984 17868 8996
rect 17920 9024 17926 9036
rect 18598 9024 18604 9036
rect 17920 8996 18604 9024
rect 17920 8984 17926 8996
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 18776 9027 18834 9033
rect 18776 8993 18788 9027
rect 18822 9024 18834 9027
rect 19518 9024 19524 9036
rect 18822 8996 19524 9024
rect 18822 8993 18834 8996
rect 18776 8987 18834 8993
rect 19518 8984 19524 8996
rect 19576 8984 19582 9036
rect 20346 9024 20352 9036
rect 20307 8996 20352 9024
rect 20346 8984 20352 8996
rect 20404 8984 20410 9036
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 20772 8996 21649 9024
rect 20772 8984 20778 8996
rect 21637 8993 21649 8996
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 21904 9027 21962 9033
rect 21904 8993 21916 9027
rect 21950 9024 21962 9027
rect 22462 9024 22468 9036
rect 21950 8996 22468 9024
rect 21950 8993 21962 8996
rect 21904 8987 21962 8993
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 15252 8928 15424 8956
rect 15252 8916 15258 8928
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16540 8928 17049 8956
rect 16540 8916 16546 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18288 8928 18521 8956
rect 18288 8916 18294 8928
rect 18509 8925 18521 8928
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20441 8959 20499 8965
rect 20441 8956 20453 8959
rect 19668 8928 20453 8956
rect 19668 8916 19674 8928
rect 20441 8925 20453 8928
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8925 20591 8959
rect 20533 8919 20591 8925
rect 14458 8848 14464 8900
rect 14516 8888 14522 8900
rect 19978 8888 19984 8900
rect 14516 8860 15332 8888
rect 14516 8848 14522 8860
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 12986 8820 12992 8832
rect 11655 8792 12992 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13170 8820 13176 8832
rect 13131 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14274 8820 14280 8832
rect 14056 8792 14280 8820
rect 14056 8780 14062 8792
rect 14274 8780 14280 8792
rect 14332 8820 14338 8832
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14332 8792 14749 8820
rect 14332 8780 14338 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 15102 8820 15108 8832
rect 15063 8792 15108 8820
rect 14737 8783 14795 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15304 8820 15332 8860
rect 16408 8860 17080 8888
rect 16408 8820 16436 8860
rect 16666 8820 16672 8832
rect 15304 8792 16436 8820
rect 16627 8792 16672 8820
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 17052 8820 17080 8860
rect 17972 8860 18552 8888
rect 19939 8860 19984 8888
rect 17972 8820 18000 8860
rect 16816 8792 16861 8820
rect 17052 8792 18000 8820
rect 16816 8780 16822 8792
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18417 8823 18475 8829
rect 18417 8820 18429 8823
rect 18104 8792 18429 8820
rect 18104 8780 18110 8792
rect 18417 8789 18429 8792
rect 18463 8789 18475 8823
rect 18524 8820 18552 8860
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 20548 8888 20576 8919
rect 20456 8860 20576 8888
rect 19889 8823 19947 8829
rect 19889 8820 19901 8823
rect 18524 8792 19901 8820
rect 18417 8783 18475 8789
rect 19889 8789 19901 8792
rect 19935 8820 19947 8823
rect 20456 8820 20484 8860
rect 19935 8792 20484 8820
rect 20993 8823 21051 8829
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20993 8789 21005 8823
rect 21039 8820 21051 8823
rect 21082 8820 21088 8832
rect 21039 8792 21088 8820
rect 21039 8789 21051 8792
rect 20993 8783 21051 8789
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 23017 8823 23075 8829
rect 23017 8820 23029 8823
rect 22336 8792 23029 8820
rect 22336 8780 22342 8792
rect 23017 8789 23029 8792
rect 23063 8789 23075 8823
rect 23017 8783 23075 8789
rect 1104 8730 23460 8752
rect 1104 8678 4714 8730
rect 4766 8678 4778 8730
rect 4830 8678 4842 8730
rect 4894 8678 4906 8730
rect 4958 8678 12178 8730
rect 12230 8678 12242 8730
rect 12294 8678 12306 8730
rect 12358 8678 12370 8730
rect 12422 8678 19642 8730
rect 19694 8678 19706 8730
rect 19758 8678 19770 8730
rect 19822 8678 19834 8730
rect 19886 8678 23460 8730
rect 1104 8656 23460 8678
rect 9582 8616 9588 8628
rect 9232 8588 9588 8616
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2866 8480 2872 8492
rect 2087 8452 2872 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 9232 8489 9260 8588
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10560 8588 10609 8616
rect 10560 8576 10566 8588
rect 10597 8585 10609 8588
rect 10643 8616 10655 8619
rect 11514 8616 11520 8628
rect 10643 8588 11192 8616
rect 11475 8588 11520 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 11164 8489 11192 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 12676 8588 13829 8616
rect 12676 8576 12682 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 13955 8588 14596 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 14568 8548 14596 8588
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 15562 8616 15568 8628
rect 14700 8588 15568 8616
rect 14700 8576 14706 8588
rect 15562 8576 15568 8588
rect 15620 8616 15626 8628
rect 16666 8616 16672 8628
rect 15620 8588 16672 8616
rect 15620 8576 15626 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 17129 8619 17187 8625
rect 17129 8585 17141 8619
rect 17175 8616 17187 8619
rect 17586 8616 17592 8628
rect 17175 8588 17592 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18748 8588 19472 8616
rect 18748 8576 18754 8588
rect 14568 8520 14688 8548
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11974 8480 11980 8492
rect 11379 8452 11980 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12158 8480 12164 8492
rect 12119 8452 12164 8480
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14660 8480 14688 8520
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 16632 8520 16957 8548
rect 16632 8508 16638 8520
rect 16945 8517 16957 8520
rect 16991 8548 17003 8551
rect 17034 8548 17040 8560
rect 16991 8520 17040 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 19444 8548 19472 8588
rect 19518 8576 19524 8628
rect 19576 8616 19582 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19576 8588 19901 8616
rect 19576 8576 19582 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22060 8588 22784 8616
rect 22060 8576 22066 8588
rect 19794 8548 19800 8560
rect 17552 8520 18092 8548
rect 19444 8520 19800 8548
rect 17552 8508 17558 8520
rect 15200 8483 15258 8489
rect 15200 8480 15212 8483
rect 14660 8452 15212 8480
rect 15200 8449 15212 8452
rect 15246 8449 15258 8483
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15200 8443 15258 8449
rect 15396 8452 16681 8480
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 2409 8415 2467 8421
rect 2409 8412 2421 8415
rect 1811 8384 2421 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2409 8381 2421 8384
rect 2455 8412 2467 8415
rect 7742 8412 7748 8424
rect 2455 8384 7748 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 9484 8415 9542 8421
rect 9484 8381 9496 8415
rect 9530 8412 9542 8415
rect 10870 8412 10876 8424
rect 9530 8384 10876 8412
rect 9530 8381 9542 8384
rect 9484 8375 9542 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11054 8412 11060 8424
rect 11015 8384 11060 8412
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11664 8384 11897 8412
rect 11664 8372 11670 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12704 8415 12762 8421
rect 12704 8381 12716 8415
rect 12750 8412 12762 8415
rect 14458 8412 14464 8424
rect 12750 8384 14464 8412
rect 12750 8381 12762 8384
rect 12704 8375 12762 8381
rect 11238 8344 11244 8356
rect 10704 8316 11244 8344
rect 10704 8285 10732 8316
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 12452 8344 12480 8375
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 14745 8415 14803 8421
rect 14745 8412 14757 8415
rect 14700 8384 14757 8412
rect 14700 8372 14706 8384
rect 14745 8381 14757 8384
rect 14791 8381 14803 8415
rect 15396 8412 15424 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17586 8480 17592 8492
rect 16908 8452 17592 8480
rect 16908 8440 16914 8452
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8480 17831 8483
rect 17954 8480 17960 8492
rect 17819 8452 17960 8480
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18064 8489 18092 8520
rect 19794 8508 19800 8520
rect 19852 8508 19858 8560
rect 21913 8551 21971 8557
rect 21913 8517 21925 8551
rect 21959 8548 21971 8551
rect 22370 8548 22376 8560
rect 21959 8520 22376 8548
rect 21959 8517 21971 8520
rect 21913 8511 21971 8517
rect 22370 8508 22376 8520
rect 22428 8508 22434 8560
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18288 8452 18521 8480
rect 18288 8440 18294 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 19702 8440 19708 8492
rect 19760 8480 19766 8492
rect 20530 8489 20536 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19760 8452 19993 8480
rect 19760 8440 19766 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20487 8483 20536 8489
rect 20487 8449 20499 8483
rect 20533 8449 20536 8483
rect 20487 8443 20536 8449
rect 20530 8440 20536 8443
rect 20588 8440 20594 8492
rect 22278 8480 22284 8492
rect 20640 8452 22284 8480
rect 14745 8375 14803 8381
rect 14844 8384 15424 8412
rect 15473 8415 15531 8421
rect 13814 8344 13820 8356
rect 12452 8316 13820 8344
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14277 8347 14335 8353
rect 14277 8313 14289 8347
rect 14323 8344 14335 8347
rect 14844 8344 14872 8384
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15562 8412 15568 8424
rect 15519 8384 15568 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15562 8372 15568 8384
rect 15620 8412 15626 8424
rect 18776 8415 18834 8421
rect 15620 8384 18552 8412
rect 15620 8372 15626 8384
rect 14323 8316 14872 8344
rect 14323 8313 14335 8316
rect 14277 8307 14335 8313
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 16448 8316 17509 8344
rect 16448 8304 16454 8316
rect 17497 8313 17509 8316
rect 17543 8313 17555 8347
rect 18524 8344 18552 8384
rect 18776 8381 18788 8415
rect 18822 8412 18834 8415
rect 20640 8412 20668 8452
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 22462 8480 22468 8492
rect 22423 8452 22468 8480
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 18822 8384 20668 8412
rect 18822 8381 18834 8384
rect 18776 8375 18834 8381
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 20772 8384 20817 8412
rect 20772 8372 20778 8384
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 22756 8421 22784 8588
rect 22741 8415 22799 8421
rect 21048 8384 21404 8412
rect 21048 8372 21054 8384
rect 19794 8344 19800 8356
rect 18524 8316 19800 8344
rect 17497 8307 17555 8313
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 21376 8344 21404 8384
rect 22741 8381 22753 8415
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 22281 8347 22339 8353
rect 22281 8344 22293 8347
rect 21376 8316 22293 8344
rect 22281 8313 22293 8316
rect 22327 8313 22339 8347
rect 22281 8307 22339 8313
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8245 10747 8279
rect 10689 8239 10747 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12032 8248 12077 8276
rect 12032 8236 12038 8248
rect 14366 8236 14372 8288
rect 14424 8276 14430 8288
rect 14424 8248 14469 8276
rect 14424 8236 14430 8248
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 15102 8276 15108 8288
rect 14700 8248 15108 8276
rect 14700 8236 14706 8248
rect 15102 8236 15108 8248
rect 15160 8276 15166 8288
rect 15203 8279 15261 8285
rect 15203 8276 15215 8279
rect 15160 8248 15215 8276
rect 15160 8236 15166 8248
rect 15203 8245 15215 8248
rect 15249 8276 15261 8279
rect 16482 8276 16488 8288
rect 15249 8248 16488 8276
rect 15249 8245 15261 8248
rect 15203 8239 15261 8245
rect 16482 8236 16488 8248
rect 16540 8236 16546 8288
rect 16577 8279 16635 8285
rect 16577 8245 16589 8279
rect 16623 8276 16635 8279
rect 16758 8276 16764 8288
rect 16623 8248 16764 8276
rect 16623 8245 16635 8248
rect 16577 8239 16635 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 18046 8236 18052 8288
rect 18104 8276 18110 8288
rect 18325 8279 18383 8285
rect 18325 8276 18337 8279
rect 18104 8248 18337 8276
rect 18104 8236 18110 8248
rect 18325 8245 18337 8248
rect 18371 8245 18383 8279
rect 18325 8239 18383 8245
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 19334 8276 19340 8288
rect 18472 8248 19340 8276
rect 18472 8236 18478 8248
rect 19334 8236 19340 8248
rect 19392 8276 19398 8288
rect 19702 8276 19708 8288
rect 19392 8248 19708 8276
rect 19392 8236 19398 8248
rect 19702 8236 19708 8248
rect 19760 8236 19766 8288
rect 19886 8236 19892 8288
rect 19944 8276 19950 8288
rect 20447 8279 20505 8285
rect 20447 8276 20459 8279
rect 19944 8248 20459 8276
rect 19944 8236 19950 8248
rect 20447 8245 20459 8248
rect 20493 8276 20505 8279
rect 21082 8276 21088 8288
rect 20493 8248 21088 8276
rect 20493 8245 20505 8248
rect 20447 8239 20505 8245
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21818 8276 21824 8288
rect 21779 8248 21824 8276
rect 21818 8236 21824 8248
rect 21876 8276 21882 8288
rect 22373 8279 22431 8285
rect 22373 8276 22385 8279
rect 21876 8248 22385 8276
rect 21876 8236 21882 8248
rect 22373 8245 22385 8248
rect 22419 8245 22431 8279
rect 22373 8239 22431 8245
rect 22462 8236 22468 8288
rect 22520 8276 22526 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 22520 8248 22937 8276
rect 22520 8236 22526 8248
rect 22925 8245 22937 8248
rect 22971 8245 22983 8279
rect 22925 8239 22983 8245
rect 1104 8186 23460 8208
rect 1104 8134 8446 8186
rect 8498 8134 8510 8186
rect 8562 8134 8574 8186
rect 8626 8134 8638 8186
rect 8690 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 23460 8186
rect 1104 8112 23460 8134
rect 9306 8072 9312 8084
rect 9219 8044 9312 8072
rect 9306 8032 9312 8044
rect 9364 8072 9370 8084
rect 9582 8072 9588 8084
rect 9364 8044 9588 8072
rect 9364 8032 9370 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12032 8044 12265 8072
rect 12032 8032 12038 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 12621 8075 12679 8081
rect 12621 8041 12633 8075
rect 12667 8072 12679 8075
rect 13170 8072 13176 8084
rect 12667 8044 13176 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 15473 8075 15531 8081
rect 15473 8041 15485 8075
rect 15519 8072 15531 8075
rect 16390 8072 16396 8084
rect 15519 8044 16396 8072
rect 15519 8041 15531 8044
rect 15473 8035 15531 8041
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 16482 8032 16488 8084
rect 16540 8081 16546 8084
rect 16540 8072 16549 8081
rect 16540 8044 17448 8072
rect 16540 8035 16549 8044
rect 16540 8032 16546 8035
rect 8573 8007 8631 8013
rect 8573 7973 8585 8007
rect 8619 8004 8631 8007
rect 9944 8007 10002 8013
rect 8619 7976 9904 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7936 7806 7948
rect 8202 7936 8208 7948
rect 7800 7908 8208 7936
rect 7800 7896 7806 7908
rect 8202 7896 8208 7908
rect 8260 7936 8266 7948
rect 8849 7939 8907 7945
rect 8849 7936 8861 7939
rect 8260 7908 8861 7936
rect 8260 7896 8266 7908
rect 8849 7905 8861 7908
rect 8895 7905 8907 7939
rect 8849 7899 8907 7905
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 9508 7868 9536 7899
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9640 7908 9689 7936
rect 9640 7896 9646 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9766 7896 9772 7948
rect 9824 7896 9830 7948
rect 9876 7936 9904 7976
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 11054 8004 11060 8016
rect 9990 7976 11060 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 13449 8007 13507 8013
rect 13449 8004 13461 8007
rect 11848 7976 13461 8004
rect 11848 7964 11854 7976
rect 13449 7973 13461 7976
rect 13495 7973 13507 8007
rect 13449 7967 13507 7973
rect 14737 8007 14795 8013
rect 14737 7973 14749 8007
rect 14783 8004 14795 8007
rect 14918 8004 14924 8016
rect 14783 7976 14924 8004
rect 14783 7973 14795 7976
rect 14737 7967 14795 7973
rect 14918 7964 14924 7976
rect 14976 7964 14982 8016
rect 17420 8004 17448 8044
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17644 8044 17877 8072
rect 17644 8032 17650 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 18064 8044 18359 8072
rect 18064 8004 18092 8044
rect 17420 7976 18092 8004
rect 18138 7964 18144 8016
rect 18196 8004 18202 8016
rect 18233 8007 18291 8013
rect 18233 8004 18245 8007
rect 18196 7976 18245 8004
rect 18196 7964 18202 7976
rect 18233 7973 18245 7976
rect 18279 7973 18291 8007
rect 18331 8004 18359 8044
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 19150 8072 19156 8084
rect 18564 8044 19156 8072
rect 18564 8032 18570 8044
rect 19150 8032 19156 8044
rect 19208 8072 19214 8084
rect 19334 8072 19340 8084
rect 19208 8044 19340 8072
rect 19208 8032 19214 8044
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 20346 8032 20352 8084
rect 20404 8072 20410 8084
rect 20441 8075 20499 8081
rect 20441 8072 20453 8075
rect 20404 8044 20453 8072
rect 20404 8032 20410 8044
rect 20441 8041 20453 8044
rect 20487 8041 20499 8075
rect 22554 8072 22560 8084
rect 22515 8044 22560 8072
rect 20441 8035 20499 8041
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 22462 8004 22468 8016
rect 18331 7976 18635 8004
rect 18233 7967 18291 7973
rect 18607 7948 18635 7976
rect 20088 7976 22468 8004
rect 9876 7908 10732 7936
rect 9784 7868 9812 7896
rect 9508 7840 9812 7868
rect 10704 7800 10732 7908
rect 10870 7896 10876 7948
rect 10928 7936 10934 7948
rect 11517 7939 11575 7945
rect 11517 7936 11529 7939
rect 10928 7908 11529 7936
rect 10928 7896 10934 7908
rect 11517 7905 11529 7908
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12676 7908 12725 7936
rect 12676 7896 12682 7908
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 13044 7908 13553 7936
rect 13044 7896 13050 7908
rect 13541 7905 13553 7908
rect 13587 7905 13599 7939
rect 13541 7899 13599 7905
rect 14001 7939 14059 7945
rect 14001 7905 14013 7939
rect 14047 7936 14059 7939
rect 14090 7936 14096 7948
rect 14047 7908 14096 7936
rect 14047 7905 14059 7908
rect 14001 7899 14059 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14458 7896 14464 7948
rect 14516 7936 14522 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14516 7908 15301 7936
rect 14516 7896 14522 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 16022 7936 16028 7948
rect 15983 7908 16028 7936
rect 15289 7899 15347 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 16758 7936 16764 7948
rect 16719 7908 16764 7936
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 18046 7936 18052 7948
rect 18003 7908 18052 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18414 7896 18420 7948
rect 18472 7936 18478 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 18472 7908 18521 7936
rect 18472 7896 18478 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 18509 7899 18567 7905
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18832 7939 18890 7945
rect 18832 7936 18844 7939
rect 18656 7908 18844 7936
rect 18656 7896 18662 7908
rect 18832 7905 18844 7908
rect 18878 7905 18890 7939
rect 19978 7936 19984 7948
rect 18832 7899 18890 7905
rect 19168 7908 19984 7936
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11020 7840 11621 7868
rect 11020 7828 11026 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 12066 7868 12072 7880
rect 11839 7840 12072 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 12066 7828 12072 7840
rect 12124 7868 12130 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12124 7840 12817 7868
rect 12124 7828 12130 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13136 7840 13737 7868
rect 13136 7828 13142 7840
rect 13725 7837 13737 7840
rect 13771 7868 13783 7871
rect 14829 7871 14887 7877
rect 13771 7840 14780 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14642 7800 14648 7812
rect 10704 7772 14648 7800
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 11020 7704 11069 7732
rect 11020 7692 11026 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 13081 7735 13139 7741
rect 11204 7704 11249 7732
rect 11204 7692 11210 7704
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13998 7732 14004 7744
rect 13127 7704 14004 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 14550 7732 14556 7744
rect 14231 7704 14556 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 14752 7732 14780 7840
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15378 7868 15384 7880
rect 15059 7840 15384 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 14844 7800 14872 7831
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15654 7868 15660 7880
rect 15615 7840 15660 7868
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 16482 7868 16488 7880
rect 16446 7840 16488 7868
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 18432 7868 18460 7896
rect 17460 7840 18460 7868
rect 19015 7871 19073 7877
rect 17460 7828 17466 7840
rect 19015 7837 19027 7871
rect 19061 7868 19073 7871
rect 19168 7868 19196 7908
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 19061 7840 19196 7868
rect 19245 7871 19303 7877
rect 19061 7837 19073 7840
rect 19015 7831 19073 7837
rect 19245 7837 19257 7871
rect 19291 7868 19303 7871
rect 19334 7868 19340 7880
rect 19291 7840 19340 7868
rect 19291 7837 19303 7840
rect 19245 7831 19303 7837
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 15286 7800 15292 7812
rect 14844 7772 15292 7800
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 20088 7732 20116 7976
rect 22462 7964 22468 7976
rect 22520 7964 22526 8016
rect 22922 8004 22928 8016
rect 22883 7976 22928 8004
rect 22922 7964 22928 7976
rect 22980 7964 22986 8016
rect 21450 7945 21456 7948
rect 21444 7899 21456 7945
rect 21508 7936 21514 7948
rect 22649 7939 22707 7945
rect 21508 7908 21544 7936
rect 21450 7896 21456 7899
rect 21508 7896 21514 7908
rect 22649 7905 22661 7939
rect 22695 7936 22707 7939
rect 23014 7936 23020 7948
rect 22695 7908 23020 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 20898 7868 20904 7880
rect 20859 7840 20904 7868
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 21140 7840 21189 7868
rect 21140 7828 21146 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 20349 7803 20407 7809
rect 20349 7769 20361 7803
rect 20395 7800 20407 7803
rect 20714 7800 20720 7812
rect 20395 7772 20720 7800
rect 20395 7769 20407 7772
rect 20349 7763 20407 7769
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 14752 7704 20116 7732
rect 1104 7642 23460 7664
rect 1104 7590 4714 7642
rect 4766 7590 4778 7642
rect 4830 7590 4842 7642
rect 4894 7590 4906 7642
rect 4958 7590 12178 7642
rect 12230 7590 12242 7642
rect 12294 7590 12306 7642
rect 12358 7590 12370 7642
rect 12422 7590 19642 7642
rect 19694 7590 19706 7642
rect 19758 7590 19770 7642
rect 19822 7590 19834 7642
rect 19886 7590 23460 7642
rect 1104 7568 23460 7590
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 10870 7528 10876 7540
rect 10735 7500 10876 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 14090 7528 14096 7540
rect 12483 7500 13952 7528
rect 14051 7500 14096 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7460 10839 7463
rect 12253 7463 12311 7469
rect 10827 7432 11652 7460
rect 10827 7429 10839 7432
rect 10781 7423 10839 7429
rect 9306 7392 9312 7404
rect 9267 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 11238 7392 11244 7404
rect 11199 7364 11244 7392
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 9576 7327 9634 7333
rect 9576 7293 9588 7327
rect 9622 7324 9634 7327
rect 10962 7324 10968 7336
rect 9622 7296 10968 7324
rect 9622 7293 9634 7296
rect 9576 7287 9634 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11146 7324 11152 7336
rect 11107 7296 11152 7324
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 11440 7268 11468 7355
rect 11624 7333 11652 7432
rect 12253 7429 12265 7463
rect 12299 7460 12311 7463
rect 13924 7460 13952 7500
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 14568 7500 16344 7528
rect 14458 7460 14464 7472
rect 12299 7432 13768 7460
rect 13924 7432 14464 7460
rect 12299 7429 12311 7432
rect 12253 7423 12311 7429
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13740 7392 13768 7432
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 14568 7392 14596 7500
rect 14734 7420 14740 7472
rect 14792 7420 14798 7472
rect 16316 7460 16344 7500
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 16448 7500 17693 7528
rect 16448 7488 16454 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 16316 7432 17540 7460
rect 13740 7364 14596 7392
rect 14752 7392 14780 7420
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14752 7364 14841 7392
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7293 11667 7327
rect 13262 7324 13268 7336
rect 13223 7296 13268 7324
rect 11609 7287 11667 7293
rect 13262 7284 13268 7296
rect 13320 7284 13326 7336
rect 13740 7333 13768 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17402 7392 17408 7404
rect 16724 7364 17408 7392
rect 16724 7352 16730 7364
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14056 7296 14657 7324
rect 14056 7284 14062 7296
rect 14645 7293 14657 7296
rect 14691 7324 14703 7327
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14691 7296 15025 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 15013 7293 15025 7296
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 15160 7296 15393 7324
rect 15160 7284 15166 7296
rect 15381 7293 15393 7296
rect 15427 7324 15439 7327
rect 16574 7324 16580 7336
rect 15427 7296 16580 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16816 7296 17325 7324
rect 16816 7284 16822 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 11422 7216 11428 7268
rect 11480 7256 11486 7268
rect 11698 7256 11704 7268
rect 11480 7228 11704 7256
rect 11480 7216 11486 7228
rect 11698 7216 11704 7228
rect 11756 7256 11762 7268
rect 12618 7256 12624 7268
rect 11756 7228 12624 7256
rect 11756 7216 11762 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 12805 7259 12863 7265
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 13909 7259 13967 7265
rect 12851 7228 13492 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13464 7197 13492 7228
rect 13909 7225 13921 7259
rect 13955 7256 13967 7259
rect 15470 7256 15476 7268
rect 13955 7228 15476 7256
rect 13955 7225 13967 7228
rect 13909 7219 13967 7225
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 15648 7259 15706 7265
rect 15648 7225 15660 7259
rect 15694 7256 15706 7259
rect 16482 7256 16488 7268
rect 15694 7228 16488 7256
rect 15694 7225 15706 7228
rect 15648 7219 15706 7225
rect 16482 7216 16488 7228
rect 16540 7216 16546 7268
rect 17221 7259 17279 7265
rect 17221 7256 17233 7259
rect 16592 7228 17233 7256
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7157 13507 7191
rect 13449 7151 13507 7157
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 14056 7160 14197 7188
rect 14056 7148 14062 7160
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 14185 7151 14243 7157
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 14553 7191 14611 7197
rect 14553 7188 14565 7191
rect 14516 7160 14565 7188
rect 14516 7148 14522 7160
rect 14553 7157 14565 7160
rect 14599 7157 14611 7191
rect 14553 7151 14611 7157
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 14792 7160 15209 7188
rect 14792 7148 14798 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 16592 7188 16620 7228
rect 17221 7225 17233 7228
rect 17267 7225 17279 7259
rect 17512 7256 17540 7432
rect 17696 7392 17724 7491
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 18012 7500 19441 7528
rect 18012 7488 18018 7500
rect 19429 7497 19441 7500
rect 19475 7497 19487 7531
rect 20714 7528 20720 7540
rect 19429 7491 19487 7497
rect 20180 7500 20720 7528
rect 19610 7460 19616 7472
rect 19571 7432 19616 7460
rect 19610 7420 19616 7432
rect 19668 7420 19674 7472
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 17696 7364 18061 7392
rect 18049 7361 18061 7364
rect 18095 7361 18107 7395
rect 19978 7392 19984 7404
rect 18049 7355 18107 7361
rect 19076 7364 19984 7392
rect 17862 7324 17868 7336
rect 17823 7296 17868 7324
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 19076 7324 19104 7364
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7392 20131 7395
rect 20180 7392 20208 7500
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 21450 7488 21456 7540
rect 21508 7528 21514 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21508 7500 21833 7528
rect 21508 7488 21514 7500
rect 21821 7497 21833 7500
rect 21867 7528 21879 7531
rect 21867 7500 22600 7528
rect 21867 7497 21879 7500
rect 21821 7491 21879 7497
rect 20119 7364 20208 7392
rect 20257 7395 20315 7401
rect 20119 7361 20131 7364
rect 20073 7355 20131 7361
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20303 7364 20576 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20548 7336 20576 7364
rect 22278 7352 22284 7404
rect 22336 7392 22342 7404
rect 22572 7401 22600 7500
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 22336 7364 22385 7392
rect 22336 7352 22342 7364
rect 22373 7361 22385 7364
rect 22419 7361 22431 7395
rect 22373 7355 22431 7361
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 17972 7296 19104 7324
rect 17972 7256 18000 7296
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19610 7324 19616 7336
rect 19484 7296 19616 7324
rect 19484 7284 19490 7296
rect 19610 7284 19616 7296
rect 19668 7324 19674 7336
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 19668 7296 20453 7324
rect 19668 7284 19674 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 17512 7228 18000 7256
rect 17221 7219 17279 7225
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 18294 7259 18352 7265
rect 18294 7256 18306 7259
rect 18196 7228 18306 7256
rect 18196 7216 18202 7228
rect 18294 7225 18306 7228
rect 18340 7225 18352 7259
rect 20456 7256 20484 7287
rect 20530 7284 20536 7336
rect 20588 7284 20594 7336
rect 21082 7324 21088 7336
rect 20640 7296 21088 7324
rect 20640 7256 20668 7296
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 22830 7324 22836 7336
rect 22787 7296 22836 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 20714 7265 20720 7268
rect 20456 7228 20668 7256
rect 18294 7219 18352 7225
rect 20708 7219 20720 7265
rect 20772 7256 20778 7268
rect 22094 7256 22100 7268
rect 20772 7228 20808 7256
rect 21928 7228 22100 7256
rect 20714 7216 20720 7219
rect 20772 7216 20778 7228
rect 15344 7160 16620 7188
rect 15344 7148 15350 7160
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 16724 7160 16773 7188
rect 16724 7148 16730 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 17586 7188 17592 7200
rect 16899 7160 17592 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 19334 7188 19340 7200
rect 18104 7160 19340 7188
rect 18104 7148 18110 7160
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19978 7188 19984 7200
rect 19939 7160 19984 7188
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 21928 7197 21956 7228
rect 22094 7216 22100 7228
rect 22152 7256 22158 7268
rect 23474 7256 23480 7268
rect 22152 7228 23480 7256
rect 22152 7216 22158 7228
rect 23474 7216 23480 7228
rect 23532 7216 23538 7268
rect 21913 7191 21971 7197
rect 21913 7157 21925 7191
rect 21959 7157 21971 7191
rect 21913 7151 21971 7157
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22281 7191 22339 7197
rect 22281 7188 22293 7191
rect 22060 7160 22293 7188
rect 22060 7148 22066 7160
rect 22281 7157 22293 7160
rect 22327 7157 22339 7191
rect 22281 7151 22339 7157
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 22925 7191 22983 7197
rect 22925 7188 22937 7191
rect 22612 7160 22937 7188
rect 22612 7148 22618 7160
rect 22925 7157 22937 7160
rect 22971 7157 22983 7191
rect 22925 7151 22983 7157
rect 1104 7098 23460 7120
rect 1104 7046 8446 7098
rect 8498 7046 8510 7098
rect 8562 7046 8574 7098
rect 8626 7046 8638 7098
rect 8690 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 23460 7098
rect 1104 7024 23460 7046
rect 8202 6944 8208 6996
rect 8260 6984 8266 6996
rect 13173 6987 13231 6993
rect 8260 6956 13124 6984
rect 8260 6944 8266 6956
rect 9944 6919 10002 6925
rect 9944 6885 9956 6919
rect 9990 6916 10002 6919
rect 10870 6916 10876 6928
rect 9990 6888 10876 6916
rect 9990 6885 10002 6888
rect 9944 6879 10002 6885
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 12066 6916 12072 6928
rect 11808 6888 12072 6916
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9364 6820 9689 6848
rect 9364 6808 9370 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 11514 6848 11520 6860
rect 11475 6820 11520 6848
rect 9677 6811 9735 6817
rect 11514 6808 11520 6820
rect 11572 6808 11578 6860
rect 11808 6789 11836 6888
rect 12066 6876 12072 6888
rect 12124 6916 12130 6928
rect 12526 6916 12532 6928
rect 12124 6888 12532 6916
rect 12124 6876 12130 6888
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13096 6916 13124 6956
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13262 6984 13268 6996
rect 13219 6956 13268 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13541 6987 13599 6993
rect 13541 6953 13553 6987
rect 13587 6984 13599 6987
rect 14366 6984 14372 6996
rect 13587 6956 14372 6984
rect 13587 6953 13599 6956
rect 13541 6947 13599 6953
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 14734 6984 14740 6996
rect 14695 6956 14740 6984
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 18138 6984 18144 6996
rect 15856 6956 16068 6984
rect 18099 6956 18144 6984
rect 15856 6916 15884 6956
rect 12676 6888 13032 6916
rect 13096 6888 15884 6916
rect 16040 6916 16068 6956
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18598 6984 18604 6996
rect 18559 6956 18604 6984
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 19150 6944 19156 6996
rect 19208 6984 19214 6996
rect 19337 6987 19395 6993
rect 19337 6984 19349 6987
rect 19208 6956 19349 6984
rect 19208 6944 19214 6956
rect 19337 6953 19349 6956
rect 19383 6953 19395 6987
rect 19337 6947 19395 6953
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 22281 6987 22339 6993
rect 22281 6984 22293 6987
rect 20956 6956 22293 6984
rect 20956 6944 20962 6956
rect 22281 6953 22293 6956
rect 22327 6953 22339 6987
rect 22281 6947 22339 6953
rect 19426 6916 19432 6928
rect 16040 6888 19432 6916
rect 12676 6876 12682 6888
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12710 6848 12716 6860
rect 12671 6820 12716 6848
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 13004 6848 13032 6888
rect 19426 6876 19432 6888
rect 19484 6876 19490 6928
rect 21910 6876 21916 6928
rect 21968 6916 21974 6928
rect 23198 6916 23204 6928
rect 21968 6888 23204 6916
rect 21968 6876 21974 6888
rect 23198 6876 23204 6888
rect 23256 6876 23262 6928
rect 13998 6848 14004 6860
rect 13004 6820 13768 6848
rect 13959 6820 14004 6848
rect 11609 6783 11667 6789
rect 11609 6780 11621 6783
rect 11072 6752 11621 6780
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 11072 6653 11100 6752
rect 11609 6749 11621 6752
rect 11655 6749 11667 6783
rect 11609 6743 11667 6749
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6749 11851 6783
rect 12802 6780 12808 6792
rect 12763 6752 12808 6780
rect 11793 6743 11851 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 12986 6780 12992 6792
rect 12947 6752 12992 6780
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13740 6789 13768 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 15556 6851 15614 6857
rect 15556 6848 15568 6851
rect 15028 6820 15568 6848
rect 15028 6789 15056 6820
rect 15556 6817 15568 6820
rect 15602 6848 15614 6851
rect 15838 6848 15844 6860
rect 15602 6820 15844 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16632 6820 16773 6848
rect 16632 6808 16638 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 17028 6851 17086 6857
rect 17028 6817 17040 6851
rect 17074 6848 17086 6851
rect 17402 6848 17408 6860
rect 17074 6820 17408 6848
rect 17074 6817 17086 6820
rect 17028 6811 17086 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 19978 6848 19984 6860
rect 19444 6820 19984 6848
rect 19444 6792 19472 6820
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20622 6848 20628 6860
rect 20211 6820 20628 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 21140 6820 21281 6848
rect 21140 6808 21146 6820
rect 21269 6817 21281 6820
rect 21315 6817 21327 6851
rect 21269 6811 21327 6817
rect 21637 6851 21695 6857
rect 21637 6817 21649 6851
rect 21683 6848 21695 6851
rect 22002 6848 22008 6860
rect 21683 6820 22008 6848
rect 21683 6817 21695 6820
rect 21637 6811 21695 6817
rect 22002 6808 22008 6820
rect 22060 6808 22066 6860
rect 22370 6848 22376 6860
rect 22331 6820 22376 6848
rect 22370 6808 22376 6820
rect 22428 6808 22434 6860
rect 22738 6848 22744 6860
rect 22699 6820 22744 6848
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 13725 6743 13783 6749
rect 14200 6752 14841 6780
rect 12345 6715 12403 6721
rect 12345 6681 12357 6715
rect 12391 6712 12403 6715
rect 13648 6712 13676 6743
rect 14200 6721 14228 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6749 15347 6783
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 15289 6743 15347 6749
rect 12391 6684 13676 6712
rect 14185 6715 14243 6721
rect 12391 6681 12403 6684
rect 12345 6675 12403 6681
rect 14185 6681 14197 6715
rect 14231 6681 14243 6715
rect 15102 6712 15108 6724
rect 14185 6675 14243 6681
rect 14292 6684 15108 6712
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10376 6616 11069 6644
rect 10376 6604 10382 6616
rect 11057 6613 11069 6616
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 11149 6647 11207 6653
rect 11149 6613 11161 6647
rect 11195 6644 11207 6647
rect 11238 6644 11244 6656
rect 11195 6616 11244 6644
rect 11195 6613 11207 6616
rect 11149 6607 11207 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 12894 6644 12900 6656
rect 12207 6616 12900 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14292 6644 14320 6684
rect 15102 6672 15108 6684
rect 15160 6712 15166 6724
rect 15304 6712 15332 6743
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 20254 6780 20260 6792
rect 19576 6752 19621 6780
rect 20215 6752 20260 6780
rect 19576 6740 19582 6752
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 15160 6684 15332 6712
rect 15160 6672 15166 6684
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16540 6684 16681 6712
rect 16540 6672 16546 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 16669 6675 16727 6681
rect 18969 6715 19027 6721
rect 18969 6681 18981 6715
rect 19015 6712 19027 6715
rect 19242 6712 19248 6724
rect 19015 6684 19248 6712
rect 19015 6681 19027 6684
rect 18969 6675 19027 6681
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 20456 6712 20484 6743
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 21818 6780 21824 6792
rect 20588 6752 21824 6780
rect 20588 6740 20594 6752
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 22186 6740 22192 6792
rect 22244 6780 22250 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22244 6752 22477 6780
rect 22244 6740 22250 6752
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 22094 6712 22100 6724
rect 20456 6684 22100 6712
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 13872 6616 14320 6644
rect 14369 6647 14427 6653
rect 13872 6604 13878 6616
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 15562 6644 15568 6656
rect 14415 6616 15568 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19208 6616 19809 6644
rect 19208 6604 19214 6616
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 19797 6607 19855 6613
rect 20438 6604 20444 6656
rect 20496 6644 20502 6656
rect 20717 6647 20775 6653
rect 20717 6644 20729 6647
rect 20496 6616 20729 6644
rect 20496 6604 20502 6616
rect 20717 6613 20729 6616
rect 20763 6613 20775 6647
rect 20717 6607 20775 6613
rect 20990 6604 20996 6656
rect 21048 6644 21054 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 21048 6616 21097 6644
rect 21048 6604 21054 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21453 6647 21511 6653
rect 21453 6644 21465 6647
rect 21324 6616 21465 6644
rect 21324 6604 21330 6616
rect 21453 6613 21465 6616
rect 21499 6613 21511 6647
rect 21910 6644 21916 6656
rect 21871 6616 21916 6644
rect 21453 6607 21511 6613
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 22925 6647 22983 6653
rect 22925 6644 22937 6647
rect 22244 6616 22937 6644
rect 22244 6604 22250 6616
rect 22925 6613 22937 6616
rect 22971 6613 22983 6647
rect 22925 6607 22983 6613
rect 1104 6554 23460 6576
rect 1104 6502 4714 6554
rect 4766 6502 4778 6554
rect 4830 6502 4842 6554
rect 4894 6502 4906 6554
rect 4958 6502 12178 6554
rect 12230 6502 12242 6554
rect 12294 6502 12306 6554
rect 12358 6502 12370 6554
rect 12422 6502 19642 6554
rect 19694 6502 19706 6554
rect 19758 6502 19770 6554
rect 19822 6502 19834 6554
rect 19886 6502 23460 6554
rect 1104 6480 23460 6502
rect 9306 6440 9312 6452
rect 8956 6412 9312 6440
rect 8956 6313 8984 6412
rect 9306 6400 9312 6412
rect 9364 6440 9370 6452
rect 10321 6443 10379 6449
rect 9364 6412 9996 6440
rect 9364 6400 9370 6412
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 9968 6304 9996 6412
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 11054 6440 11060 6452
rect 10367 6412 11060 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 11054 6400 11060 6412
rect 11112 6440 11118 6452
rect 11514 6440 11520 6452
rect 11112 6412 11520 6440
rect 11112 6400 11118 6412
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12986 6440 12992 6452
rect 12584 6412 12992 6440
rect 12584 6400 12590 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15528 6412 15577 6440
rect 15528 6400 15534 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 9968 6276 10425 6304
rect 8941 6267 8999 6273
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 15580 6304 15608 6403
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 17037 6443 17095 6449
rect 17037 6440 17049 6443
rect 15896 6412 17049 6440
rect 15896 6400 15902 6412
rect 17037 6409 17049 6412
rect 17083 6409 17095 6443
rect 23109 6443 23167 6449
rect 23109 6440 23121 6443
rect 17037 6403 17095 6409
rect 18340 6412 23121 6440
rect 17586 6304 17592 6316
rect 15580 6276 15792 6304
rect 17547 6276 17592 6304
rect 10413 6267 10471 6273
rect 9208 6239 9266 6245
rect 9208 6205 9220 6239
rect 9254 6236 9266 6239
rect 10318 6236 10324 6248
rect 9254 6208 10324 6236
rect 9254 6205 9266 6208
rect 9208 6199 9266 6205
rect 10318 6196 10324 6208
rect 10376 6196 10382 6248
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 13814 6236 13820 6248
rect 12759 6208 13820 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 10680 6171 10738 6177
rect 10680 6137 10692 6171
rect 10726 6168 10738 6171
rect 11330 6168 11336 6180
rect 10726 6140 11336 6168
rect 10726 6137 10738 6140
rect 10680 6131 10738 6137
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 12912 6112 12940 6208
rect 13814 6196 13820 6208
rect 13872 6236 13878 6248
rect 14182 6236 14188 6248
rect 13872 6208 14188 6236
rect 13872 6196 13878 6208
rect 14182 6196 14188 6208
rect 14240 6236 14246 6248
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 14240 6208 15669 6236
rect 14240 6196 14246 6208
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 15764 6236 15792 6276
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17773 6307 17831 6313
rect 17773 6273 17785 6307
rect 17819 6304 17831 6307
rect 18138 6304 18144 6316
rect 17819 6276 18144 6304
rect 17819 6273 17831 6276
rect 17773 6267 17831 6273
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 15913 6239 15971 6245
rect 15913 6236 15925 6239
rect 15764 6208 15925 6236
rect 15657 6199 15715 6205
rect 15913 6205 15925 6208
rect 15959 6205 15971 6239
rect 15913 6199 15971 6205
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6236 17555 6239
rect 18230 6236 18236 6248
rect 17543 6208 18236 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 18230 6196 18236 6208
rect 18288 6196 18294 6248
rect 18340 6245 18368 6412
rect 23109 6409 23121 6412
rect 23155 6409 23167 6443
rect 23109 6403 23167 6409
rect 18509 6375 18567 6381
rect 18509 6341 18521 6375
rect 18555 6341 18567 6375
rect 18509 6335 18567 6341
rect 18693 6375 18751 6381
rect 18693 6341 18705 6375
rect 18739 6372 18751 6375
rect 19426 6372 19432 6384
rect 18739 6344 19432 6372
rect 18739 6341 18751 6344
rect 18693 6335 18751 6341
rect 18325 6239 18383 6245
rect 18325 6205 18337 6239
rect 18371 6205 18383 6239
rect 18524 6236 18552 6335
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 20714 6332 20720 6384
rect 20772 6372 20778 6384
rect 20901 6375 20959 6381
rect 20901 6372 20913 6375
rect 20772 6344 20913 6372
rect 20772 6332 20778 6344
rect 20901 6341 20913 6344
rect 20947 6341 20959 6375
rect 20901 6335 20959 6341
rect 19150 6304 19156 6316
rect 19111 6276 19156 6304
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 19392 6276 19437 6304
rect 19392 6264 19398 6276
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 21545 6307 21603 6313
rect 21545 6304 21557 6307
rect 20588 6276 21557 6304
rect 20588 6264 20594 6276
rect 21545 6273 21557 6276
rect 21591 6273 21603 6307
rect 22462 6304 22468 6316
rect 22423 6276 22468 6304
rect 21545 6267 21603 6273
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 19426 6236 19432 6248
rect 18524 6208 19432 6236
rect 18325 6199 18383 6205
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 19525 6196 19531 6248
rect 19583 6236 19589 6248
rect 19794 6245 19800 6248
rect 19788 6236 19800 6245
rect 19583 6208 19628 6236
rect 19707 6208 19800 6236
rect 19583 6196 19589 6208
rect 19788 6199 19800 6208
rect 19852 6236 19858 6248
rect 20346 6236 20352 6248
rect 19852 6208 20352 6236
rect 19794 6196 19800 6199
rect 19852 6196 19858 6208
rect 20346 6196 20352 6208
rect 20404 6196 20410 6248
rect 20898 6196 20904 6248
rect 20956 6236 20962 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 20956 6208 21373 6236
rect 20956 6196 20962 6208
rect 21361 6205 21373 6208
rect 21407 6205 21419 6239
rect 21818 6236 21824 6248
rect 21779 6208 21824 6236
rect 21361 6199 21419 6205
rect 21818 6196 21824 6208
rect 21876 6196 21882 6248
rect 22189 6239 22247 6245
rect 22189 6205 22201 6239
rect 22235 6236 22247 6239
rect 22278 6236 22284 6248
rect 22235 6208 22284 6236
rect 22235 6205 22247 6208
rect 22189 6199 22247 6205
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22388 6208 22753 6236
rect 12980 6171 13038 6177
rect 12980 6137 12992 6171
rect 13026 6168 13038 6171
rect 13998 6168 14004 6180
rect 13026 6140 14004 6168
rect 13026 6137 13038 6140
rect 12980 6131 13038 6137
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 14430 6171 14488 6177
rect 14430 6168 14442 6171
rect 14108 6140 14442 6168
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12894 6060 12900 6112
rect 12952 6060 12958 6112
rect 14108 6109 14136 6140
rect 14430 6137 14442 6140
rect 14476 6168 14488 6171
rect 14734 6168 14740 6180
rect 14476 6140 14740 6168
rect 14476 6137 14488 6140
rect 14430 6131 14488 6137
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 18049 6171 18107 6177
rect 18049 6137 18061 6171
rect 18095 6168 18107 6171
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 18095 6140 19073 6168
rect 18095 6137 18107 6140
rect 18049 6131 18107 6137
rect 19061 6137 19073 6140
rect 19107 6137 19119 6171
rect 19061 6131 19119 6137
rect 20714 6128 20720 6180
rect 20772 6168 20778 6180
rect 21453 6171 21511 6177
rect 21453 6168 21465 6171
rect 20772 6140 21465 6168
rect 20772 6128 20778 6140
rect 21453 6137 21465 6140
rect 21499 6137 21511 6171
rect 21453 6131 21511 6137
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 22388 6168 22416 6208
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 22922 6168 22928 6180
rect 21692 6140 22416 6168
rect 22883 6140 22928 6168
rect 21692 6128 21698 6140
rect 22922 6128 22928 6140
rect 22980 6128 22986 6180
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6069 14151 6103
rect 14093 6063 14151 6069
rect 17129 6103 17187 6109
rect 17129 6069 17141 6103
rect 17175 6100 17187 6103
rect 19334 6100 19340 6112
rect 17175 6072 19340 6100
rect 17175 6069 17187 6072
rect 17129 6063 17187 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 20990 6060 20996 6112
rect 21048 6100 21054 6112
rect 22002 6100 22008 6112
rect 21048 6072 21093 6100
rect 21963 6072 22008 6100
rect 21048 6060 21054 6072
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 1104 6010 23460 6032
rect 1104 5958 8446 6010
rect 8498 5958 8510 6010
rect 8562 5958 8574 6010
rect 8626 5958 8638 6010
rect 8690 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 23460 6010
rect 1104 5936 23460 5958
rect 11330 5896 11336 5908
rect 11291 5868 11336 5896
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14056 5868 14289 5896
rect 14056 5856 14062 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 10220 5831 10278 5837
rect 10220 5797 10232 5831
rect 10266 5828 10278 5831
rect 11054 5828 11060 5840
rect 10266 5800 11060 5828
rect 10266 5797 10278 5800
rect 10220 5791 10278 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11692 5831 11750 5837
rect 11692 5797 11704 5831
rect 11738 5828 11750 5831
rect 11790 5828 11796 5840
rect 11738 5800 11796 5828
rect 11738 5797 11750 5800
rect 11692 5791 11750 5797
rect 11790 5788 11796 5800
rect 11848 5788 11854 5840
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 13142 5831 13200 5837
rect 13142 5828 13154 5831
rect 12768 5800 13154 5828
rect 12768 5788 12774 5800
rect 13142 5797 13154 5800
rect 13188 5828 13200 5831
rect 13722 5828 13728 5840
rect 13188 5800 13728 5828
rect 13188 5797 13200 5800
rect 13142 5791 13200 5797
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 14292 5828 14320 5859
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14734 5896 14740 5908
rect 14424 5868 14469 5896
rect 14695 5868 14740 5896
rect 14424 5856 14430 5868
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 19518 5896 19524 5908
rect 18984 5868 19524 5896
rect 14829 5831 14887 5837
rect 14829 5828 14841 5831
rect 14292 5800 14841 5828
rect 14829 5797 14841 5800
rect 14875 5797 14887 5831
rect 14829 5791 14887 5797
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 15749 5831 15807 5837
rect 15749 5828 15761 5831
rect 15620 5800 15761 5828
rect 15620 5788 15626 5800
rect 15749 5797 15761 5800
rect 15795 5797 15807 5831
rect 15749 5791 15807 5797
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 9953 5763 10011 5769
rect 9953 5760 9965 5763
rect 9364 5732 9965 5760
rect 9364 5720 9370 5732
rect 9953 5729 9965 5732
rect 9999 5760 10011 5763
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 9999 5732 11437 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 11425 5729 11437 5732
rect 11471 5729 11483 5763
rect 12894 5760 12900 5772
rect 12855 5732 12900 5760
rect 11425 5723 11483 5729
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 16482 5760 16488 5772
rect 13044 5732 14964 5760
rect 13044 5720 13050 5732
rect 14936 5701 14964 5732
rect 15948 5732 16488 5760
rect 15948 5701 15976 5732
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16660 5763 16718 5769
rect 16660 5729 16672 5763
rect 16706 5760 16718 5763
rect 17218 5760 17224 5772
rect 16706 5732 17224 5760
rect 16706 5729 16718 5732
rect 16660 5723 16718 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 18230 5760 18236 5772
rect 18191 5732 18236 5760
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 18984 5769 19012 5868
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20346 5896 20352 5908
rect 20307 5868 20352 5896
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 20622 5896 20628 5908
rect 20583 5868 20628 5896
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 20898 5896 20904 5908
rect 20859 5868 20904 5896
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 21266 5896 21272 5908
rect 21227 5868 21272 5896
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 21450 5856 21456 5908
rect 21508 5896 21514 5908
rect 22554 5896 22560 5908
rect 21508 5868 22560 5896
rect 21508 5856 21514 5868
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 23109 5899 23167 5905
rect 23109 5865 23121 5899
rect 23155 5865 23167 5899
rect 23109 5859 23167 5865
rect 19236 5831 19294 5837
rect 19236 5797 19248 5831
rect 19282 5828 19294 5831
rect 22094 5828 22100 5840
rect 19282 5800 22100 5828
rect 19282 5797 19294 5800
rect 19236 5791 19294 5797
rect 22094 5788 22100 5800
rect 22152 5828 22158 5840
rect 23124 5828 23152 5859
rect 22152 5800 23152 5828
rect 22152 5788 22158 5800
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5729 19027 5763
rect 18969 5723 19027 5729
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 20441 5763 20499 5769
rect 20441 5760 20453 5763
rect 19576 5732 20453 5760
rect 19576 5720 19582 5732
rect 20441 5729 20453 5732
rect 20487 5760 20499 5763
rect 20622 5760 20628 5772
rect 20487 5732 20628 5760
rect 20487 5729 20499 5732
rect 20441 5723 20499 5729
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 21996 5763 22054 5769
rect 21996 5729 22008 5763
rect 22042 5760 22054 5763
rect 22922 5760 22928 5772
rect 22042 5732 22928 5760
rect 22042 5729 22054 5732
rect 21996 5723 22054 5729
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 16390 5692 16396 5704
rect 16351 5664 16396 5692
rect 15933 5655 15991 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 17770 5556 17776 5568
rect 17731 5528 17776 5556
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18524 5556 18552 5655
rect 20530 5652 20536 5704
rect 20588 5692 20594 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 20588 5664 21373 5692
rect 20588 5652 20594 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 21450 5652 21456 5704
rect 21508 5692 21514 5704
rect 21729 5695 21787 5701
rect 21508 5664 21553 5692
rect 21508 5652 21514 5664
rect 21729 5661 21741 5695
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 19242 5556 19248 5568
rect 17920 5528 17965 5556
rect 18524 5528 19248 5556
rect 17920 5516 17926 5528
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 21358 5516 21364 5568
rect 21416 5556 21422 5568
rect 21744 5556 21772 5655
rect 21416 5528 21772 5556
rect 21416 5516 21422 5528
rect 1104 5466 23460 5488
rect 1104 5414 4714 5466
rect 4766 5414 4778 5466
rect 4830 5414 4842 5466
rect 4894 5414 4906 5466
rect 4958 5414 12178 5466
rect 12230 5414 12242 5466
rect 12294 5414 12306 5466
rect 12358 5414 12370 5466
rect 12422 5414 19642 5466
rect 19694 5414 19706 5466
rect 19758 5414 19770 5466
rect 19822 5414 19834 5466
rect 19886 5414 23460 5466
rect 1104 5392 23460 5414
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13780 5324 13829 5352
rect 13780 5312 13786 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 13817 5315 13875 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 17276 5324 17325 5352
rect 17276 5312 17282 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18322 5352 18328 5364
rect 18095 5324 18328 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 11388 5188 11437 5216
rect 11388 5176 11394 5188
rect 11425 5185 11437 5188
rect 11471 5185 11483 5219
rect 11425 5179 11483 5185
rect 11609 5219 11667 5225
rect 11609 5185 11621 5219
rect 11655 5216 11667 5219
rect 17328 5216 17356 5315
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 18877 5355 18935 5361
rect 18877 5321 18889 5355
rect 18923 5352 18935 5355
rect 19426 5352 19432 5364
rect 18923 5324 19432 5352
rect 18923 5321 18935 5324
rect 18877 5315 18935 5321
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 20717 5355 20775 5361
rect 19536 5324 20668 5352
rect 18509 5219 18567 5225
rect 18509 5216 18521 5219
rect 11655 5188 12572 5216
rect 17328 5188 18521 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12544 5148 12572 5188
rect 18509 5185 18521 5188
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 19334 5216 19340 5228
rect 18739 5188 19340 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 19536 5225 19564 5324
rect 19705 5287 19763 5293
rect 19705 5253 19717 5287
rect 19751 5284 19763 5287
rect 20346 5284 20352 5296
rect 19751 5256 20352 5284
rect 19751 5253 19763 5256
rect 19705 5247 19763 5253
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 20640 5284 20668 5324
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 21082 5352 21088 5364
rect 20763 5324 21088 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 22186 5352 22192 5364
rect 21560 5324 22192 5352
rect 21450 5284 21456 5296
rect 20640 5256 21456 5284
rect 21450 5244 21456 5256
rect 21508 5244 21514 5296
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5185 19579 5219
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 19521 5179 19579 5185
rect 19904 5188 20269 5216
rect 12986 5148 12992 5160
rect 12544 5120 12992 5148
rect 12437 5111 12495 5117
rect 11333 5083 11391 5089
rect 11333 5049 11345 5083
rect 11379 5080 11391 5083
rect 11790 5080 11796 5092
rect 11379 5052 11796 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11146 5012 11152 5024
rect 11011 4984 11152 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 12452 5012 12480 5111
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 14274 5108 14280 5160
rect 14332 5148 14338 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 14332 5120 14381 5148
rect 14332 5108 14338 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 17589 5151 17647 5157
rect 15979 5120 16436 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 16408 5092 16436 5120
rect 17589 5117 17601 5151
rect 17635 5148 17647 5151
rect 17862 5148 17868 5160
rect 17635 5120 17868 5148
rect 17635 5117 17647 5120
rect 17589 5111 17647 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 19245 5151 19303 5157
rect 19245 5117 19257 5151
rect 19291 5148 19303 5151
rect 19291 5120 19564 5148
rect 19291 5117 19303 5120
rect 19245 5111 19303 5117
rect 19536 5092 19564 5120
rect 12704 5083 12762 5089
rect 12704 5049 12716 5083
rect 12750 5080 12762 5083
rect 12802 5080 12808 5092
rect 12750 5052 12808 5080
rect 12750 5049 12762 5052
rect 12704 5043 12762 5049
rect 12802 5040 12808 5052
rect 12860 5040 12866 5092
rect 16200 5083 16258 5089
rect 16200 5049 16212 5083
rect 16246 5080 16258 5083
rect 16298 5080 16304 5092
rect 16246 5052 16304 5080
rect 16246 5049 16258 5052
rect 16200 5043 16258 5049
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 16390 5040 16396 5092
rect 16448 5040 16454 5092
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 17788 5052 19349 5080
rect 12894 5012 12900 5024
rect 12452 4984 12900 5012
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 17788 5021 17816 5052
rect 19337 5049 19349 5052
rect 19383 5049 19395 5083
rect 19337 5043 19395 5049
rect 19518 5040 19524 5092
rect 19576 5040 19582 5092
rect 17773 5015 17831 5021
rect 17773 4981 17785 5015
rect 17819 4981 17831 5015
rect 17773 4975 17831 4981
rect 17862 4972 17868 5024
rect 17920 5012 17926 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 17920 4984 18429 5012
rect 17920 4972 17926 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 19904 5012 19932 5188
rect 20257 5185 20269 5188
rect 20303 5216 20315 5219
rect 21269 5219 21327 5225
rect 21269 5216 21281 5219
rect 20303 5188 21281 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 21269 5185 21281 5188
rect 21315 5216 21327 5219
rect 21560 5216 21588 5324
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22922 5352 22928 5364
rect 22336 5324 22784 5352
rect 22883 5324 22928 5352
rect 22336 5312 22342 5324
rect 22756 5284 22784 5324
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 23017 5287 23075 5293
rect 23017 5284 23029 5287
rect 22756 5256 23029 5284
rect 23017 5253 23029 5256
rect 23063 5253 23075 5287
rect 23017 5247 23075 5253
rect 21315 5188 21588 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21358 5108 21364 5160
rect 21416 5148 21422 5160
rect 21545 5151 21603 5157
rect 21545 5148 21557 5151
rect 21416 5120 21557 5148
rect 21416 5108 21422 5120
rect 21545 5117 21557 5120
rect 21591 5117 21603 5151
rect 22278 5148 22284 5160
rect 21545 5111 21603 5117
rect 21652 5120 22284 5148
rect 21085 5083 21143 5089
rect 21085 5049 21097 5083
rect 21131 5080 21143 5083
rect 21652 5080 21680 5120
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 21131 5052 21680 5080
rect 21812 5083 21870 5089
rect 21131 5049 21143 5052
rect 21085 5043 21143 5049
rect 21812 5049 21824 5083
rect 21858 5080 21870 5083
rect 22646 5080 22652 5092
rect 21858 5052 22652 5080
rect 21858 5049 21870 5052
rect 21812 5043 21870 5049
rect 22646 5040 22652 5052
rect 22704 5080 22710 5092
rect 22922 5080 22928 5092
rect 22704 5052 22928 5080
rect 22704 5040 22710 5052
rect 22922 5040 22928 5052
rect 22980 5040 22986 5092
rect 20070 5012 20076 5024
rect 19300 4984 19932 5012
rect 20031 4984 20076 5012
rect 19300 4972 19306 4984
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 21177 5015 21235 5021
rect 20220 4984 20265 5012
rect 20220 4972 20226 4984
rect 21177 4981 21189 5015
rect 21223 5012 21235 5015
rect 22370 5012 22376 5024
rect 21223 4984 22376 5012
rect 21223 4981 21235 4984
rect 21177 4975 21235 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 1104 4922 23460 4944
rect 1104 4870 8446 4922
rect 8498 4870 8510 4922
rect 8562 4870 8574 4922
rect 8626 4870 8638 4922
rect 8690 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 23460 4922
rect 1104 4848 23460 4870
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 17865 4811 17923 4817
rect 17865 4777 17877 4811
rect 17911 4808 17923 4811
rect 18230 4808 18236 4820
rect 17911 4780 18236 4808
rect 17911 4777 17923 4780
rect 17865 4771 17923 4777
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 19521 4811 19579 4817
rect 19521 4777 19533 4811
rect 19567 4808 19579 4811
rect 20162 4808 20168 4820
rect 19567 4780 20168 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20533 4811 20591 4817
rect 20533 4808 20545 4811
rect 20312 4780 20545 4808
rect 20312 4768 20318 4780
rect 20533 4777 20545 4780
rect 20579 4777 20591 4811
rect 20533 4771 20591 4777
rect 21453 4811 21511 4817
rect 21453 4777 21465 4811
rect 21499 4808 21511 4811
rect 21634 4808 21640 4820
rect 21499 4780 21640 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 22922 4808 22928 4820
rect 22883 4780 22928 4808
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 11146 4740 11152 4752
rect 11107 4712 11152 4740
rect 11146 4700 11152 4712
rect 11204 4700 11210 4752
rect 16660 4743 16718 4749
rect 16660 4709 16672 4743
rect 16706 4740 16718 4743
rect 17770 4740 17776 4752
rect 16706 4712 17776 4740
rect 16706 4709 16718 4712
rect 16660 4703 16718 4709
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 19334 4740 19340 4752
rect 18984 4712 19340 4740
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4672 16451 4675
rect 16482 4672 16488 4684
rect 16439 4644 16488 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 11422 4604 11428 4616
rect 11383 4576 11428 4604
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 17788 4576 18337 4604
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 11974 4536 11980 4548
rect 10827 4508 11980 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 17788 4480 17816 4576
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4604 18567 4607
rect 18984 4604 19012 4712
rect 19334 4700 19340 4712
rect 19392 4740 19398 4752
rect 20990 4740 20996 4752
rect 19392 4712 20300 4740
rect 19392 4700 19398 4712
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4672 19119 4675
rect 19426 4672 19432 4684
rect 19107 4644 19432 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4672 19947 4675
rect 20162 4672 20168 4684
rect 19935 4644 20168 4672
rect 19935 4641 19947 4644
rect 19889 4635 19947 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 20272 4616 20300 4712
rect 20364 4712 20996 4740
rect 20364 4681 20392 4712
rect 20990 4700 20996 4712
rect 21048 4700 21054 4752
rect 22738 4700 22744 4752
rect 22796 4740 22802 4752
rect 23017 4743 23075 4749
rect 23017 4740 23029 4743
rect 22796 4712 23029 4740
rect 22796 4700 22802 4712
rect 23017 4709 23029 4712
rect 23063 4709 23075 4743
rect 23017 4703 23075 4709
rect 20349 4675 20407 4681
rect 20349 4641 20361 4675
rect 20395 4641 20407 4675
rect 20349 4635 20407 4641
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4641 20959 4675
rect 20901 4635 20959 4641
rect 19150 4604 19156 4616
rect 18555 4576 19012 4604
rect 19111 4576 19156 4604
rect 18555 4573 18567 4576
rect 18509 4567 18567 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19242 4564 19248 4616
rect 19300 4604 19306 4616
rect 19978 4604 19984 4616
rect 19300 4576 19345 4604
rect 19939 4576 19984 4604
rect 19300 4564 19306 4576
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20254 4604 20260 4616
rect 20119 4576 20260 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 20916 4536 20944 4635
rect 21358 4632 21364 4684
rect 21416 4672 21422 4684
rect 21545 4675 21603 4681
rect 21545 4672 21557 4675
rect 21416 4644 21557 4672
rect 21416 4632 21422 4644
rect 21545 4641 21557 4644
rect 21591 4641 21603 4675
rect 21545 4635 21603 4641
rect 21812 4675 21870 4681
rect 21812 4641 21824 4675
rect 21858 4672 21870 4675
rect 22830 4672 22836 4684
rect 21858 4644 22836 4672
rect 21858 4641 21870 4644
rect 21812 4635 21870 4641
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 18739 4508 20944 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 17770 4468 17776 4480
rect 17731 4440 17776 4468
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 19518 4428 19524 4480
rect 19576 4468 19582 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 19576 4440 21097 4468
rect 19576 4428 19582 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 23460 4400
rect 1104 4326 4714 4378
rect 4766 4326 4778 4378
rect 4830 4326 4842 4378
rect 4894 4326 4906 4378
rect 4958 4326 12178 4378
rect 12230 4326 12242 4378
rect 12294 4326 12306 4378
rect 12358 4326 12370 4378
rect 12422 4326 19642 4378
rect 19694 4326 19706 4378
rect 19758 4326 19770 4378
rect 19822 4326 19834 4378
rect 19886 4326 23460 4378
rect 1104 4304 23460 4326
rect 19613 4267 19671 4273
rect 19613 4233 19625 4267
rect 19659 4264 19671 4267
rect 19978 4264 19984 4276
rect 19659 4236 19984 4264
rect 19659 4233 19671 4236
rect 19613 4227 19671 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 22830 4264 22836 4276
rect 22791 4236 22836 4264
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 21358 4128 21364 4140
rect 20956 4100 21364 4128
rect 20956 4088 20962 4100
rect 21358 4088 21364 4100
rect 21416 4128 21422 4140
rect 21453 4131 21511 4137
rect 21453 4128 21465 4131
rect 21416 4100 21465 4128
rect 21416 4088 21422 4100
rect 21453 4097 21465 4100
rect 21499 4097 21511 4131
rect 23014 4128 23020 4140
rect 22975 4100 23020 4128
rect 21453 4091 21511 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 16301 4063 16359 4069
rect 16301 4029 16313 4063
rect 16347 4060 16359 4063
rect 16568 4063 16626 4069
rect 16347 4032 16528 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16500 4004 16528 4032
rect 16568 4029 16580 4063
rect 16614 4060 16626 4063
rect 17770 4060 17776 4072
rect 16614 4032 17776 4060
rect 16614 4029 16626 4032
rect 16568 4023 16626 4029
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 19978 4069 19984 4072
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 18279 4032 19717 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 19705 4029 19717 4032
rect 19751 4060 19763 4063
rect 19751 4032 19932 4060
rect 19751 4029 19763 4032
rect 19705 4023 19763 4029
rect 16482 3952 16488 4004
rect 16540 3952 16546 4004
rect 18500 3995 18558 4001
rect 18500 3961 18512 3995
rect 18546 3992 18558 3995
rect 19518 3992 19524 4004
rect 18546 3964 19524 3992
rect 18546 3961 18558 3964
rect 18500 3955 18558 3961
rect 19518 3952 19524 3964
rect 19576 3992 19582 4004
rect 19794 3992 19800 4004
rect 19576 3964 19800 3992
rect 19576 3952 19582 3964
rect 19794 3952 19800 3964
rect 19852 3952 19858 4004
rect 19904 3992 19932 4032
rect 19972 4023 19984 4069
rect 20036 4060 20042 4072
rect 20036 4032 20072 4060
rect 19978 4020 19984 4023
rect 20036 4020 20042 4032
rect 20898 3992 20904 4004
rect 19904 3964 20904 3992
rect 20898 3952 20904 3964
rect 20956 3952 20962 4004
rect 21720 3995 21778 4001
rect 21720 3961 21732 3995
rect 21766 3992 21778 3995
rect 22738 3992 22744 4004
rect 21766 3964 22744 3992
rect 21766 3961 21778 3964
rect 21720 3955 21778 3961
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 17681 3927 17739 3933
rect 17681 3893 17693 3927
rect 17727 3924 17739 3927
rect 17954 3924 17960 3936
rect 17727 3896 17960 3924
rect 17727 3893 17739 3896
rect 17681 3887 17739 3893
rect 17954 3884 17960 3896
rect 18012 3924 18018 3936
rect 18230 3924 18236 3936
rect 18012 3896 18236 3924
rect 18012 3884 18018 3896
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20220 3896 21097 3924
rect 20220 3884 20226 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 1104 3834 23460 3856
rect 1104 3782 8446 3834
rect 8498 3782 8510 3834
rect 8562 3782 8574 3834
rect 8626 3782 8638 3834
rect 8690 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 23460 3834
rect 1104 3760 23460 3782
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 2332 3692 3525 3720
rect 2332 3596 2360 3692
rect 3513 3689 3525 3692
rect 3559 3720 3571 3723
rect 18046 3720 18052 3732
rect 3559 3692 18052 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 19426 3720 19432 3732
rect 19387 3692 19432 3720
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19794 3720 19800 3732
rect 19755 3692 19800 3720
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20530 3720 20536 3732
rect 20487 3692 20536 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 20530 3680 20536 3692
rect 20588 3680 20594 3732
rect 22186 3680 22192 3732
rect 22244 3720 22250 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22244 3692 22293 3720
rect 22244 3680 22250 3692
rect 22281 3689 22293 3692
rect 22327 3720 22339 3723
rect 22833 3723 22891 3729
rect 22833 3720 22845 3723
rect 22327 3692 22845 3720
rect 22327 3689 22339 3692
rect 22281 3683 22339 3689
rect 22833 3689 22845 3692
rect 22879 3689 22891 3723
rect 22833 3683 22891 3689
rect 3142 3652 3148 3664
rect 3103 3624 3148 3652
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 16752 3655 16810 3661
rect 16752 3621 16764 3655
rect 16798 3652 16810 3655
rect 17954 3652 17960 3664
rect 16798 3624 17960 3652
rect 16798 3621 16810 3624
rect 16752 3615 16810 3621
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 20272 3652 20300 3680
rect 22002 3652 22008 3664
rect 20088 3624 22008 3652
rect 2314 3584 2320 3596
rect 2227 3556 2320 3584
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18213 3587 18271 3593
rect 18213 3584 18225 3587
rect 17920 3556 18225 3584
rect 17920 3544 17926 3556
rect 18213 3553 18225 3556
rect 18259 3553 18271 3587
rect 18213 3547 18271 3553
rect 16482 3516 16488 3528
rect 16443 3488 16488 3516
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17954 3516 17960 3528
rect 17915 3488 17960 3516
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 20088 3525 20116 3624
rect 22002 3612 22008 3624
rect 22060 3652 22066 3664
rect 22060 3624 22968 3652
rect 22060 3612 22066 3624
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20346 3584 20352 3596
rect 20303 3556 20352 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 21157 3587 21215 3593
rect 21157 3584 21169 3587
rect 21048 3556 21169 3584
rect 21048 3544 21054 3556
rect 21157 3553 21169 3556
rect 21203 3553 21215 3587
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 21157 3547 21215 3553
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 22940 3528 22968 3624
rect 19889 3519 19947 3525
rect 19889 3516 19901 3519
rect 19352 3488 19901 3516
rect 19352 3460 19380 3488
rect 19889 3485 19901 3488
rect 19935 3485 19947 3519
rect 19889 3479 19947 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3485 20131 3519
rect 22922 3516 22928 3528
rect 22835 3488 22928 3516
rect 20073 3479 20131 3485
rect 22922 3476 22928 3488
rect 22980 3476 22986 3528
rect 19334 3448 19340 3460
rect 19247 3420 19340 3448
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 22370 3408 22376 3460
rect 22428 3448 22434 3460
rect 22428 3420 22473 3448
rect 22428 3408 22434 3420
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 17865 3383 17923 3389
rect 17865 3380 17877 3383
rect 17828 3352 17877 3380
rect 17828 3340 17834 3352
rect 17865 3349 17877 3352
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22186 3380 22192 3392
rect 22060 3352 22192 3380
rect 22060 3340 22066 3352
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 1104 3290 23460 3312
rect 1104 3238 4714 3290
rect 4766 3238 4778 3290
rect 4830 3238 4842 3290
rect 4894 3238 4906 3290
rect 4958 3238 12178 3290
rect 12230 3238 12242 3290
rect 12294 3238 12306 3290
rect 12358 3238 12370 3290
rect 12422 3238 19642 3290
rect 19694 3238 19706 3290
rect 19758 3238 19770 3290
rect 19822 3238 19834 3290
rect 19886 3238 23460 3290
rect 1104 3216 23460 3238
rect 2314 3176 2320 3188
rect 1780 3148 2320 3176
rect 1780 2981 1808 3148
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 2498 3136 2504 3188
rect 2556 3176 2562 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2556 3148 2973 3176
rect 2556 3136 2562 3148
rect 2961 3145 2973 3148
rect 3007 3176 3019 3179
rect 10226 3176 10232 3188
rect 3007 3148 10232 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 10226 3136 10232 3148
rect 10284 3176 10290 3188
rect 17862 3176 17868 3188
rect 10284 3148 17448 3176
rect 17823 3148 17868 3176
rect 10284 3136 10290 3148
rect 2038 3068 2044 3120
rect 2096 3108 2102 3120
rect 2685 3111 2743 3117
rect 2685 3108 2697 3111
rect 2096 3080 2697 3108
rect 2096 3068 2102 3080
rect 2685 3077 2697 3080
rect 2731 3077 2743 3111
rect 17420 3108 17448 3148
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 19150 3176 19156 3188
rect 18095 3148 19156 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 20990 3136 20996 3188
rect 21048 3176 21054 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 21048 3148 22201 3176
rect 21048 3136 21054 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 22189 3139 22247 3145
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 22336 3148 22381 3176
rect 22336 3136 22342 3148
rect 18874 3108 18880 3120
rect 17420 3080 18880 3108
rect 2685 3071 2743 3077
rect 18874 3068 18880 3080
rect 18932 3068 18938 3120
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 22922 3040 22928 3052
rect 18739 3012 19472 3040
rect 22883 3012 22928 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 2498 2981 2504 2984
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2941 1823 2975
rect 1765 2935 1823 2941
rect 2489 2975 2504 2981
rect 2489 2941 2501 2975
rect 2489 2935 2504 2941
rect 2498 2932 2504 2935
rect 2556 2932 2562 2984
rect 6086 2972 6092 2984
rect 6047 2944 6092 2972
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 16482 2972 16488 2984
rect 16395 2944 16488 2972
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 17862 2932 17868 2984
rect 17920 2972 17926 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17920 2944 18429 2972
rect 17920 2932 17926 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 16500 2836 16528 2932
rect 16752 2907 16810 2913
rect 16752 2873 16764 2907
rect 16798 2904 16810 2907
rect 17770 2904 17776 2916
rect 16798 2876 17776 2904
rect 16798 2873 16810 2876
rect 16752 2867 16810 2873
rect 17770 2864 17776 2876
rect 17828 2904 17834 2916
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 17828 2876 18521 2904
rect 17828 2864 17834 2876
rect 18509 2873 18521 2876
rect 18555 2873 18567 2907
rect 18509 2867 18567 2873
rect 18046 2836 18052 2848
rect 16500 2808 18052 2836
rect 18046 2796 18052 2808
rect 18104 2836 18110 2848
rect 19352 2836 19380 2935
rect 19444 2904 19472 3012
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 19604 2975 19662 2981
rect 19604 2941 19616 2975
rect 19650 2972 19662 2975
rect 20162 2972 20168 2984
rect 19650 2944 20168 2972
rect 19650 2941 19662 2944
rect 19604 2935 19662 2941
rect 20162 2932 20168 2944
rect 20220 2932 20226 2984
rect 20809 2975 20867 2981
rect 20809 2972 20821 2975
rect 20364 2944 20821 2972
rect 20254 2904 20260 2916
rect 19444 2876 20260 2904
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 20364 2836 20392 2944
rect 20809 2941 20821 2944
rect 20855 2972 20867 2975
rect 20898 2972 20904 2984
rect 20855 2944 20904 2972
rect 20855 2941 20867 2944
rect 20809 2935 20867 2941
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 22646 2972 22652 2984
rect 22607 2944 22652 2972
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 22741 2975 22799 2981
rect 22741 2941 22753 2975
rect 22787 2972 22799 2975
rect 22830 2972 22836 2984
rect 22787 2944 22836 2972
rect 22787 2941 22799 2944
rect 22741 2935 22799 2941
rect 22830 2932 22836 2944
rect 22888 2932 22894 2984
rect 21054 2907 21112 2913
rect 21054 2904 21066 2907
rect 20732 2876 21066 2904
rect 20732 2848 20760 2876
rect 21054 2873 21066 2876
rect 21100 2873 21112 2907
rect 21054 2867 21112 2873
rect 20714 2836 20720 2848
rect 18104 2808 20392 2836
rect 20627 2808 20720 2836
rect 18104 2796 18110 2808
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 22646 2796 22652 2848
rect 22704 2836 22710 2848
rect 23014 2836 23020 2848
rect 22704 2808 23020 2836
rect 22704 2796 22710 2808
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 1104 2746 23460 2768
rect 1104 2694 8446 2746
rect 8498 2694 8510 2746
rect 8562 2694 8574 2746
rect 8626 2694 8638 2746
rect 8690 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 23460 2746
rect 1104 2672 23460 2694
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19576 2604 19717 2632
rect 19576 2592 19582 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 20070 2592 20076 2644
rect 20128 2632 20134 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 20128 2604 20269 2632
rect 20128 2592 20134 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20257 2595 20315 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22557 2635 22615 2641
rect 22557 2601 22569 2635
rect 22603 2632 22615 2635
rect 22738 2632 22744 2644
rect 22603 2604 22744 2632
rect 22603 2601 22615 2604
rect 22557 2595 22615 2601
rect 22738 2592 22744 2604
rect 22796 2592 22802 2644
rect 18592 2567 18650 2573
rect 18592 2533 18604 2567
rect 18638 2564 18650 2567
rect 19334 2564 19340 2576
rect 18638 2536 19340 2564
rect 18638 2533 18650 2536
rect 18592 2527 18650 2533
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 20990 2564 20996 2576
rect 20671 2536 20996 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 20990 2524 20996 2536
rect 21048 2524 21054 2576
rect 21444 2567 21502 2573
rect 21444 2533 21456 2567
rect 21490 2564 21502 2567
rect 22002 2564 22008 2576
rect 21490 2536 22008 2564
rect 21490 2533 21502 2536
rect 21444 2527 21502 2533
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18104 2468 18337 2496
rect 18104 2456 18110 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20956 2468 21189 2496
rect 20956 2456 20962 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 22646 2496 22652 2508
rect 22607 2468 22652 2496
rect 21177 2459 21235 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20809 2431 20867 2437
rect 20809 2428 20821 2431
rect 20312 2400 20821 2428
rect 20312 2388 20318 2400
rect 20809 2397 20821 2400
rect 20855 2397 20867 2431
rect 20809 2391 20867 2397
rect 22462 2388 22468 2440
rect 22520 2428 22526 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22520 2400 22845 2428
rect 22520 2388 22526 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 1104 2202 23460 2224
rect 1104 2150 4714 2202
rect 4766 2150 4778 2202
rect 4830 2150 4842 2202
rect 4894 2150 4906 2202
rect 4958 2150 12178 2202
rect 12230 2150 12242 2202
rect 12294 2150 12306 2202
rect 12358 2150 12370 2202
rect 12422 2150 19642 2202
rect 19694 2150 19706 2202
rect 19758 2150 19770 2202
rect 19822 2150 19834 2202
rect 19886 2150 23460 2202
rect 1104 2128 23460 2150
<< via1 >>
rect 5540 22448 5592 22500
rect 6920 22448 6972 22500
rect 8668 22448 8720 22500
rect 5448 22380 5500 22432
rect 6644 22380 6696 22432
rect 13820 22380 13872 22432
rect 14832 22380 14884 22432
rect 8446 22278 8498 22330
rect 8510 22278 8562 22330
rect 8574 22278 8626 22330
rect 8638 22278 8690 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 5356 22108 5408 22160
rect 6920 22151 6972 22160
rect 6920 22117 6929 22151
rect 6929 22117 6963 22151
rect 6963 22117 6972 22151
rect 6920 22108 6972 22117
rect 5264 22040 5316 22092
rect 5540 22083 5592 22092
rect 5540 22049 5549 22083
rect 5549 22049 5583 22083
rect 5583 22049 5592 22083
rect 6276 22083 6328 22092
rect 5540 22040 5592 22049
rect 6276 22049 6285 22083
rect 6285 22049 6319 22083
rect 6319 22049 6328 22083
rect 6276 22040 6328 22049
rect 7564 22176 7616 22228
rect 8024 22176 8076 22228
rect 8392 22108 8444 22160
rect 10600 22151 10652 22160
rect 2412 21972 2464 22024
rect 5908 21972 5960 22024
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 7840 22015 7892 22024
rect 6460 21972 6512 21981
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 10140 22083 10192 22092
rect 10140 22049 10149 22083
rect 10149 22049 10183 22083
rect 10183 22049 10192 22083
rect 10140 22040 10192 22049
rect 10600 22117 10609 22151
rect 10609 22117 10643 22151
rect 10643 22117 10652 22151
rect 10600 22108 10652 22117
rect 13084 22108 13136 22160
rect 14188 22108 14240 22160
rect 12624 22040 12676 22092
rect 13176 22040 13228 22092
rect 13728 22040 13780 22092
rect 14832 22083 14884 22092
rect 14832 22049 14841 22083
rect 14841 22049 14875 22083
rect 14875 22049 14884 22083
rect 14832 22040 14884 22049
rect 15292 22040 15344 22092
rect 18052 22108 18104 22160
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 11060 21972 11112 22024
rect 11980 21972 12032 22024
rect 13360 21972 13412 22024
rect 4160 21904 4212 21956
rect 5264 21904 5316 21956
rect 5816 21904 5868 21956
rect 12900 21947 12952 21956
rect 12900 21913 12909 21947
rect 12909 21913 12943 21947
rect 12943 21913 12952 21947
rect 12900 21904 12952 21913
rect 14464 21972 14516 22024
rect 14924 21972 14976 22024
rect 15200 21904 15252 21956
rect 19432 22040 19484 22092
rect 23572 22083 23624 22092
rect 23572 22049 23581 22083
rect 23581 22049 23615 22083
rect 23615 22049 23624 22083
rect 23572 22040 23624 22049
rect 17868 21904 17920 21956
rect 2320 21879 2372 21888
rect 2320 21845 2329 21879
rect 2329 21845 2363 21879
rect 2363 21845 2372 21879
rect 2320 21836 2372 21845
rect 4528 21879 4580 21888
rect 4528 21845 4537 21879
rect 4537 21845 4571 21879
rect 4571 21845 4580 21879
rect 4528 21836 4580 21845
rect 5540 21836 5592 21888
rect 5724 21879 5776 21888
rect 5724 21845 5733 21879
rect 5733 21845 5767 21879
rect 5767 21845 5776 21879
rect 5724 21836 5776 21845
rect 7196 21836 7248 21888
rect 7656 21836 7708 21888
rect 7840 21836 7892 21888
rect 13820 21836 13872 21888
rect 14004 21879 14056 21888
rect 14004 21845 14013 21879
rect 14013 21845 14047 21879
rect 14047 21845 14056 21879
rect 14004 21836 14056 21845
rect 14740 21836 14792 21888
rect 14924 21836 14976 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 16304 21836 16356 21888
rect 17408 21879 17460 21888
rect 17408 21845 17417 21879
rect 17417 21845 17451 21879
rect 17451 21845 17460 21879
rect 24124 21904 24176 21956
rect 17408 21836 17460 21845
rect 18236 21836 18288 21888
rect 4714 21734 4766 21786
rect 4778 21734 4830 21786
rect 4842 21734 4894 21786
rect 4906 21734 4958 21786
rect 12178 21734 12230 21786
rect 12242 21734 12294 21786
rect 12306 21734 12358 21786
rect 12370 21734 12422 21786
rect 19642 21734 19694 21786
rect 19706 21734 19758 21786
rect 19770 21734 19822 21786
rect 19834 21734 19886 21786
rect 296 21632 348 21684
rect 2872 21632 2924 21684
rect 5172 21632 5224 21684
rect 6736 21632 6788 21684
rect 7564 21675 7616 21684
rect 7564 21641 7573 21675
rect 7573 21641 7607 21675
rect 7607 21641 7616 21675
rect 7564 21632 7616 21641
rect 7656 21632 7708 21684
rect 11796 21632 11848 21684
rect 940 21564 992 21616
rect 2320 21496 2372 21548
rect 2412 21428 2464 21480
rect 2596 21471 2648 21480
rect 2596 21437 2605 21471
rect 2605 21437 2639 21471
rect 2639 21437 2648 21471
rect 2596 21428 2648 21437
rect 4620 21428 4672 21480
rect 5080 21428 5132 21480
rect 5908 21496 5960 21548
rect 7840 21496 7892 21548
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 4344 21360 4396 21412
rect 4528 21360 4580 21412
rect 5448 21360 5500 21412
rect 6736 21428 6788 21480
rect 8024 21428 8076 21480
rect 9036 21471 9088 21480
rect 9036 21437 9045 21471
rect 9045 21437 9079 21471
rect 9079 21437 9088 21471
rect 9036 21428 9088 21437
rect 10048 21428 10100 21480
rect 10508 21471 10560 21480
rect 10508 21437 10517 21471
rect 10517 21437 10551 21471
rect 10551 21437 10560 21471
rect 10508 21428 10560 21437
rect 12624 21632 12676 21684
rect 13728 21632 13780 21684
rect 13912 21632 13964 21684
rect 12072 21564 12124 21616
rect 14924 21632 14976 21684
rect 17684 21675 17736 21684
rect 13912 21471 13964 21480
rect 4160 21292 4212 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 6920 21292 6972 21344
rect 7288 21292 7340 21344
rect 7748 21292 7800 21344
rect 8208 21292 8260 21344
rect 8300 21292 8352 21344
rect 10048 21292 10100 21344
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 10692 21360 10744 21412
rect 13912 21437 13921 21471
rect 13921 21437 13955 21471
rect 13955 21437 13964 21471
rect 13912 21428 13964 21437
rect 14004 21428 14056 21480
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 21916 21632 21968 21684
rect 20260 21564 20312 21616
rect 21824 21564 21876 21616
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 18604 21496 18656 21548
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 18236 21428 18288 21480
rect 18328 21428 18380 21480
rect 12532 21360 12584 21412
rect 13084 21360 13136 21412
rect 14188 21403 14240 21412
rect 14188 21369 14222 21403
rect 14222 21369 14240 21403
rect 14188 21360 14240 21369
rect 19248 21360 19300 21412
rect 11060 21292 11112 21344
rect 11152 21292 11204 21344
rect 14464 21292 14516 21344
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 15752 21292 15804 21344
rect 16580 21292 16632 21344
rect 16856 21292 16908 21344
rect 17040 21335 17092 21344
rect 17040 21301 17049 21335
rect 17049 21301 17083 21335
rect 17083 21301 17092 21335
rect 17040 21292 17092 21301
rect 17132 21335 17184 21344
rect 17132 21301 17141 21335
rect 17141 21301 17175 21335
rect 17175 21301 17184 21335
rect 17132 21292 17184 21301
rect 23296 21428 23348 21480
rect 22560 21292 22612 21344
rect 8446 21190 8498 21242
rect 8510 21190 8562 21242
rect 8574 21190 8626 21242
rect 8638 21190 8690 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 1584 21088 1636 21140
rect 2228 21088 2280 21140
rect 2596 21020 2648 21072
rect 2964 20952 3016 21004
rect 5080 21088 5132 21140
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 4160 21020 4212 21072
rect 4528 21020 4580 21072
rect 5816 21088 5868 21140
rect 6000 21088 6052 21140
rect 6644 21088 6696 21140
rect 3976 20884 4028 20936
rect 5172 20952 5224 21004
rect 6460 21063 6512 21072
rect 6460 21029 6494 21063
rect 6494 21029 6512 21063
rect 6460 21020 6512 21029
rect 10140 21088 10192 21140
rect 11060 21131 11112 21140
rect 11060 21097 11069 21131
rect 11069 21097 11103 21131
rect 11103 21097 11112 21131
rect 11060 21088 11112 21097
rect 8116 21020 8168 21072
rect 9036 21020 9088 21072
rect 9220 21020 9272 21072
rect 5816 20884 5868 20936
rect 6184 20927 6236 20936
rect 6184 20893 6200 20927
rect 6200 20893 6234 20927
rect 6234 20893 6236 20927
rect 6184 20884 6236 20893
rect 7196 20884 7248 20936
rect 3792 20748 3844 20800
rect 4344 20748 4396 20800
rect 5172 20748 5224 20800
rect 6184 20748 6236 20800
rect 8392 20748 8444 20800
rect 9772 20952 9824 21004
rect 10508 20952 10560 21004
rect 11888 21088 11940 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 14188 21088 14240 21140
rect 13176 21020 13228 21072
rect 13728 21020 13780 21072
rect 11796 20952 11848 21004
rect 15108 21020 15160 21072
rect 15568 20995 15620 21004
rect 15568 20961 15602 20995
rect 15602 20961 15620 20995
rect 15568 20952 15620 20961
rect 17316 21088 17368 21140
rect 17224 21020 17276 21072
rect 22008 21088 22060 21140
rect 21548 20952 21600 21004
rect 11612 20816 11664 20868
rect 11336 20791 11388 20800
rect 11336 20757 11345 20791
rect 11345 20757 11379 20791
rect 11379 20757 11388 20791
rect 11336 20748 11388 20757
rect 12624 20748 12676 20800
rect 15200 20884 15252 20936
rect 13912 20748 13964 20800
rect 14372 20748 14424 20800
rect 17408 20748 17460 20800
rect 18052 20884 18104 20936
rect 19524 20748 19576 20800
rect 23664 20952 23716 21004
rect 23204 20748 23256 20800
rect 4714 20646 4766 20698
rect 4778 20646 4830 20698
rect 4842 20646 4894 20698
rect 4906 20646 4958 20698
rect 12178 20646 12230 20698
rect 12242 20646 12294 20698
rect 12306 20646 12358 20698
rect 12370 20646 12422 20698
rect 19642 20646 19694 20698
rect 19706 20646 19758 20698
rect 19770 20646 19822 20698
rect 19834 20646 19886 20698
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 3516 20544 3568 20596
rect 1584 20451 1636 20460
rect 1584 20417 1593 20451
rect 1593 20417 1627 20451
rect 1627 20417 1636 20451
rect 1584 20408 1636 20417
rect 3148 20408 3200 20460
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 4344 20451 4396 20460
rect 4344 20417 4353 20451
rect 4353 20417 4387 20451
rect 4387 20417 4396 20451
rect 4344 20408 4396 20417
rect 6460 20544 6512 20596
rect 6644 20544 6696 20596
rect 10692 20587 10744 20596
rect 6920 20476 6972 20528
rect 10692 20553 10701 20587
rect 10701 20553 10735 20587
rect 10735 20553 10744 20587
rect 10692 20544 10744 20553
rect 10784 20544 10836 20596
rect 13084 20544 13136 20596
rect 13176 20544 13228 20596
rect 13728 20544 13780 20596
rect 11888 20476 11940 20528
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 6276 20408 6328 20460
rect 9220 20408 9272 20460
rect 10876 20408 10928 20460
rect 15384 20544 15436 20596
rect 15568 20544 15620 20596
rect 17132 20544 17184 20596
rect 19432 20544 19484 20596
rect 22468 20587 22520 20596
rect 22468 20553 22477 20587
rect 22477 20553 22511 20587
rect 22511 20553 22520 20587
rect 22468 20544 22520 20553
rect 16856 20476 16908 20528
rect 17684 20476 17736 20528
rect 2964 20340 3016 20392
rect 4160 20340 4212 20392
rect 4988 20340 5040 20392
rect 5908 20340 5960 20392
rect 6184 20340 6236 20392
rect 6736 20340 6788 20392
rect 7196 20340 7248 20392
rect 7932 20340 7984 20392
rect 8392 20340 8444 20392
rect 5632 20272 5684 20324
rect 10416 20340 10468 20392
rect 10600 20340 10652 20392
rect 2964 20204 3016 20256
rect 3056 20247 3108 20256
rect 3056 20213 3065 20247
rect 3065 20213 3099 20247
rect 3099 20213 3108 20247
rect 3884 20247 3936 20256
rect 3056 20204 3108 20213
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 7012 20204 7064 20256
rect 9312 20272 9364 20324
rect 9680 20272 9732 20324
rect 8852 20204 8904 20256
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 13544 20340 13596 20392
rect 15660 20408 15712 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 14188 20340 14240 20392
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 16580 20340 16632 20392
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 10048 20204 10100 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 14556 20272 14608 20324
rect 19064 20476 19116 20528
rect 23480 20476 23532 20528
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 19524 20340 19576 20392
rect 22376 20408 22428 20460
rect 22928 20408 22980 20460
rect 16488 20204 16540 20256
rect 22192 20272 22244 20324
rect 22744 20272 22796 20324
rect 17868 20204 17920 20256
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 22100 20247 22152 20256
rect 22100 20213 22109 20247
rect 22109 20213 22143 20247
rect 22143 20213 22152 20247
rect 22652 20247 22704 20256
rect 22100 20204 22152 20213
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23572 20204 23624 20256
rect 8446 20102 8498 20154
rect 8510 20102 8562 20154
rect 8574 20102 8626 20154
rect 8638 20102 8690 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 3884 20000 3936 20052
rect 2872 19932 2924 19984
rect 3056 19932 3108 19984
rect 6092 19975 6144 19984
rect 6092 19941 6101 19975
rect 6101 19941 6135 19975
rect 6135 19941 6144 19975
rect 6092 19932 6144 19941
rect 7012 19975 7064 19984
rect 7012 19941 7046 19975
rect 7046 19941 7064 19975
rect 7012 19932 7064 19941
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 2780 19864 2832 19916
rect 3608 19864 3660 19916
rect 5264 19907 5316 19916
rect 3516 19839 3568 19848
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 3976 19796 4028 19848
rect 5264 19873 5273 19907
rect 5273 19873 5307 19907
rect 5307 19873 5316 19907
rect 5264 19864 5316 19873
rect 5540 19864 5592 19916
rect 8852 20000 8904 20052
rect 10232 20000 10284 20052
rect 13544 20000 13596 20052
rect 13820 20043 13872 20052
rect 13820 20009 13829 20043
rect 13829 20009 13863 20043
rect 13863 20009 13872 20043
rect 13820 20000 13872 20009
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 14556 20043 14608 20052
rect 14556 20009 14565 20043
rect 14565 20009 14599 20043
rect 14599 20009 14608 20043
rect 14556 20000 14608 20009
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 15200 20000 15252 20052
rect 16212 20000 16264 20052
rect 12532 19932 12584 19984
rect 22284 20000 22336 20052
rect 22468 20043 22520 20052
rect 22468 20009 22477 20043
rect 22477 20009 22511 20043
rect 22511 20009 22520 20043
rect 22468 20000 22520 20009
rect 22836 20043 22888 20052
rect 22836 20009 22845 20043
rect 22845 20009 22879 20043
rect 22879 20009 22888 20043
rect 22836 20000 22888 20009
rect 16580 19975 16632 19984
rect 16580 19941 16589 19975
rect 16589 19941 16623 19975
rect 16623 19941 16632 19975
rect 16580 19932 16632 19941
rect 17040 19932 17092 19984
rect 17868 19975 17920 19984
rect 17868 19941 17902 19975
rect 17902 19941 17920 19975
rect 17868 19932 17920 19941
rect 18052 19932 18104 19984
rect 20904 19932 20956 19984
rect 22376 19932 22428 19984
rect 3792 19728 3844 19780
rect 5632 19796 5684 19848
rect 6184 19839 6236 19848
rect 6184 19805 6193 19839
rect 6193 19805 6227 19839
rect 6227 19805 6236 19839
rect 6184 19796 6236 19805
rect 3056 19703 3108 19712
rect 3056 19669 3065 19703
rect 3065 19669 3099 19703
rect 3099 19669 3108 19703
rect 4068 19703 4120 19712
rect 3056 19660 3108 19669
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 5540 19728 5592 19780
rect 5724 19728 5776 19780
rect 5816 19728 5868 19780
rect 6736 19839 6788 19848
rect 6736 19805 6745 19839
rect 6745 19805 6779 19839
rect 6779 19805 6788 19839
rect 8852 19864 8904 19916
rect 9312 19864 9364 19916
rect 9220 19839 9272 19848
rect 6736 19796 6788 19805
rect 7840 19728 7892 19780
rect 6736 19660 6788 19712
rect 7104 19660 7156 19712
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 9680 19796 9732 19848
rect 9956 19796 10008 19848
rect 9128 19728 9180 19780
rect 9772 19728 9824 19780
rect 12716 19864 12768 19916
rect 11152 19839 11204 19848
rect 11152 19805 11161 19839
rect 11161 19805 11195 19839
rect 11195 19805 11204 19839
rect 11152 19796 11204 19805
rect 11244 19796 11296 19848
rect 12808 19796 12860 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13360 19864 13412 19916
rect 13728 19907 13780 19916
rect 13728 19873 13737 19907
rect 13737 19873 13771 19907
rect 13771 19873 13780 19907
rect 13728 19864 13780 19873
rect 15476 19864 15528 19916
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 16488 19907 16540 19916
rect 16488 19873 16497 19907
rect 16497 19873 16531 19907
rect 16531 19873 16540 19907
rect 16488 19864 16540 19873
rect 13912 19839 13964 19848
rect 13912 19805 13921 19839
rect 13921 19805 13955 19839
rect 13955 19805 13964 19839
rect 13912 19796 13964 19805
rect 14556 19728 14608 19780
rect 9864 19660 9916 19712
rect 11244 19660 11296 19712
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 15844 19839 15896 19848
rect 14740 19796 14792 19805
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 16580 19796 16632 19848
rect 16304 19728 16356 19780
rect 19064 19864 19116 19916
rect 20076 19864 20128 19916
rect 21364 19907 21416 19916
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 22284 19907 22336 19916
rect 17408 19796 17460 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 19432 19796 19484 19848
rect 15844 19660 15896 19712
rect 21916 19728 21968 19780
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 22652 19907 22704 19916
rect 22652 19873 22661 19907
rect 22661 19873 22695 19907
rect 22695 19873 22704 19907
rect 22652 19864 22704 19873
rect 23388 19864 23440 19916
rect 17132 19703 17184 19712
rect 17132 19669 17141 19703
rect 17141 19669 17175 19703
rect 17175 19669 17184 19703
rect 17132 19660 17184 19669
rect 17960 19660 18012 19712
rect 20444 19660 20496 19712
rect 20996 19703 21048 19712
rect 20996 19669 21005 19703
rect 21005 19669 21039 19703
rect 21039 19669 21048 19703
rect 20996 19660 21048 19669
rect 22284 19660 22336 19712
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 4714 19558 4766 19610
rect 4778 19558 4830 19610
rect 4842 19558 4894 19610
rect 4906 19558 4958 19610
rect 12178 19558 12230 19610
rect 12242 19558 12294 19610
rect 12306 19558 12358 19610
rect 12370 19558 12422 19610
rect 19642 19558 19694 19610
rect 19706 19558 19758 19610
rect 19770 19558 19822 19610
rect 19834 19558 19886 19610
rect 5264 19456 5316 19508
rect 6736 19456 6788 19508
rect 10692 19456 10744 19508
rect 10784 19456 10836 19508
rect 13084 19456 13136 19508
rect 13820 19499 13872 19508
rect 3608 19388 3660 19440
rect 3792 19388 3844 19440
rect 12440 19388 12492 19440
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 14372 19456 14424 19508
rect 15016 19456 15068 19508
rect 18052 19456 18104 19508
rect 18144 19456 18196 19508
rect 18972 19456 19024 19508
rect 19156 19456 19208 19508
rect 22836 19499 22888 19508
rect 15292 19388 15344 19440
rect 15844 19388 15896 19440
rect 17592 19388 17644 19440
rect 22836 19465 22845 19499
rect 22845 19465 22879 19499
rect 22879 19465 22888 19499
rect 22836 19456 22888 19465
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3056 19252 3108 19304
rect 3976 19363 4028 19372
rect 3976 19329 3985 19363
rect 3985 19329 4019 19363
rect 4019 19329 4028 19363
rect 3976 19320 4028 19329
rect 5632 19320 5684 19372
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6184 19295 6236 19304
rect 6184 19261 6193 19295
rect 6193 19261 6227 19295
rect 6227 19261 6236 19295
rect 7012 19320 7064 19372
rect 7840 19320 7892 19372
rect 8024 19320 8076 19372
rect 7656 19295 7708 19304
rect 6184 19252 6236 19261
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 14372 19320 14424 19372
rect 14740 19320 14792 19372
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 15752 19320 15804 19372
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 4068 19184 4120 19236
rect 2780 19116 2832 19168
rect 2872 19116 2924 19168
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3424 19159 3476 19168
rect 3056 19116 3108 19125
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 3608 19116 3660 19168
rect 4620 19116 4672 19168
rect 5172 19116 5224 19168
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 8208 19252 8260 19304
rect 6184 19116 6236 19168
rect 7012 19116 7064 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 9864 19184 9916 19236
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 11152 19252 11204 19304
rect 12532 19252 12584 19304
rect 14280 19252 14332 19304
rect 16304 19252 16356 19304
rect 16396 19252 16448 19304
rect 10968 19184 11020 19236
rect 11704 19227 11756 19236
rect 11704 19193 11713 19227
rect 11713 19193 11747 19227
rect 11747 19193 11756 19227
rect 11704 19184 11756 19193
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 9680 19116 9732 19125
rect 11152 19116 11204 19168
rect 11428 19159 11480 19168
rect 11428 19125 11437 19159
rect 11437 19125 11471 19159
rect 11471 19125 11480 19159
rect 11428 19116 11480 19125
rect 14004 19159 14056 19168
rect 14004 19125 14013 19159
rect 14013 19125 14047 19159
rect 14047 19125 14056 19159
rect 14004 19116 14056 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 16580 19184 16632 19236
rect 17960 19252 18012 19304
rect 22744 19388 22796 19440
rect 18972 19252 19024 19304
rect 20812 19252 20864 19304
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 17040 19116 17092 19168
rect 19340 19184 19392 19236
rect 20352 19184 20404 19236
rect 22284 19184 22336 19236
rect 23388 19252 23440 19304
rect 19524 19116 19576 19168
rect 21088 19159 21140 19168
rect 21088 19125 21097 19159
rect 21097 19125 21131 19159
rect 21131 19125 21140 19159
rect 21088 19116 21140 19125
rect 21640 19116 21692 19168
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 8446 19014 8498 19066
rect 8510 19014 8562 19066
rect 8574 19014 8626 19066
rect 8638 19014 8690 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 2872 18912 2924 18964
rect 3516 18912 3568 18964
rect 4620 18912 4672 18964
rect 6736 18912 6788 18964
rect 7012 18955 7064 18964
rect 7012 18921 7021 18955
rect 7021 18921 7055 18955
rect 7055 18921 7064 18955
rect 7012 18912 7064 18921
rect 8208 18912 8260 18964
rect 9956 18912 10008 18964
rect 12992 18955 13044 18964
rect 12992 18921 13001 18955
rect 13001 18921 13035 18955
rect 13035 18921 13044 18955
rect 12992 18912 13044 18921
rect 14464 18912 14516 18964
rect 15568 18912 15620 18964
rect 16580 18912 16632 18964
rect 19984 18912 20036 18964
rect 20352 18955 20404 18964
rect 20352 18921 20361 18955
rect 20361 18921 20395 18955
rect 20395 18921 20404 18955
rect 20352 18912 20404 18921
rect 22284 18955 22336 18964
rect 22284 18921 22293 18955
rect 22293 18921 22327 18955
rect 22327 18921 22336 18955
rect 22284 18912 22336 18921
rect 3424 18844 3476 18896
rect 1584 18776 1636 18828
rect 3056 18776 3108 18828
rect 3516 18819 3568 18828
rect 3516 18785 3525 18819
rect 3525 18785 3559 18819
rect 3559 18785 3568 18819
rect 3516 18776 3568 18785
rect 6828 18844 6880 18896
rect 9128 18844 9180 18896
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 8024 18776 8076 18828
rect 9220 18776 9272 18828
rect 9496 18776 9548 18828
rect 9680 18844 9732 18896
rect 11520 18776 11572 18828
rect 12532 18844 12584 18896
rect 14004 18844 14056 18896
rect 14280 18776 14332 18828
rect 14556 18819 14608 18828
rect 14556 18785 14565 18819
rect 14565 18785 14599 18819
rect 14599 18785 14608 18819
rect 14556 18776 14608 18785
rect 15476 18776 15528 18828
rect 3700 18751 3752 18760
rect 3700 18717 3709 18751
rect 3709 18717 3743 18751
rect 3743 18717 3752 18751
rect 3700 18708 3752 18717
rect 4252 18640 4304 18692
rect 5540 18708 5592 18760
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 7196 18640 7248 18692
rect 6184 18572 6236 18624
rect 7564 18708 7616 18760
rect 9588 18708 9640 18760
rect 8760 18640 8812 18692
rect 10048 18708 10100 18760
rect 10784 18708 10836 18760
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 15200 18640 15252 18692
rect 15568 18640 15620 18692
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 21088 18844 21140 18896
rect 18972 18819 19024 18828
rect 17316 18776 17368 18785
rect 18972 18785 18981 18819
rect 18981 18785 19015 18819
rect 19015 18785 19024 18819
rect 18972 18776 19024 18785
rect 19984 18776 20036 18828
rect 20996 18776 21048 18828
rect 16304 18708 16356 18760
rect 16856 18708 16908 18760
rect 17132 18708 17184 18760
rect 20812 18708 20864 18760
rect 22468 18708 22520 18760
rect 7656 18572 7708 18624
rect 9404 18572 9456 18624
rect 11796 18572 11848 18624
rect 12716 18572 12768 18624
rect 15108 18615 15160 18624
rect 15108 18581 15117 18615
rect 15117 18581 15151 18615
rect 15151 18581 15160 18615
rect 15108 18572 15160 18581
rect 22376 18683 22428 18692
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 22744 18572 22796 18624
rect 4714 18470 4766 18522
rect 4778 18470 4830 18522
rect 4842 18470 4894 18522
rect 4906 18470 4958 18522
rect 12178 18470 12230 18522
rect 12242 18470 12294 18522
rect 12306 18470 12358 18522
rect 12370 18470 12422 18522
rect 19642 18470 19694 18522
rect 19706 18470 19758 18522
rect 19770 18470 19822 18522
rect 19834 18470 19886 18522
rect 3056 18368 3108 18420
rect 3516 18368 3568 18420
rect 5172 18368 5224 18420
rect 10784 18411 10836 18420
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 3884 18164 3936 18216
rect 8024 18232 8076 18284
rect 4252 18096 4304 18148
rect 6184 18164 6236 18216
rect 7104 18207 7156 18216
rect 7104 18173 7138 18207
rect 7138 18173 7156 18207
rect 7104 18164 7156 18173
rect 8760 18164 8812 18216
rect 9312 18275 9364 18284
rect 9312 18241 9324 18275
rect 9324 18241 9358 18275
rect 9358 18241 9364 18275
rect 9312 18232 9364 18241
rect 10048 18232 10100 18284
rect 10784 18377 10793 18411
rect 10793 18377 10827 18411
rect 10827 18377 10836 18411
rect 10784 18368 10836 18377
rect 10968 18368 11020 18420
rect 14556 18368 14608 18420
rect 15292 18368 15344 18420
rect 10692 18300 10744 18352
rect 11244 18275 11296 18284
rect 11244 18241 11253 18275
rect 11253 18241 11287 18275
rect 11287 18241 11296 18275
rect 11244 18232 11296 18241
rect 11428 18300 11480 18352
rect 16396 18368 16448 18420
rect 9956 18164 10008 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 14372 18164 14424 18216
rect 15016 18164 15068 18216
rect 16396 18207 16448 18216
rect 16396 18173 16405 18207
rect 16405 18173 16439 18207
rect 16439 18173 16448 18207
rect 16396 18164 16448 18173
rect 18052 18232 18104 18284
rect 18972 18368 19024 18420
rect 19984 18411 20036 18420
rect 19984 18377 19993 18411
rect 19993 18377 20027 18411
rect 20027 18377 20036 18411
rect 19984 18368 20036 18377
rect 20076 18411 20128 18420
rect 20076 18377 20085 18411
rect 20085 18377 20119 18411
rect 20119 18377 20128 18411
rect 20076 18368 20128 18377
rect 20628 18368 20680 18420
rect 22376 18368 22428 18420
rect 20444 18300 20496 18352
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 20352 18164 20404 18216
rect 7564 18096 7616 18148
rect 8024 18096 8076 18148
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 6276 18028 6328 18080
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 9128 18028 9180 18080
rect 9496 18028 9548 18080
rect 12532 18028 12584 18080
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 14004 18096 14056 18148
rect 15660 18096 15712 18148
rect 19524 18096 19576 18148
rect 20812 18096 20864 18148
rect 21456 18164 21508 18216
rect 21640 18207 21692 18216
rect 21640 18173 21674 18207
rect 21674 18173 21692 18207
rect 21640 18164 21692 18173
rect 21916 18164 21968 18216
rect 23112 18164 23164 18216
rect 12900 18028 12952 18037
rect 14096 18028 14148 18080
rect 14464 18028 14516 18080
rect 16672 18028 16724 18080
rect 22468 18096 22520 18148
rect 21824 18028 21876 18080
rect 8446 17926 8498 17978
rect 8510 17926 8562 17978
rect 8574 17926 8626 17978
rect 8638 17926 8690 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 7748 17824 7800 17876
rect 9588 17824 9640 17876
rect 10048 17867 10100 17876
rect 10048 17833 10057 17867
rect 10057 17833 10091 17867
rect 10091 17833 10100 17867
rect 10048 17824 10100 17833
rect 12900 17824 12952 17876
rect 14004 17867 14056 17876
rect 14004 17833 14013 17867
rect 14013 17833 14047 17867
rect 14047 17833 14056 17867
rect 14004 17824 14056 17833
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14464 17867 14516 17876
rect 14096 17824 14148 17833
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 15016 17824 15068 17876
rect 16672 17867 16724 17876
rect 16672 17833 16681 17867
rect 16681 17833 16715 17867
rect 16715 17833 16724 17867
rect 16672 17824 16724 17833
rect 17132 17824 17184 17876
rect 19432 17867 19484 17876
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 19524 17824 19576 17876
rect 1768 17756 1820 17808
rect 3240 17756 3292 17808
rect 3884 17756 3936 17808
rect 4620 17756 4672 17808
rect 3332 17688 3384 17740
rect 5724 17756 5776 17808
rect 6184 17756 6236 17808
rect 8576 17756 8628 17808
rect 9036 17756 9088 17808
rect 12072 17756 12124 17808
rect 9128 17688 9180 17740
rect 9680 17688 9732 17740
rect 15476 17756 15528 17808
rect 18420 17756 18472 17808
rect 21180 17756 21232 17808
rect 21732 17824 21784 17876
rect 21824 17799 21876 17808
rect 21824 17765 21858 17799
rect 21858 17765 21876 17799
rect 21824 17756 21876 17765
rect 13820 17688 13872 17740
rect 15108 17731 15160 17740
rect 15108 17697 15117 17731
rect 15117 17697 15151 17731
rect 15151 17697 15160 17731
rect 15108 17688 15160 17697
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 16396 17688 16448 17740
rect 18052 17688 18104 17740
rect 19432 17688 19484 17740
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 3148 17620 3200 17672
rect 3608 17620 3660 17672
rect 6920 17620 6972 17672
rect 8208 17620 8260 17672
rect 8944 17552 8996 17604
rect 3608 17484 3660 17536
rect 6184 17527 6236 17536
rect 6184 17493 6193 17527
rect 6193 17493 6227 17527
rect 6227 17493 6236 17527
rect 6184 17484 6236 17493
rect 8116 17484 8168 17536
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 12440 17663 12492 17672
rect 12440 17629 12449 17663
rect 12449 17629 12483 17663
rect 12483 17629 12492 17663
rect 12440 17620 12492 17629
rect 14648 17663 14700 17672
rect 9404 17484 9456 17536
rect 10048 17484 10100 17536
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 17868 17620 17920 17672
rect 17040 17552 17092 17604
rect 19340 17595 19392 17604
rect 19340 17561 19349 17595
rect 19349 17561 19383 17595
rect 19383 17561 19392 17595
rect 20168 17620 20220 17672
rect 20628 17620 20680 17672
rect 21456 17620 21508 17672
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 19340 17552 19392 17561
rect 13268 17484 13320 17536
rect 20444 17527 20496 17536
rect 20444 17493 20453 17527
rect 20453 17493 20487 17527
rect 20487 17493 20496 17527
rect 20444 17484 20496 17493
rect 22836 17484 22888 17536
rect 4714 17382 4766 17434
rect 4778 17382 4830 17434
rect 4842 17382 4894 17434
rect 4906 17382 4958 17434
rect 12178 17382 12230 17434
rect 12242 17382 12294 17434
rect 12306 17382 12358 17434
rect 12370 17382 12422 17434
rect 19642 17382 19694 17434
rect 19706 17382 19758 17434
rect 19770 17382 19822 17434
rect 19834 17382 19886 17434
rect 4252 17280 4304 17332
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 6368 17280 6420 17332
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 8576 17280 8628 17332
rect 9496 17280 9548 17332
rect 9772 17280 9824 17332
rect 10968 17280 11020 17332
rect 12072 17323 12124 17332
rect 12072 17289 12081 17323
rect 12081 17289 12115 17323
rect 12115 17289 12124 17323
rect 12072 17280 12124 17289
rect 12716 17280 12768 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 15476 17280 15528 17332
rect 19432 17323 19484 17332
rect 19432 17289 19441 17323
rect 19441 17289 19475 17323
rect 19475 17289 19484 17323
rect 19432 17280 19484 17289
rect 21364 17280 21416 17332
rect 1584 17144 1636 17196
rect 3240 17144 3292 17196
rect 4620 17144 4672 17196
rect 3608 17119 3660 17128
rect 3608 17085 3642 17119
rect 3642 17085 3660 17119
rect 3608 17076 3660 17085
rect 3056 17008 3108 17060
rect 7012 17144 7064 17196
rect 18052 17187 18104 17196
rect 5632 17076 5684 17128
rect 6184 17076 6236 17128
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 9772 17076 9824 17128
rect 9864 17076 9916 17128
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 18052 17153 18061 17187
rect 18061 17153 18095 17187
rect 18095 17153 18104 17187
rect 18052 17144 18104 17153
rect 11244 17076 11296 17128
rect 12716 17119 12768 17128
rect 12716 17085 12750 17119
rect 12750 17085 12768 17119
rect 5264 17008 5316 17060
rect 3424 16940 3476 16992
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 6276 16940 6328 16992
rect 8300 17008 8352 17060
rect 8944 17008 8996 17060
rect 10140 17008 10192 17060
rect 9864 16940 9916 16992
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 11060 17008 11112 17060
rect 12716 17076 12768 17085
rect 13268 17076 13320 17128
rect 13544 17076 13596 17128
rect 15292 17076 15344 17128
rect 20168 17187 20220 17196
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 22192 17212 22244 17264
rect 22376 17144 22428 17196
rect 22468 17144 22520 17196
rect 20444 17076 20496 17128
rect 21824 17076 21876 17128
rect 22744 17119 22796 17128
rect 22744 17085 22753 17119
rect 22753 17085 22787 17119
rect 22787 17085 22796 17119
rect 22744 17076 22796 17085
rect 12532 17008 12584 17060
rect 14464 17008 14516 17060
rect 19064 17008 19116 17060
rect 10324 16940 10376 16949
rect 12716 16940 12768 16992
rect 19708 16940 19760 16992
rect 21548 17008 21600 17060
rect 21640 17008 21692 17060
rect 20996 16983 21048 16992
rect 20996 16949 21005 16983
rect 21005 16949 21039 16983
rect 21039 16949 21048 16983
rect 20996 16940 21048 16949
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 8446 16838 8498 16890
rect 8510 16838 8562 16890
rect 8574 16838 8626 16890
rect 8638 16838 8690 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 3056 16779 3108 16788
rect 3056 16745 3065 16779
rect 3065 16745 3099 16779
rect 3099 16745 3108 16779
rect 3056 16736 3108 16745
rect 4068 16736 4120 16788
rect 4712 16736 4764 16788
rect 6460 16736 6512 16788
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 8208 16736 8260 16788
rect 11060 16736 11112 16788
rect 11244 16736 11296 16788
rect 19064 16779 19116 16788
rect 2688 16668 2740 16720
rect 6184 16668 6236 16720
rect 1584 16600 1636 16652
rect 3148 16600 3200 16652
rect 3516 16643 3568 16652
rect 3516 16609 3525 16643
rect 3525 16609 3559 16643
rect 3559 16609 3568 16643
rect 3516 16600 3568 16609
rect 3700 16575 3752 16584
rect 3700 16541 3709 16575
rect 3709 16541 3743 16575
rect 3743 16541 3752 16575
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 6368 16600 6420 16652
rect 7196 16643 7248 16652
rect 7196 16609 7230 16643
rect 7230 16609 7248 16643
rect 7196 16600 7248 16609
rect 3700 16532 3752 16541
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 6184 16507 6236 16516
rect 6184 16473 6193 16507
rect 6193 16473 6227 16507
rect 6227 16473 6236 16507
rect 6184 16464 6236 16473
rect 8852 16668 8904 16720
rect 14096 16668 14148 16720
rect 15108 16668 15160 16720
rect 16212 16668 16264 16720
rect 19064 16745 19073 16779
rect 19073 16745 19107 16779
rect 19107 16745 19116 16779
rect 19064 16736 19116 16745
rect 22468 16736 22520 16788
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 9036 16600 9088 16652
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 13544 16643 13596 16652
rect 13544 16609 13553 16643
rect 13553 16609 13587 16643
rect 13587 16609 13596 16643
rect 13544 16600 13596 16609
rect 14188 16600 14240 16652
rect 17224 16600 17276 16652
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 18052 16668 18104 16720
rect 18696 16668 18748 16720
rect 19708 16668 19760 16720
rect 21732 16668 21784 16720
rect 19432 16600 19484 16652
rect 21180 16643 21232 16652
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 21456 16600 21508 16652
rect 8852 16575 8904 16584
rect 8852 16541 8861 16575
rect 8861 16541 8895 16575
rect 8895 16541 8904 16575
rect 8852 16532 8904 16541
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 9772 16575 9824 16584
rect 8944 16532 8996 16541
rect 9772 16541 9781 16575
rect 9781 16541 9815 16575
rect 9815 16541 9824 16575
rect 9772 16532 9824 16541
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 15292 16532 15344 16584
rect 19340 16532 19392 16584
rect 20168 16532 20220 16584
rect 12716 16464 12768 16516
rect 5816 16396 5868 16448
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 11888 16396 11940 16448
rect 20260 16464 20312 16516
rect 15200 16396 15252 16448
rect 17040 16439 17092 16448
rect 17040 16405 17049 16439
rect 17049 16405 17083 16439
rect 17083 16405 17092 16439
rect 17040 16396 17092 16405
rect 20904 16396 20956 16448
rect 21916 16396 21968 16448
rect 22928 16439 22980 16448
rect 22928 16405 22937 16439
rect 22937 16405 22971 16439
rect 22971 16405 22980 16439
rect 22928 16396 22980 16405
rect 4714 16294 4766 16346
rect 4778 16294 4830 16346
rect 4842 16294 4894 16346
rect 4906 16294 4958 16346
rect 12178 16294 12230 16346
rect 12242 16294 12294 16346
rect 12306 16294 12358 16346
rect 12370 16294 12422 16346
rect 19642 16294 19694 16346
rect 19706 16294 19758 16346
rect 19770 16294 19822 16346
rect 19834 16294 19886 16346
rect 3332 16192 3384 16244
rect 3792 16192 3844 16244
rect 8024 16192 8076 16244
rect 8852 16192 8904 16244
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 11796 16192 11848 16244
rect 14924 16192 14976 16244
rect 17316 16192 17368 16244
rect 19432 16235 19484 16244
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 21180 16235 21232 16244
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 3700 16124 3752 16176
rect 4620 16056 4672 16108
rect 5816 16056 5868 16108
rect 1676 15988 1728 16040
rect 2044 16031 2096 16040
rect 2044 15997 2053 16031
rect 2053 15997 2087 16031
rect 2087 15997 2096 16031
rect 2044 15988 2096 15997
rect 3516 15988 3568 16040
rect 3608 15988 3660 16040
rect 5080 15988 5132 16040
rect 5356 15988 5408 16040
rect 6552 16056 6604 16108
rect 5724 15920 5776 15972
rect 6644 15988 6696 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 8300 16056 8352 16108
rect 7380 15988 7432 16040
rect 8760 15988 8812 16040
rect 9864 16056 9916 16108
rect 10048 16056 10100 16108
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 6920 15920 6972 15972
rect 8392 15920 8444 15972
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 7196 15852 7248 15904
rect 8852 15920 8904 15972
rect 11060 15988 11112 16040
rect 14188 16056 14240 16108
rect 14556 16056 14608 16108
rect 15660 16099 15712 16108
rect 15660 16065 15672 16099
rect 15672 16065 15706 16099
rect 15706 16065 15712 16099
rect 15660 16056 15712 16065
rect 17040 16056 17092 16108
rect 20168 16099 20220 16108
rect 20168 16065 20177 16099
rect 20177 16065 20211 16099
rect 20211 16065 20220 16099
rect 20168 16056 20220 16065
rect 20904 16099 20956 16108
rect 20904 16065 20913 16099
rect 20913 16065 20947 16099
rect 20947 16065 20956 16099
rect 20904 16056 20956 16065
rect 12072 15988 12124 16040
rect 12532 15988 12584 16040
rect 15292 15988 15344 16040
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 10324 15852 10376 15904
rect 11980 15920 12032 15972
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14188 15852 14240 15904
rect 15200 15852 15252 15904
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17684 15920 17736 15972
rect 20352 15988 20404 16040
rect 19340 15920 19392 15972
rect 22376 16192 22428 16244
rect 21640 16099 21692 16108
rect 21640 16065 21649 16099
rect 21649 16065 21683 16099
rect 21683 16065 21692 16099
rect 21640 16056 21692 16065
rect 22284 16056 22336 16108
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22928 16056 22980 16108
rect 17132 15852 17184 15861
rect 19892 15895 19944 15904
rect 19892 15861 19901 15895
rect 19901 15861 19935 15895
rect 19935 15861 19944 15895
rect 19892 15852 19944 15861
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 20444 15852 20496 15904
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 21548 15895 21600 15904
rect 21548 15861 21557 15895
rect 21557 15861 21591 15895
rect 21591 15861 21600 15895
rect 21548 15852 21600 15861
rect 22192 15852 22244 15904
rect 8446 15750 8498 15802
rect 8510 15750 8562 15802
rect 8574 15750 8626 15802
rect 8638 15750 8690 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 1676 15512 1728 15564
rect 3056 15512 3108 15564
rect 3424 15555 3476 15564
rect 3424 15521 3433 15555
rect 3433 15521 3467 15555
rect 3467 15521 3476 15555
rect 3424 15512 3476 15521
rect 2964 15444 3016 15496
rect 4528 15580 4580 15632
rect 7472 15648 7524 15700
rect 9036 15691 9088 15700
rect 9036 15657 9045 15691
rect 9045 15657 9079 15691
rect 9079 15657 9088 15691
rect 9036 15648 9088 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10324 15648 10376 15700
rect 11980 15648 12032 15700
rect 12716 15691 12768 15700
rect 12716 15657 12731 15691
rect 12731 15657 12765 15691
rect 12765 15657 12768 15691
rect 14188 15691 14240 15700
rect 12716 15648 12768 15657
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 7196 15580 7248 15632
rect 8300 15580 8352 15632
rect 4620 15512 4672 15564
rect 5264 15512 5316 15564
rect 6368 15512 6420 15564
rect 9220 15512 9272 15564
rect 9404 15512 9456 15564
rect 10048 15512 10100 15564
rect 11060 15555 11112 15564
rect 11060 15521 11094 15555
rect 11094 15521 11112 15555
rect 11060 15512 11112 15521
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 7012 15444 7064 15496
rect 2780 15308 2832 15360
rect 3516 15308 3568 15360
rect 5264 15308 5316 15360
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 8944 15419 8996 15428
rect 8944 15385 8953 15419
rect 8953 15385 8987 15419
rect 8987 15385 8996 15419
rect 8944 15376 8996 15385
rect 9772 15376 9824 15428
rect 11888 15512 11940 15564
rect 12440 15444 12492 15496
rect 13452 15444 13504 15496
rect 11428 15308 11480 15360
rect 12072 15308 12124 15360
rect 13820 15376 13872 15428
rect 13912 15308 13964 15360
rect 15292 15648 15344 15700
rect 19340 15648 19392 15700
rect 17040 15580 17092 15632
rect 19892 15580 19944 15632
rect 20996 15648 21048 15700
rect 22560 15648 22612 15700
rect 22928 15580 22980 15632
rect 16396 15512 16448 15564
rect 17224 15555 17276 15564
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 18052 15512 18104 15564
rect 18512 15512 18564 15564
rect 19984 15512 20036 15564
rect 20444 15555 20496 15564
rect 20444 15521 20453 15555
rect 20453 15521 20487 15555
rect 20487 15521 20496 15555
rect 20444 15512 20496 15521
rect 23112 15512 23164 15564
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 17592 15308 17644 15360
rect 17684 15308 17736 15360
rect 19340 15308 19392 15360
rect 22376 15308 22428 15360
rect 4714 15206 4766 15258
rect 4778 15206 4830 15258
rect 4842 15206 4894 15258
rect 4906 15206 4958 15258
rect 12178 15206 12230 15258
rect 12242 15206 12294 15258
rect 12306 15206 12358 15258
rect 12370 15206 12422 15258
rect 19642 15206 19694 15258
rect 19706 15206 19758 15258
rect 19770 15206 19822 15258
rect 19834 15206 19886 15258
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 6460 15147 6512 15156
rect 6460 15113 6469 15147
rect 6469 15113 6503 15147
rect 6503 15113 6512 15147
rect 7656 15147 7708 15156
rect 6460 15104 6512 15113
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 7656 15104 7708 15113
rect 8760 15104 8812 15156
rect 4620 15036 4672 15088
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 1768 14900 1820 14952
rect 2044 14943 2096 14952
rect 2044 14909 2053 14943
rect 2053 14909 2087 14943
rect 2087 14909 2096 14943
rect 2044 14900 2096 14909
rect 4068 14900 4120 14952
rect 5264 14943 5316 14952
rect 5264 14909 5298 14943
rect 5298 14909 5316 14943
rect 5264 14900 5316 14909
rect 8024 14943 8076 14952
rect 3148 14832 3200 14884
rect 4436 14832 4488 14884
rect 5172 14832 5224 14884
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 9128 15104 9180 15156
rect 10508 15104 10560 15156
rect 11060 15104 11112 15156
rect 12532 15104 12584 15156
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 9680 14900 9732 14952
rect 11336 14900 11388 14952
rect 12624 15036 12676 15088
rect 16212 15036 16264 15088
rect 15384 14968 15436 15020
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 16672 14968 16724 15020
rect 10416 14875 10468 14884
rect 10416 14841 10450 14875
rect 10450 14841 10468 14875
rect 10416 14832 10468 14841
rect 11980 14875 12032 14884
rect 11980 14841 11989 14875
rect 11989 14841 12023 14875
rect 12023 14841 12032 14875
rect 11980 14832 12032 14841
rect 13268 14900 13320 14952
rect 13820 14900 13872 14952
rect 16764 14900 16816 14952
rect 19340 15104 19392 15156
rect 19984 15104 20036 15156
rect 20812 15104 20864 15156
rect 22284 15104 22336 15156
rect 17960 15036 18012 15088
rect 18604 15036 18656 15088
rect 18696 15011 18748 15020
rect 18696 14977 18705 15011
rect 18705 14977 18739 15011
rect 18739 14977 18748 15011
rect 18696 14968 18748 14977
rect 20168 14968 20220 15020
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 21364 14943 21416 14952
rect 21364 14909 21373 14943
rect 21373 14909 21407 14943
rect 21407 14909 21416 14943
rect 21364 14900 21416 14909
rect 22376 14900 22428 14952
rect 22836 14943 22888 14952
rect 22836 14909 22845 14943
rect 22845 14909 22879 14943
rect 22879 14909 22888 14943
rect 22836 14900 22888 14909
rect 14464 14832 14516 14884
rect 7012 14764 7064 14816
rect 7472 14764 7524 14816
rect 9404 14764 9456 14816
rect 9864 14764 9916 14816
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 15660 14832 15712 14884
rect 17132 14832 17184 14884
rect 14740 14764 14792 14816
rect 15108 14807 15160 14816
rect 15108 14773 15117 14807
rect 15117 14773 15151 14807
rect 15151 14773 15160 14807
rect 16488 14807 16540 14816
rect 15108 14764 15160 14773
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 17224 14764 17276 14816
rect 18788 14832 18840 14884
rect 19800 14832 19852 14884
rect 19340 14764 19392 14816
rect 19432 14764 19484 14816
rect 22284 14764 22336 14816
rect 22928 14764 22980 14816
rect 8446 14662 8498 14714
rect 8510 14662 8562 14714
rect 8574 14662 8626 14714
rect 8638 14662 8690 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 3424 14560 3476 14612
rect 4436 14603 4488 14612
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 5080 14560 5132 14612
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 6368 14560 6420 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10416 14560 10468 14612
rect 2780 14492 2832 14544
rect 4620 14492 4672 14544
rect 6920 14492 6972 14544
rect 8116 14492 8168 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 7380 14424 7432 14476
rect 9772 14424 9824 14476
rect 12716 14560 12768 14612
rect 15660 14603 15712 14612
rect 10324 14424 10376 14476
rect 6552 14356 6604 14408
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 10876 14424 10928 14476
rect 14556 14492 14608 14544
rect 15108 14492 15160 14544
rect 11428 14424 11480 14476
rect 11980 14424 12032 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 17040 14560 17092 14612
rect 19800 14603 19852 14612
rect 16396 14424 16448 14476
rect 16580 14467 16632 14476
rect 16580 14433 16614 14467
rect 16614 14433 16632 14467
rect 19340 14492 19392 14544
rect 19800 14569 19809 14603
rect 19809 14569 19843 14603
rect 19843 14569 19852 14603
rect 19800 14560 19852 14569
rect 20260 14603 20312 14612
rect 20260 14569 20269 14603
rect 20269 14569 20303 14603
rect 20303 14569 20312 14603
rect 20260 14560 20312 14569
rect 16580 14424 16632 14433
rect 18236 14424 18288 14476
rect 18512 14424 18564 14476
rect 19432 14424 19484 14476
rect 21548 14424 21600 14476
rect 22928 14424 22980 14476
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 5356 14288 5408 14340
rect 15660 14288 15712 14340
rect 16212 14356 16264 14408
rect 17316 14288 17368 14340
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 9404 14220 9456 14272
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 14004 14220 14056 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 17040 14220 17092 14272
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 17868 14220 17920 14272
rect 18604 14220 18656 14272
rect 21364 14356 21416 14408
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 20536 14220 20588 14272
rect 22652 14220 22704 14272
rect 4714 14118 4766 14170
rect 4778 14118 4830 14170
rect 4842 14118 4894 14170
rect 4906 14118 4958 14170
rect 12178 14118 12230 14170
rect 12242 14118 12294 14170
rect 12306 14118 12358 14170
rect 12370 14118 12422 14170
rect 19642 14118 19694 14170
rect 19706 14118 19758 14170
rect 19770 14118 19822 14170
rect 19834 14118 19886 14170
rect 1768 14016 1820 14068
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 5172 14016 5224 14068
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 11796 14016 11848 14068
rect 13452 14059 13504 14068
rect 3056 13948 3108 14000
rect 3608 13923 3660 13932
rect 3608 13889 3617 13923
rect 3617 13889 3651 13923
rect 3651 13889 3660 13923
rect 3608 13880 3660 13889
rect 4528 13880 4580 13932
rect 6736 13948 6788 14000
rect 10140 13948 10192 14000
rect 10324 13948 10376 14000
rect 5540 13880 5592 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 10876 13880 10928 13932
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 8668 13812 8720 13864
rect 9680 13812 9732 13864
rect 9956 13812 10008 13864
rect 11336 13812 11388 13864
rect 11428 13812 11480 13864
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 14464 14016 14516 14068
rect 15016 14016 15068 14068
rect 17960 14016 18012 14068
rect 18052 14016 18104 14068
rect 19432 14059 19484 14068
rect 12624 13880 12676 13932
rect 17776 13948 17828 14000
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 20444 14016 20496 14068
rect 23112 13948 23164 14000
rect 14740 13880 14792 13932
rect 2688 13744 2740 13796
rect 2780 13744 2832 13796
rect 3516 13744 3568 13796
rect 6092 13744 6144 13796
rect 6276 13787 6328 13796
rect 6276 13753 6285 13787
rect 6285 13753 6319 13787
rect 6319 13753 6328 13787
rect 6276 13744 6328 13753
rect 10692 13744 10744 13796
rect 12624 13744 12676 13796
rect 12900 13787 12952 13796
rect 12900 13753 12909 13787
rect 12909 13753 12943 13787
rect 12943 13753 12952 13787
rect 12900 13744 12952 13753
rect 15292 13744 15344 13796
rect 16488 13812 16540 13864
rect 17592 13812 17644 13864
rect 18328 13855 18380 13864
rect 18328 13821 18362 13855
rect 18362 13821 18380 13855
rect 16396 13744 16448 13796
rect 18328 13812 18380 13821
rect 20260 13880 20312 13932
rect 20536 13880 20588 13932
rect 22192 13880 22244 13932
rect 20076 13812 20128 13864
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 22468 13812 22520 13864
rect 18512 13744 18564 13796
rect 19616 13744 19668 13796
rect 4068 13676 4120 13728
rect 5264 13676 5316 13728
rect 6184 13676 6236 13728
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 8760 13719 8812 13728
rect 6368 13676 6420 13685
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 10416 13676 10468 13728
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 13360 13676 13412 13728
rect 17040 13719 17092 13728
rect 17040 13685 17049 13719
rect 17049 13685 17083 13719
rect 17083 13685 17092 13719
rect 17040 13676 17092 13685
rect 17316 13719 17368 13728
rect 17316 13685 17325 13719
rect 17325 13685 17359 13719
rect 17359 13685 17368 13719
rect 17316 13676 17368 13685
rect 20260 13676 20312 13728
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 8446 13574 8498 13626
rect 8510 13574 8562 13626
rect 8574 13574 8626 13626
rect 8638 13574 8690 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 3516 13472 3568 13524
rect 4068 13515 4120 13524
rect 4068 13481 4077 13515
rect 4077 13481 4111 13515
rect 4111 13481 4120 13515
rect 4068 13472 4120 13481
rect 6828 13472 6880 13524
rect 10140 13515 10192 13524
rect 3424 13404 3476 13456
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3976 13268 4028 13320
rect 5448 13404 5500 13456
rect 6736 13404 6788 13456
rect 8760 13404 8812 13456
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 10876 13472 10928 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 16580 13472 16632 13524
rect 16948 13472 17000 13524
rect 18512 13472 18564 13524
rect 18880 13472 18932 13524
rect 19248 13472 19300 13524
rect 5080 13336 5132 13388
rect 6092 13336 6144 13388
rect 6184 13336 6236 13388
rect 12440 13404 12492 13456
rect 13360 13404 13412 13456
rect 17684 13404 17736 13456
rect 20536 13472 20588 13524
rect 20444 13447 20496 13456
rect 10508 13379 10560 13388
rect 7380 13311 7432 13320
rect 3608 13200 3660 13252
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 8944 13268 8996 13320
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 11888 13336 11940 13388
rect 12992 13336 13044 13388
rect 14372 13336 14424 13388
rect 14464 13336 14516 13388
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 15384 13336 15436 13388
rect 15844 13336 15896 13388
rect 20444 13413 20453 13447
rect 20453 13413 20487 13447
rect 20487 13413 20496 13447
rect 20444 13404 20496 13413
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 10692 13268 10744 13320
rect 12348 13268 12400 13320
rect 4528 13132 4580 13184
rect 9864 13200 9916 13252
rect 11980 13200 12032 13252
rect 12532 13200 12584 13252
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 8760 13175 8812 13184
rect 8760 13141 8769 13175
rect 8769 13141 8803 13175
rect 8803 13141 8812 13175
rect 8760 13132 8812 13141
rect 10600 13132 10652 13184
rect 14832 13200 14884 13252
rect 16212 13132 16264 13184
rect 17960 13132 18012 13184
rect 20352 13336 20404 13388
rect 22560 13472 22612 13524
rect 22652 13404 22704 13456
rect 23112 13404 23164 13456
rect 20720 13336 20772 13388
rect 22008 13336 22060 13388
rect 20904 13311 20956 13320
rect 18512 13132 18564 13184
rect 19524 13132 19576 13184
rect 20168 13132 20220 13184
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 20812 13132 20864 13184
rect 22468 13132 22520 13184
rect 4714 13030 4766 13082
rect 4778 13030 4830 13082
rect 4842 13030 4894 13082
rect 4906 13030 4958 13082
rect 12178 13030 12230 13082
rect 12242 13030 12294 13082
rect 12306 13030 12358 13082
rect 12370 13030 12422 13082
rect 19642 13030 19694 13082
rect 19706 13030 19758 13082
rect 19770 13030 19822 13082
rect 19834 13030 19886 13082
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 4068 12903 4120 12912
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 5080 12928 5132 12980
rect 6092 12971 6144 12980
rect 6092 12937 6101 12971
rect 6101 12937 6135 12971
rect 6135 12937 6144 12971
rect 6092 12928 6144 12937
rect 4068 12860 4120 12869
rect 2044 12724 2096 12776
rect 3424 12656 3476 12708
rect 4068 12588 4120 12640
rect 5264 12724 5316 12776
rect 9128 12928 9180 12980
rect 9772 12928 9824 12980
rect 8944 12860 8996 12912
rect 9404 12860 9456 12912
rect 10968 12928 11020 12980
rect 11888 12928 11940 12980
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 15752 12928 15804 12980
rect 16856 12928 16908 12980
rect 17592 12928 17644 12980
rect 20352 12928 20404 12980
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7380 12724 7432 12776
rect 8760 12724 8812 12776
rect 10692 12724 10744 12776
rect 11796 12792 11848 12844
rect 12992 12835 13044 12844
rect 11704 12724 11756 12776
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 14004 12792 14056 12844
rect 17224 12860 17276 12912
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 16396 12792 16448 12844
rect 17868 12860 17920 12912
rect 20168 12835 20220 12844
rect 20168 12801 20177 12835
rect 20177 12801 20211 12835
rect 20211 12801 20220 12835
rect 20168 12792 20220 12801
rect 20444 12792 20496 12844
rect 7012 12588 7064 12597
rect 8300 12588 8352 12640
rect 9772 12656 9824 12708
rect 12072 12656 12124 12708
rect 9864 12588 9916 12640
rect 10600 12588 10652 12640
rect 16580 12724 16632 12776
rect 17960 12724 18012 12776
rect 14648 12656 14700 12708
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 14832 12656 14884 12665
rect 17684 12656 17736 12708
rect 19524 12724 19576 12776
rect 20904 12928 20956 12980
rect 21180 12928 21232 12980
rect 23296 12928 23348 12980
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 22652 12835 22704 12844
rect 22652 12801 22661 12835
rect 22661 12801 22695 12835
rect 22695 12801 22704 12835
rect 22652 12792 22704 12801
rect 18512 12656 18564 12708
rect 20812 12767 20864 12776
rect 20812 12733 20846 12767
rect 20846 12733 20864 12767
rect 20812 12724 20864 12733
rect 22744 12724 22796 12776
rect 20444 12656 20496 12708
rect 20996 12656 21048 12708
rect 13912 12588 13964 12640
rect 15108 12588 15160 12640
rect 17040 12588 17092 12640
rect 19616 12588 19668 12640
rect 21824 12588 21876 12640
rect 22744 12588 22796 12640
rect 23112 12588 23164 12640
rect 8446 12486 8498 12538
rect 8510 12486 8562 12538
rect 8574 12486 8626 12538
rect 8638 12486 8690 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 5264 12384 5316 12436
rect 6276 12384 6328 12436
rect 9036 12384 9088 12436
rect 10048 12384 10100 12436
rect 10140 12384 10192 12436
rect 10692 12384 10744 12436
rect 12072 12384 12124 12436
rect 14648 12384 14700 12436
rect 15108 12384 15160 12436
rect 15568 12384 15620 12436
rect 16212 12384 16264 12436
rect 2780 12316 2832 12368
rect 3332 12316 3384 12368
rect 4436 12316 4488 12368
rect 6368 12316 6420 12368
rect 8300 12316 8352 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 8208 12248 8260 12300
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 11520 12248 11572 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 6920 12180 6972 12232
rect 8300 12112 8352 12164
rect 9404 12180 9456 12232
rect 14280 12248 14332 12300
rect 15016 12316 15068 12368
rect 16672 12316 16724 12368
rect 16488 12248 16540 12300
rect 17316 12384 17368 12436
rect 23020 12384 23072 12436
rect 17132 12316 17184 12368
rect 20444 12359 20496 12368
rect 20444 12325 20453 12359
rect 20453 12325 20487 12359
rect 20487 12325 20496 12359
rect 20444 12316 20496 12325
rect 20996 12316 21048 12368
rect 21824 12316 21876 12368
rect 23204 12316 23256 12368
rect 19248 12248 19300 12300
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 22928 12248 22980 12300
rect 9772 12112 9824 12164
rect 3148 12044 3200 12096
rect 12624 12180 12676 12232
rect 12992 12180 13044 12232
rect 15660 12180 15712 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 17776 12223 17828 12232
rect 15384 12112 15436 12164
rect 15476 12112 15528 12164
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 17960 12180 18012 12232
rect 18236 12180 18288 12232
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 19524 12223 19576 12232
rect 18788 12180 18840 12189
rect 19524 12189 19533 12223
rect 19533 12189 19567 12223
rect 19567 12189 19576 12223
rect 19524 12180 19576 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 20536 12223 20588 12232
rect 19616 12180 19668 12189
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 20904 12180 20956 12232
rect 19340 12112 19392 12164
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 17132 12044 17184 12096
rect 18052 12044 18104 12096
rect 18972 12044 19024 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 22652 12044 22704 12096
rect 4714 11942 4766 11994
rect 4778 11942 4830 11994
rect 4842 11942 4894 11994
rect 4906 11942 4958 11994
rect 12178 11942 12230 11994
rect 12242 11942 12294 11994
rect 12306 11942 12358 11994
rect 12370 11942 12422 11994
rect 19642 11942 19694 11994
rect 19706 11942 19758 11994
rect 19770 11942 19822 11994
rect 19834 11942 19886 11994
rect 4436 11840 4488 11892
rect 8760 11840 8812 11892
rect 10324 11840 10376 11892
rect 11520 11840 11572 11892
rect 12624 11883 12676 11892
rect 12624 11849 12633 11883
rect 12633 11849 12667 11883
rect 12667 11849 12676 11883
rect 12624 11840 12676 11849
rect 2044 11704 2096 11756
rect 3976 11636 4028 11688
rect 6920 11636 6972 11688
rect 10140 11704 10192 11756
rect 9680 11636 9732 11688
rect 14096 11840 14148 11892
rect 14280 11883 14332 11892
rect 14280 11849 14289 11883
rect 14289 11849 14323 11883
rect 14323 11849 14332 11883
rect 14280 11840 14332 11849
rect 15476 11883 15528 11892
rect 15476 11849 15485 11883
rect 15485 11849 15519 11883
rect 15519 11849 15528 11883
rect 15476 11840 15528 11849
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 19432 11840 19484 11892
rect 20444 11840 20496 11892
rect 12900 11679 12952 11688
rect 12900 11645 12909 11679
rect 12909 11645 12943 11679
rect 12943 11645 12952 11679
rect 15384 11772 15436 11824
rect 17960 11772 18012 11824
rect 22008 11815 22060 11824
rect 22008 11781 22017 11815
rect 22017 11781 22051 11815
rect 22051 11781 22060 11815
rect 22008 11772 22060 11781
rect 15200 11704 15252 11756
rect 16396 11704 16448 11756
rect 19248 11704 19300 11756
rect 12900 11636 12952 11645
rect 15568 11636 15620 11688
rect 8208 11568 8260 11620
rect 9312 11568 9364 11620
rect 11796 11568 11848 11620
rect 14188 11568 14240 11620
rect 14924 11568 14976 11620
rect 15752 11568 15804 11620
rect 16120 11636 16172 11688
rect 17132 11636 17184 11688
rect 17960 11636 18012 11688
rect 19340 11636 19392 11688
rect 19984 11704 20036 11756
rect 20720 11704 20772 11756
rect 22376 11704 22428 11756
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 22928 11747 22980 11756
rect 22928 11713 22937 11747
rect 22937 11713 22971 11747
rect 22971 11713 22980 11747
rect 22928 11704 22980 11713
rect 20076 11636 20128 11688
rect 20260 11636 20312 11688
rect 16396 11568 16448 11620
rect 18696 11568 18748 11620
rect 22744 11636 22796 11688
rect 21640 11568 21692 11620
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 14556 11500 14608 11552
rect 16212 11500 16264 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 19064 11500 19116 11552
rect 19892 11500 19944 11552
rect 8446 11398 8498 11450
rect 8510 11398 8562 11450
rect 8574 11398 8626 11450
rect 8638 11398 8690 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 8208 11339 8260 11348
rect 2780 11296 2832 11305
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 1400 11228 1452 11280
rect 8300 11228 8352 11280
rect 2044 11160 2096 11212
rect 6920 11160 6972 11212
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8760 11135 8812 11144
rect 8760 11101 8769 11135
rect 8769 11101 8803 11135
rect 8803 11101 8812 11135
rect 8760 11092 8812 11101
rect 10048 11296 10100 11348
rect 10140 11296 10192 11348
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 11520 11296 11572 11348
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 16948 11296 17000 11348
rect 9036 11160 9088 11212
rect 10692 11160 10744 11212
rect 14004 11228 14056 11280
rect 20720 11296 20772 11348
rect 22468 11296 22520 11348
rect 19064 11271 19116 11280
rect 19064 11237 19098 11271
rect 19098 11237 19116 11271
rect 19064 11228 19116 11237
rect 19340 11228 19392 11280
rect 21364 11271 21416 11280
rect 21364 11237 21373 11271
rect 21373 11237 21407 11271
rect 21407 11237 21416 11271
rect 21364 11228 21416 11237
rect 21640 11228 21692 11280
rect 22652 11228 22704 11280
rect 14096 11160 14148 11212
rect 14280 11160 14332 11212
rect 15108 11160 15160 11212
rect 16396 11160 16448 11212
rect 17960 11160 18012 11212
rect 19892 11160 19944 11212
rect 21456 11160 21508 11212
rect 9772 11092 9824 11144
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 9680 11024 9732 11076
rect 10048 10956 10100 11008
rect 10968 11092 11020 11144
rect 12532 11092 12584 11144
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 15200 11092 15252 11144
rect 21640 11092 21692 11144
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 18328 11024 18380 11076
rect 18696 11067 18748 11076
rect 18696 11033 18705 11067
rect 18705 11033 18739 11067
rect 18739 11033 18748 11067
rect 18696 11024 18748 11033
rect 20260 11024 20312 11076
rect 20536 11024 20588 11076
rect 11060 10956 11112 11008
rect 14372 10999 14424 11008
rect 14372 10965 14381 10999
rect 14381 10965 14415 10999
rect 14415 10965 14424 10999
rect 14372 10956 14424 10965
rect 14648 10956 14700 11008
rect 19432 10956 19484 11008
rect 20168 10999 20220 11008
rect 20168 10965 20177 10999
rect 20177 10965 20211 10999
rect 20211 10965 20220 10999
rect 20168 10956 20220 10965
rect 4714 10854 4766 10906
rect 4778 10854 4830 10906
rect 4842 10854 4894 10906
rect 4906 10854 4958 10906
rect 12178 10854 12230 10906
rect 12242 10854 12294 10906
rect 12306 10854 12358 10906
rect 12370 10854 12422 10906
rect 19642 10854 19694 10906
rect 19706 10854 19758 10906
rect 19770 10854 19822 10906
rect 19834 10854 19886 10906
rect 8300 10752 8352 10804
rect 8668 10795 8720 10804
rect 8668 10761 8677 10795
rect 8677 10761 8711 10795
rect 8711 10761 8720 10795
rect 8668 10752 8720 10761
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 11796 10752 11848 10804
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14464 10752 14516 10804
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 6920 10616 6972 10668
rect 14372 10616 14424 10668
rect 14924 10616 14976 10668
rect 19064 10659 19116 10668
rect 19064 10625 19073 10659
rect 19073 10625 19107 10659
rect 19107 10625 19116 10659
rect 19064 10616 19116 10625
rect 8760 10548 8812 10600
rect 9956 10548 10008 10600
rect 10140 10548 10192 10600
rect 11060 10591 11112 10600
rect 11060 10557 11094 10591
rect 11094 10557 11112 10591
rect 11060 10548 11112 10557
rect 12808 10548 12860 10600
rect 14556 10591 14608 10600
rect 14556 10557 14565 10591
rect 14565 10557 14599 10591
rect 14599 10557 14608 10591
rect 14556 10548 14608 10557
rect 15108 10548 15160 10600
rect 16488 10591 16540 10600
rect 16488 10557 16497 10591
rect 16497 10557 16531 10591
rect 16531 10557 16540 10591
rect 16488 10548 16540 10557
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18972 10591 19024 10600
rect 18972 10557 18981 10591
rect 18981 10557 19015 10591
rect 19015 10557 19024 10591
rect 18972 10548 19024 10557
rect 20076 10752 20128 10804
rect 21364 10752 21416 10804
rect 22376 10752 22428 10804
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19984 10616 20036 10668
rect 19524 10548 19576 10600
rect 20076 10548 20128 10600
rect 20904 10548 20956 10600
rect 21456 10548 21508 10600
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 16212 10480 16264 10532
rect 16396 10480 16448 10532
rect 16948 10480 17000 10532
rect 17040 10480 17092 10532
rect 16856 10412 16908 10464
rect 19340 10480 19392 10532
rect 21640 10523 21692 10532
rect 21640 10489 21674 10523
rect 21674 10489 21692 10523
rect 21640 10480 21692 10489
rect 18604 10412 18656 10464
rect 18696 10412 18748 10464
rect 22836 10455 22888 10464
rect 22836 10421 22845 10455
rect 22845 10421 22879 10455
rect 22879 10421 22888 10455
rect 22836 10412 22888 10421
rect 8446 10310 8498 10362
rect 8510 10310 8562 10362
rect 8574 10310 8626 10362
rect 8638 10310 8690 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9864 10208 9916 10260
rect 9956 10208 10008 10260
rect 10416 10208 10468 10260
rect 11060 10208 11112 10260
rect 8300 10140 8352 10192
rect 10692 10140 10744 10192
rect 14280 10140 14332 10192
rect 9588 10072 9640 10124
rect 14648 10072 14700 10124
rect 15384 10072 15436 10124
rect 15568 10115 15620 10124
rect 15568 10081 15602 10115
rect 15602 10081 15620 10115
rect 15568 10072 15620 10081
rect 16672 10072 16724 10124
rect 20076 10208 20128 10260
rect 21640 10208 21692 10260
rect 22836 10208 22888 10260
rect 18972 10140 19024 10192
rect 19432 10140 19484 10192
rect 10048 10004 10100 10056
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15108 10004 15160 10056
rect 17040 10004 17092 10056
rect 14188 9936 14240 9988
rect 16396 9936 16448 9988
rect 16856 9936 16908 9988
rect 17408 10004 17460 10056
rect 18604 10072 18656 10124
rect 20720 10072 20772 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21180 10115 21232 10124
rect 21180 10081 21214 10115
rect 21214 10081 21232 10115
rect 21180 10072 21232 10081
rect 22468 10072 22520 10124
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 20168 10047 20220 10056
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 20812 10004 20864 10056
rect 22376 10004 22428 10056
rect 12072 9868 12124 9920
rect 20076 9936 20128 9988
rect 20628 9936 20680 9988
rect 18236 9868 18288 9920
rect 21548 9868 21600 9920
rect 23112 9868 23164 9920
rect 4714 9766 4766 9818
rect 4778 9766 4830 9818
rect 4842 9766 4894 9818
rect 4906 9766 4958 9818
rect 12178 9766 12230 9818
rect 12242 9766 12294 9818
rect 12306 9766 12358 9818
rect 12370 9766 12422 9818
rect 19642 9766 19694 9818
rect 19706 9766 19758 9818
rect 19770 9766 19822 9818
rect 19834 9766 19886 9818
rect 17960 9664 18012 9716
rect 18236 9664 18288 9716
rect 21180 9707 21232 9716
rect 21180 9673 21189 9707
rect 21189 9673 21223 9707
rect 21223 9673 21232 9707
rect 21180 9664 21232 9673
rect 9772 9596 9824 9648
rect 11704 9596 11756 9648
rect 15384 9596 15436 9648
rect 12072 9571 12124 9580
rect 12072 9537 12081 9571
rect 12081 9537 12115 9571
rect 12115 9537 12124 9571
rect 12072 9528 12124 9537
rect 18052 9596 18104 9648
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 9680 9460 9732 9512
rect 12992 9460 13044 9512
rect 13820 9460 13872 9512
rect 10876 9392 10928 9444
rect 13176 9392 13228 9444
rect 15476 9392 15528 9444
rect 16856 9460 16908 9512
rect 22652 9596 22704 9648
rect 22928 9639 22980 9648
rect 22928 9605 22937 9639
rect 22937 9605 22971 9639
rect 22971 9605 22980 9639
rect 22928 9596 22980 9605
rect 17960 9460 18012 9512
rect 18328 9503 18380 9512
rect 18328 9469 18362 9503
rect 18362 9469 18380 9503
rect 18328 9460 18380 9469
rect 18604 9460 18656 9512
rect 16948 9392 17000 9444
rect 11612 9324 11664 9376
rect 13544 9324 13596 9376
rect 15384 9324 15436 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16396 9324 16448 9376
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 18420 9392 18472 9444
rect 20812 9460 20864 9512
rect 23020 9528 23072 9580
rect 20168 9392 20220 9444
rect 20720 9392 20772 9444
rect 21548 9392 21600 9444
rect 17592 9324 17644 9333
rect 19340 9324 19392 9376
rect 19432 9324 19484 9376
rect 19800 9324 19852 9376
rect 23020 9367 23072 9376
rect 23020 9333 23029 9367
rect 23029 9333 23063 9367
rect 23063 9333 23072 9367
rect 23020 9324 23072 9333
rect 23664 9528 23716 9580
rect 23664 9392 23716 9444
rect 8446 9222 8498 9274
rect 8510 9222 8562 9274
rect 8574 9222 8626 9274
rect 8638 9222 8690 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 10876 9120 10928 9172
rect 15752 9120 15804 9172
rect 19800 9120 19852 9172
rect 21916 9120 21968 9172
rect 13544 9095 13596 9104
rect 9588 8984 9640 9036
rect 10508 8984 10560 9036
rect 11520 8984 11572 9036
rect 13544 9061 13578 9095
rect 13578 9061 13596 9095
rect 13544 9052 13596 9061
rect 12624 8984 12676 9036
rect 12900 8984 12952 9036
rect 16764 9052 16816 9104
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 15108 8984 15160 9036
rect 15200 8916 15252 8968
rect 16396 8984 16448 9036
rect 17960 9052 18012 9104
rect 19340 9052 19392 9104
rect 23664 9052 23716 9104
rect 17868 8984 17920 9036
rect 18604 8984 18656 9036
rect 19524 8984 19576 9036
rect 20352 9027 20404 9036
rect 20352 8993 20361 9027
rect 20361 8993 20395 9027
rect 20395 8993 20404 9027
rect 20352 8984 20404 8993
rect 20720 8984 20772 9036
rect 22468 8984 22520 9036
rect 16488 8916 16540 8968
rect 18236 8916 18288 8968
rect 19616 8916 19668 8968
rect 14464 8848 14516 8900
rect 19984 8891 20036 8900
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 12992 8780 13044 8832
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 14004 8780 14056 8832
rect 14280 8780 14332 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 18052 8780 18104 8832
rect 19984 8857 19993 8891
rect 19993 8857 20027 8891
rect 20027 8857 20036 8891
rect 19984 8848 20036 8857
rect 21088 8780 21140 8832
rect 22284 8780 22336 8832
rect 4714 8678 4766 8730
rect 4778 8678 4830 8730
rect 4842 8678 4894 8730
rect 4906 8678 4958 8730
rect 12178 8678 12230 8730
rect 12242 8678 12294 8730
rect 12306 8678 12358 8730
rect 12370 8678 12422 8730
rect 19642 8678 19694 8730
rect 19706 8678 19758 8730
rect 19770 8678 19822 8730
rect 19834 8678 19886 8730
rect 2872 8440 2924 8492
rect 9588 8576 9640 8628
rect 10508 8576 10560 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 12624 8576 12676 8628
rect 14648 8576 14700 8628
rect 15568 8576 15620 8628
rect 16672 8576 16724 8628
rect 17592 8576 17644 8628
rect 18696 8576 18748 8628
rect 11980 8440 12032 8492
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 16580 8508 16632 8560
rect 17040 8508 17092 8560
rect 17500 8508 17552 8560
rect 19524 8576 19576 8628
rect 22008 8576 22060 8628
rect 7748 8372 7800 8424
rect 10876 8372 10928 8424
rect 11060 8415 11112 8424
rect 11060 8381 11069 8415
rect 11069 8381 11103 8415
rect 11103 8381 11112 8415
rect 11060 8372 11112 8381
rect 11612 8372 11664 8424
rect 11244 8304 11296 8356
rect 14464 8372 14516 8424
rect 14648 8372 14700 8424
rect 16856 8440 16908 8492
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 17960 8440 18012 8492
rect 19800 8508 19852 8560
rect 22376 8508 22428 8560
rect 18236 8440 18288 8492
rect 19708 8440 19760 8492
rect 20536 8440 20588 8492
rect 13820 8304 13872 8356
rect 15568 8372 15620 8424
rect 16396 8304 16448 8356
rect 22284 8440 22336 8492
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 20996 8372 21048 8424
rect 19800 8304 19852 8356
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 14372 8279 14424 8288
rect 14372 8245 14381 8279
rect 14381 8245 14415 8279
rect 14415 8245 14424 8279
rect 14372 8236 14424 8245
rect 14648 8236 14700 8288
rect 15108 8236 15160 8288
rect 16488 8236 16540 8288
rect 16764 8236 16816 8288
rect 18052 8236 18104 8288
rect 18420 8236 18472 8288
rect 19340 8236 19392 8288
rect 19708 8236 19760 8288
rect 19892 8236 19944 8288
rect 21088 8236 21140 8288
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 21824 8236 21876 8245
rect 22468 8236 22520 8288
rect 8446 8134 8498 8186
rect 8510 8134 8562 8186
rect 8574 8134 8626 8186
rect 8638 8134 8690 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 9588 8032 9640 8084
rect 11980 8032 12032 8084
rect 13176 8032 13228 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 16396 8032 16448 8084
rect 16488 8075 16540 8084
rect 16488 8041 16503 8075
rect 16503 8041 16537 8075
rect 16537 8041 16540 8075
rect 16488 8032 16540 8041
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8208 7896 8260 7948
rect 9588 7896 9640 7948
rect 9772 7896 9824 7948
rect 11060 7964 11112 8016
rect 11796 7964 11848 8016
rect 14924 7964 14976 8016
rect 17592 8032 17644 8084
rect 18144 7964 18196 8016
rect 18512 8032 18564 8084
rect 19156 8032 19208 8084
rect 19340 8032 19392 8084
rect 20352 8032 20404 8084
rect 22560 8075 22612 8084
rect 22560 8041 22569 8075
rect 22569 8041 22603 8075
rect 22603 8041 22612 8075
rect 22560 8032 22612 8041
rect 10876 7896 10928 7948
rect 12624 7896 12676 7948
rect 12992 7896 13044 7948
rect 14096 7896 14148 7948
rect 14464 7896 14516 7948
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 18052 7896 18104 7948
rect 18420 7896 18472 7948
rect 18604 7896 18656 7948
rect 10968 7828 11020 7880
rect 12072 7828 12124 7880
rect 13084 7828 13136 7880
rect 14648 7760 14700 7812
rect 10968 7692 11020 7744
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 14004 7692 14056 7744
rect 14556 7692 14608 7744
rect 15384 7828 15436 7880
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 16488 7871 16540 7880
rect 16488 7837 16500 7871
rect 16500 7837 16534 7871
rect 16534 7837 16540 7871
rect 16488 7828 16540 7837
rect 17408 7828 17460 7880
rect 19984 7896 20036 7948
rect 19340 7828 19392 7880
rect 15292 7760 15344 7812
rect 22468 7964 22520 8016
rect 22928 8007 22980 8016
rect 22928 7973 22937 8007
rect 22937 7973 22971 8007
rect 22971 7973 22980 8007
rect 22928 7964 22980 7973
rect 21456 7939 21508 7948
rect 21456 7905 21490 7939
rect 21490 7905 21508 7939
rect 21456 7896 21508 7905
rect 23020 7896 23072 7948
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 21088 7828 21140 7880
rect 20720 7760 20772 7812
rect 4714 7590 4766 7642
rect 4778 7590 4830 7642
rect 4842 7590 4894 7642
rect 4906 7590 4958 7642
rect 12178 7590 12230 7642
rect 12242 7590 12294 7642
rect 12306 7590 12358 7642
rect 12370 7590 12422 7642
rect 19642 7590 19694 7642
rect 19706 7590 19758 7642
rect 19770 7590 19822 7642
rect 19834 7590 19886 7642
rect 10876 7488 10928 7540
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 14096 7531 14148 7540
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 10968 7284 11020 7336
rect 11152 7327 11204 7336
rect 11152 7293 11161 7327
rect 11161 7293 11195 7327
rect 11195 7293 11204 7327
rect 11152 7284 11204 7293
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 14464 7420 14516 7472
rect 14740 7420 14792 7472
rect 16396 7488 16448 7540
rect 13268 7327 13320 7336
rect 13268 7293 13277 7327
rect 13277 7293 13311 7327
rect 13311 7293 13320 7327
rect 13268 7284 13320 7293
rect 16672 7352 16724 7404
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 14004 7284 14056 7336
rect 15108 7284 15160 7336
rect 16580 7284 16632 7336
rect 16764 7284 16816 7336
rect 11428 7216 11480 7268
rect 11704 7216 11756 7268
rect 12624 7216 12676 7268
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 15476 7216 15528 7268
rect 16488 7216 16540 7268
rect 14004 7148 14056 7200
rect 14464 7148 14516 7200
rect 14740 7148 14792 7200
rect 15292 7148 15344 7200
rect 17960 7488 18012 7540
rect 19616 7463 19668 7472
rect 19616 7429 19625 7463
rect 19625 7429 19659 7463
rect 19659 7429 19668 7463
rect 19616 7420 19668 7429
rect 17868 7327 17920 7336
rect 17868 7293 17877 7327
rect 17877 7293 17911 7327
rect 17911 7293 17920 7327
rect 17868 7284 17920 7293
rect 19984 7352 20036 7404
rect 20720 7488 20772 7540
rect 21456 7488 21508 7540
rect 22284 7352 22336 7404
rect 19432 7284 19484 7336
rect 19616 7284 19668 7336
rect 18144 7216 18196 7268
rect 20536 7284 20588 7336
rect 21088 7284 21140 7336
rect 22836 7284 22888 7336
rect 20720 7259 20772 7268
rect 20720 7225 20754 7259
rect 20754 7225 20772 7259
rect 20720 7216 20772 7225
rect 16672 7148 16724 7200
rect 17592 7148 17644 7200
rect 18052 7148 18104 7200
rect 19340 7148 19392 7200
rect 19984 7191 20036 7200
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 22100 7216 22152 7268
rect 23480 7216 23532 7268
rect 22008 7148 22060 7200
rect 22560 7148 22612 7200
rect 8446 7046 8498 7098
rect 8510 7046 8562 7098
rect 8574 7046 8626 7098
rect 8638 7046 8690 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 8208 6944 8260 6996
rect 10876 6876 10928 6928
rect 9312 6808 9364 6860
rect 11520 6851 11572 6860
rect 11520 6817 11529 6851
rect 11529 6817 11563 6851
rect 11563 6817 11572 6851
rect 11520 6808 11572 6817
rect 12072 6876 12124 6928
rect 12532 6876 12584 6928
rect 12624 6876 12676 6928
rect 13268 6944 13320 6996
rect 14372 6944 14424 6996
rect 14740 6987 14792 6996
rect 14740 6953 14749 6987
rect 14749 6953 14783 6987
rect 14783 6953 14792 6987
rect 14740 6944 14792 6953
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 19156 6944 19208 6996
rect 20904 6944 20956 6996
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 19432 6876 19484 6928
rect 21916 6876 21968 6928
rect 23204 6876 23256 6928
rect 14004 6851 14056 6860
rect 10324 6604 10376 6656
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 15844 6808 15896 6860
rect 16580 6808 16632 6860
rect 17408 6808 17460 6860
rect 19984 6808 20036 6860
rect 20628 6808 20680 6860
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 21088 6808 21140 6860
rect 22008 6808 22060 6860
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 18236 6783 18288 6792
rect 11244 6604 11296 6656
rect 12900 6604 12952 6656
rect 13820 6604 13872 6656
rect 15108 6672 15160 6724
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 20260 6783 20312 6792
rect 19524 6740 19576 6749
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 16488 6672 16540 6724
rect 19248 6672 19300 6724
rect 20536 6740 20588 6792
rect 21824 6740 21876 6792
rect 22192 6740 22244 6792
rect 22100 6672 22152 6724
rect 15568 6604 15620 6656
rect 19156 6604 19208 6656
rect 20444 6604 20496 6656
rect 20996 6604 21048 6656
rect 21272 6604 21324 6656
rect 21916 6647 21968 6656
rect 21916 6613 21925 6647
rect 21925 6613 21959 6647
rect 21959 6613 21968 6647
rect 21916 6604 21968 6613
rect 22192 6604 22244 6656
rect 4714 6502 4766 6554
rect 4778 6502 4830 6554
rect 4842 6502 4894 6554
rect 4906 6502 4958 6554
rect 12178 6502 12230 6554
rect 12242 6502 12294 6554
rect 12306 6502 12358 6554
rect 12370 6502 12422 6554
rect 19642 6502 19694 6554
rect 19706 6502 19758 6554
rect 19770 6502 19822 6554
rect 19834 6502 19886 6554
rect 9312 6400 9364 6452
rect 11060 6400 11112 6452
rect 11520 6400 11572 6452
rect 12532 6400 12584 6452
rect 12992 6400 13044 6452
rect 15476 6400 15528 6452
rect 15844 6400 15896 6452
rect 17592 6307 17644 6316
rect 10324 6196 10376 6248
rect 11336 6128 11388 6180
rect 13820 6196 13872 6248
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 18144 6264 18196 6316
rect 18236 6196 18288 6248
rect 19432 6332 19484 6384
rect 20720 6332 20772 6384
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 20536 6264 20588 6316
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 19432 6196 19484 6248
rect 19531 6239 19583 6248
rect 19531 6205 19540 6239
rect 19540 6205 19574 6239
rect 19574 6205 19583 6239
rect 19800 6239 19852 6248
rect 19531 6196 19583 6205
rect 19800 6205 19834 6239
rect 19834 6205 19852 6239
rect 19800 6196 19852 6205
rect 20352 6196 20404 6248
rect 20904 6196 20956 6248
rect 21824 6239 21876 6248
rect 21824 6205 21833 6239
rect 21833 6205 21867 6239
rect 21867 6205 21876 6239
rect 21824 6196 21876 6205
rect 22284 6196 22336 6248
rect 14004 6128 14056 6180
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 12900 6060 12952 6112
rect 14740 6128 14792 6180
rect 20720 6128 20772 6180
rect 21640 6128 21692 6180
rect 22928 6171 22980 6180
rect 22928 6137 22937 6171
rect 22937 6137 22971 6171
rect 22971 6137 22980 6171
rect 22928 6128 22980 6137
rect 19340 6060 19392 6112
rect 20996 6103 21048 6112
rect 20996 6069 21005 6103
rect 21005 6069 21039 6103
rect 21039 6069 21048 6103
rect 22008 6103 22060 6112
rect 20996 6060 21048 6069
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 8446 5958 8498 6010
rect 8510 5958 8562 6010
rect 8574 5958 8626 6010
rect 8638 5958 8690 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 11336 5899 11388 5908
rect 11336 5865 11345 5899
rect 11345 5865 11379 5899
rect 11379 5865 11388 5899
rect 11336 5856 11388 5865
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 14004 5856 14056 5908
rect 11060 5788 11112 5840
rect 11796 5788 11848 5840
rect 12716 5788 12768 5840
rect 13728 5788 13780 5840
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14740 5899 14792 5908
rect 14372 5856 14424 5865
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 15568 5788 15620 5840
rect 9312 5720 9364 5772
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 12992 5720 13044 5772
rect 16488 5720 16540 5772
rect 17224 5720 17276 5772
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 19524 5856 19576 5908
rect 20352 5899 20404 5908
rect 20352 5865 20361 5899
rect 20361 5865 20395 5899
rect 20395 5865 20404 5899
rect 20352 5856 20404 5865
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 20904 5899 20956 5908
rect 20904 5865 20913 5899
rect 20913 5865 20947 5899
rect 20947 5865 20956 5899
rect 20904 5856 20956 5865
rect 21272 5899 21324 5908
rect 21272 5865 21281 5899
rect 21281 5865 21315 5899
rect 21315 5865 21324 5899
rect 21272 5856 21324 5865
rect 21456 5856 21508 5908
rect 22560 5856 22612 5908
rect 22100 5788 22152 5840
rect 19524 5720 19576 5772
rect 20628 5720 20680 5772
rect 22928 5720 22980 5772
rect 16396 5695 16448 5704
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 20536 5652 20588 5704
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 17868 5516 17920 5525
rect 19248 5516 19300 5568
rect 21364 5516 21416 5568
rect 4714 5414 4766 5466
rect 4778 5414 4830 5466
rect 4842 5414 4894 5466
rect 4906 5414 4958 5466
rect 12178 5414 12230 5466
rect 12242 5414 12294 5466
rect 12306 5414 12358 5466
rect 12370 5414 12422 5466
rect 19642 5414 19694 5466
rect 19706 5414 19758 5466
rect 19770 5414 19822 5466
rect 19834 5414 19886 5466
rect 13728 5312 13780 5364
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 17224 5312 17276 5364
rect 11336 5176 11388 5228
rect 18328 5312 18380 5364
rect 19432 5312 19484 5364
rect 19340 5176 19392 5228
rect 20352 5244 20404 5296
rect 21088 5312 21140 5364
rect 21456 5244 21508 5296
rect 11796 5040 11848 5092
rect 11152 4972 11204 5024
rect 12992 5108 13044 5160
rect 14280 5108 14332 5160
rect 17868 5108 17920 5160
rect 12808 5040 12860 5092
rect 16304 5040 16356 5092
rect 16396 5040 16448 5092
rect 12900 4972 12952 5024
rect 19524 5040 19576 5092
rect 17868 4972 17920 5024
rect 19248 4972 19300 5024
rect 22192 5312 22244 5364
rect 22284 5312 22336 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 21364 5108 21416 5160
rect 22284 5108 22336 5160
rect 22652 5040 22704 5092
rect 22928 5040 22980 5092
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 22376 4972 22428 5024
rect 8446 4870 8498 4922
rect 8510 4870 8562 4922
rect 8574 4870 8626 4922
rect 8638 4870 8690 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 18236 4768 18288 4820
rect 20168 4768 20220 4820
rect 20260 4768 20312 4820
rect 21640 4768 21692 4820
rect 22928 4811 22980 4820
rect 22928 4777 22937 4811
rect 22937 4777 22971 4811
rect 22971 4777 22980 4811
rect 22928 4768 22980 4777
rect 11152 4743 11204 4752
rect 11152 4709 11161 4743
rect 11161 4709 11195 4743
rect 11195 4709 11204 4743
rect 11152 4700 11204 4709
rect 17776 4700 17828 4752
rect 16488 4632 16540 4684
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11980 4496 12032 4548
rect 19340 4700 19392 4752
rect 19432 4632 19484 4684
rect 20168 4632 20220 4684
rect 20996 4700 21048 4752
rect 22744 4700 22796 4752
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19984 4607 20036 4616
rect 19248 4564 19300 4573
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 20260 4564 20312 4616
rect 21364 4632 21416 4684
rect 22836 4632 22888 4684
rect 17776 4471 17828 4480
rect 17776 4437 17785 4471
rect 17785 4437 17819 4471
rect 17819 4437 17828 4471
rect 17776 4428 17828 4437
rect 19524 4428 19576 4480
rect 4714 4326 4766 4378
rect 4778 4326 4830 4378
rect 4842 4326 4894 4378
rect 4906 4326 4958 4378
rect 12178 4326 12230 4378
rect 12242 4326 12294 4378
rect 12306 4326 12358 4378
rect 12370 4326 12422 4378
rect 19642 4326 19694 4378
rect 19706 4326 19758 4378
rect 19770 4326 19822 4378
rect 19834 4326 19886 4378
rect 19984 4224 20036 4276
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 20904 4088 20956 4140
rect 21364 4088 21416 4140
rect 23020 4131 23072 4140
rect 23020 4097 23029 4131
rect 23029 4097 23063 4131
rect 23063 4097 23072 4131
rect 23020 4088 23072 4097
rect 17776 4020 17828 4072
rect 16488 3952 16540 4004
rect 19524 3952 19576 4004
rect 19800 3952 19852 4004
rect 19984 4063 20036 4072
rect 19984 4029 20018 4063
rect 20018 4029 20036 4063
rect 19984 4020 20036 4029
rect 20904 3952 20956 4004
rect 22744 3952 22796 4004
rect 17960 3884 18012 3936
rect 18236 3884 18288 3936
rect 20168 3884 20220 3936
rect 8446 3782 8498 3834
rect 8510 3782 8562 3834
rect 8574 3782 8626 3834
rect 8638 3782 8690 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 18052 3680 18104 3732
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 19800 3723 19852 3732
rect 19800 3689 19809 3723
rect 19809 3689 19843 3723
rect 19843 3689 19852 3723
rect 19800 3680 19852 3689
rect 20260 3680 20312 3732
rect 20536 3680 20588 3732
rect 22192 3680 22244 3732
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 3148 3612 3200 3621
rect 17960 3612 18012 3664
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 17868 3544 17920 3596
rect 16488 3519 16540 3528
rect 16488 3485 16497 3519
rect 16497 3485 16531 3519
rect 16531 3485 16540 3519
rect 16488 3476 16540 3485
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 22008 3612 22060 3664
rect 20352 3544 20404 3596
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 20996 3544 21048 3596
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 22928 3519 22980 3528
rect 22928 3485 22937 3519
rect 22937 3485 22971 3519
rect 22971 3485 22980 3519
rect 22928 3476 22980 3485
rect 19340 3451 19392 3460
rect 19340 3417 19349 3451
rect 19349 3417 19383 3451
rect 19383 3417 19392 3451
rect 19340 3408 19392 3417
rect 22376 3451 22428 3460
rect 22376 3417 22385 3451
rect 22385 3417 22419 3451
rect 22419 3417 22428 3451
rect 22376 3408 22428 3417
rect 17776 3340 17828 3392
rect 22008 3340 22060 3392
rect 22192 3340 22244 3392
rect 4714 3238 4766 3290
rect 4778 3238 4830 3290
rect 4842 3238 4894 3290
rect 4906 3238 4958 3290
rect 12178 3238 12230 3290
rect 12242 3238 12294 3290
rect 12306 3238 12358 3290
rect 12370 3238 12422 3290
rect 19642 3238 19694 3290
rect 19706 3238 19758 3290
rect 19770 3238 19822 3290
rect 19834 3238 19886 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 2504 3136 2556 3188
rect 10232 3136 10284 3188
rect 17868 3179 17920 3188
rect 2044 3068 2096 3120
rect 17868 3145 17877 3179
rect 17877 3145 17911 3179
rect 17911 3145 17920 3179
rect 17868 3136 17920 3145
rect 19156 3136 19208 3188
rect 20996 3136 21048 3188
rect 22284 3179 22336 3188
rect 22284 3145 22293 3179
rect 22293 3145 22327 3179
rect 22327 3145 22336 3179
rect 22284 3136 22336 3145
rect 18880 3068 18932 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 22928 3043 22980 3052
rect 2504 2975 2556 2984
rect 2504 2941 2535 2975
rect 2535 2941 2556 2975
rect 2504 2932 2556 2941
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 16488 2975 16540 2984
rect 16488 2941 16497 2975
rect 16497 2941 16531 2975
rect 16531 2941 16540 2975
rect 16488 2932 16540 2941
rect 17868 2932 17920 2984
rect 17776 2864 17828 2916
rect 18052 2796 18104 2848
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 20168 2932 20220 2984
rect 20260 2864 20312 2916
rect 20904 2932 20956 2984
rect 22652 2975 22704 2984
rect 22652 2941 22661 2975
rect 22661 2941 22695 2975
rect 22695 2941 22704 2975
rect 22652 2932 22704 2941
rect 22836 2932 22888 2984
rect 20720 2839 20772 2848
rect 20720 2805 20729 2839
rect 20729 2805 20763 2839
rect 20763 2805 20772 2839
rect 20720 2796 20772 2805
rect 22652 2796 22704 2848
rect 23020 2796 23072 2848
rect 8446 2694 8498 2746
rect 8510 2694 8562 2746
rect 8574 2694 8626 2746
rect 8638 2694 8690 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 19524 2592 19576 2644
rect 20076 2592 20128 2644
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 22744 2592 22796 2644
rect 19340 2524 19392 2576
rect 20996 2524 21048 2576
rect 22008 2524 22060 2576
rect 18052 2456 18104 2508
rect 20904 2456 20956 2508
rect 22652 2499 22704 2508
rect 22652 2465 22661 2499
rect 22661 2465 22695 2499
rect 22695 2465 22704 2499
rect 22652 2456 22704 2465
rect 20260 2388 20312 2440
rect 22468 2388 22520 2440
rect 4714 2150 4766 2202
rect 4778 2150 4830 2202
rect 4842 2150 4894 2202
rect 4906 2150 4958 2202
rect 12178 2150 12230 2202
rect 12242 2150 12294 2202
rect 12306 2150 12358 2202
rect 12370 2150 12422 2202
rect 19642 2150 19694 2202
rect 19706 2150 19758 2202
rect 19770 2150 19822 2202
rect 19834 2150 19886 2202
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 15106 23800 15162 24600
rect 15750 23800 15806 24600
rect 16394 23800 16450 24600
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21546 23800 21602 24600
rect 21822 24304 21878 24313
rect 21822 24239 21878 24248
rect 308 21690 336 23800
rect 296 21684 348 21690
rect 296 21626 348 21632
rect 952 21622 980 23800
rect 940 21616 992 21622
rect 940 21558 992 21564
rect 1596 21146 1624 23800
rect 2240 21146 2268 23800
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2332 21593 2360 21830
rect 2318 21584 2374 21593
rect 2318 21519 2320 21528
rect 2372 21519 2374 21528
rect 2320 21490 2372 21496
rect 2332 21459 2360 21490
rect 2424 21486 2452 21966
rect 2884 21690 2912 23800
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 2608 21078 2636 21422
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2976 20602 3004 20946
rect 3528 20602 3556 23800
rect 4172 21962 4200 23800
rect 4816 22930 4844 23800
rect 4816 22902 5212 22930
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21418 4568 21830
rect 4688 21788 4984 21808
rect 4744 21786 4768 21788
rect 4824 21786 4848 21788
rect 4904 21786 4928 21788
rect 4766 21734 4768 21786
rect 4830 21734 4842 21786
rect 4904 21734 4906 21786
rect 4744 21732 4768 21734
rect 4824 21732 4848 21734
rect 4904 21732 4928 21734
rect 4688 21712 4984 21732
rect 5184 21690 5212 22902
rect 5460 22438 5488 23800
rect 6104 22930 6132 23800
rect 6104 22902 6408 22930
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5264 22092 5316 22098
rect 5264 22034 5316 22040
rect 5276 21962 5304 22034
rect 5264 21956 5316 21962
rect 5264 21898 5316 21904
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 4344 21412 4396 21418
rect 4344 21354 4396 21360
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 4172 21078 4200 21286
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 1582 20496 1638 20505
rect 1582 20431 1584 20440
rect 1636 20431 1638 20440
rect 1584 20402 1636 20408
rect 1596 19922 1624 20402
rect 2976 20398 3004 20538
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 2976 20058 3004 20198
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3068 19990 3096 20198
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 3056 19984 3108 19990
rect 3056 19926 3108 19932
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 1596 18834 1624 19858
rect 2792 19174 2820 19858
rect 2884 19174 2912 19926
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3068 19310 3096 19654
rect 3160 19378 3188 20402
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 2884 18970 2912 19110
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 3068 18834 3096 19110
rect 3436 18902 3464 19110
rect 3528 18970 3556 19790
rect 3620 19446 3648 19858
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 3516 18828 3568 18834
rect 3516 18770 3568 18776
rect 1596 17202 1624 18770
rect 3068 18426 3096 18770
rect 3528 18426 3556 18770
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 17814 1808 18158
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1596 16658 1624 17138
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 3068 16794 3096 17002
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 1584 16652 1636 16658
rect 1636 16612 1716 16640
rect 1584 16594 1636 16600
rect 1688 16046 1716 16612
rect 2700 16561 2728 16662
rect 3160 16658 3188 17614
rect 3252 17202 3280 17750
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 3344 16250 3372 17682
rect 3620 17678 3648 19110
rect 3712 18766 3740 20402
rect 3804 19786 3832 20742
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 20058 3924 20198
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3988 19938 4016 20878
rect 4172 20398 4200 21014
rect 4356 20806 4384 21354
rect 4540 21078 4568 21354
rect 4528 21072 4580 21078
rect 4528 21014 4580 21020
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4356 20466 4384 20742
rect 4632 20505 4660 21422
rect 5092 21146 5120 21422
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5184 20806 5212 20946
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 4688 20700 4984 20720
rect 4744 20698 4768 20700
rect 4824 20698 4848 20700
rect 4904 20698 4928 20700
rect 4766 20646 4768 20698
rect 4830 20646 4842 20698
rect 4904 20646 4906 20698
rect 4744 20644 4768 20646
rect 4824 20644 4848 20646
rect 4904 20644 4928 20646
rect 4688 20624 4984 20644
rect 4618 20496 4674 20505
rect 4344 20460 4396 20466
rect 4618 20431 4674 20440
rect 4986 20496 5042 20505
rect 5184 20466 5212 20742
rect 4986 20431 5042 20440
rect 5172 20460 5224 20466
rect 4344 20402 4396 20408
rect 5000 20398 5028 20431
rect 5172 20402 5224 20408
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 3896 19910 4016 19938
rect 5264 19916 5316 19922
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17134 3648 17478
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 3424 16992 3476 16998
rect 3476 16940 3556 16946
rect 3424 16934 3556 16940
rect 3436 16918 3556 16934
rect 3528 16658 3556 16918
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3528 16046 3556 16594
rect 3620 16046 3648 17070
rect 3712 16590 3740 18702
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3712 16182 3740 16526
rect 3804 16250 3832 19382
rect 3896 18222 3924 19910
rect 5264 19858 5316 19864
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3988 19378 4016 19790
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 4080 19242 4108 19654
rect 4688 19612 4984 19632
rect 4744 19610 4768 19612
rect 4824 19610 4848 19612
rect 4904 19610 4928 19612
rect 4766 19558 4768 19610
rect 4830 19558 4842 19610
rect 4904 19558 4906 19610
rect 4744 19556 4768 19558
rect 4824 19556 4848 19558
rect 4904 19556 4928 19558
rect 4688 19536 4984 19556
rect 5276 19514 5304 19858
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 5368 19174 5396 22102
rect 5552 22098 5580 22442
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5460 21146 5488 21354
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5552 19922 5580 21830
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5644 19854 5672 20266
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 4632 18970 4660 19110
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 17814 3924 18158
rect 4264 18154 4292 18634
rect 4688 18524 4984 18544
rect 4744 18522 4768 18524
rect 4824 18522 4848 18524
rect 4904 18522 4928 18524
rect 4766 18470 4768 18522
rect 4830 18470 4842 18522
rect 4904 18470 4906 18522
rect 4744 18468 4768 18470
rect 4824 18468 4848 18470
rect 4904 18468 4928 18470
rect 4688 18448 4984 18468
rect 5184 18426 5212 19110
rect 5552 18766 5580 19722
rect 5644 19378 5672 19790
rect 5736 19786 5764 21830
rect 5828 21146 5856 21898
rect 5920 21554 5948 21966
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5828 19786 5856 20878
rect 5920 20398 5948 21286
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 6012 20505 6040 21082
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 20806 6224 20878
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 5998 20496 6054 20505
rect 5998 20431 6054 20440
rect 6196 20398 6224 20742
rect 6288 20466 6316 22034
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5920 19378 5948 20334
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6104 18834 6132 19926
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 19310 6224 19790
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6196 19174 6224 19246
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 3884 17808 3936 17814
rect 3884 17750 3936 17756
rect 4264 17338 4292 18090
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4632 17202 4660 17750
rect 4688 17436 4984 17456
rect 4744 17434 4768 17436
rect 4824 17434 4848 17436
rect 4904 17434 4928 17436
rect 4766 17382 4768 17434
rect 4830 17382 4842 17434
rect 4904 17382 4906 17434
rect 4744 17380 4768 17382
rect 4824 17380 4848 17382
rect 4904 17380 4928 17382
rect 4688 17360 4984 17380
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 5644 17134 5672 18770
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5736 17814 5764 18702
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 18222 6224 18566
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6196 17814 6224 18022
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 17134 6224 17478
rect 6288 17338 6316 18022
rect 6380 17338 6408 22902
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 21078 6500 21966
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6656 21298 6684 22374
rect 6748 21690 6776 23800
rect 7392 22930 7420 23800
rect 7392 22902 7512 22930
rect 6920 22500 6972 22506
rect 6920 22442 6972 22448
rect 6932 22166 6960 22442
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 7196 21888 7248 21894
rect 7248 21836 7328 21842
rect 7196 21830 7328 21836
rect 7208 21814 7328 21830
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6748 21486 6776 21626
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 7300 21350 7328 21814
rect 6920 21344 6972 21350
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6472 20602 6500 21014
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 1688 15570 1716 15982
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 2056 14958 2084 15982
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2870 15328 2926 15337
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1780 14482 1808 14894
rect 2792 14550 2820 15302
rect 2870 15263 2926 15272
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1780 14074 1808 14418
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 2686 13832 2742 13841
rect 2792 13802 2820 14486
rect 2686 13767 2688 13776
rect 2740 13767 2742 13776
rect 2780 13796 2832 13802
rect 2688 13738 2740 13744
rect 2780 13738 2832 13744
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12238 2084 12718
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11762 2084 12174
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1412 10470 1440 11222
rect 2056 11218 2084 11698
rect 2792 11354 2820 12310
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 9217 1440 10406
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 2884 8498 2912 15263
rect 2976 14074 3004 15438
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3068 14006 3096 15506
rect 3148 14884 3200 14890
rect 3148 14826 3200 14832
rect 3160 14618 3188 14826
rect 3436 14618 3464 15506
rect 4080 15502 4108 16730
rect 4724 16658 4752 16730
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4688 16348 4984 16368
rect 4744 16346 4768 16348
rect 4824 16346 4848 16348
rect 4904 16346 4928 16348
rect 4766 16294 4768 16346
rect 4830 16294 4842 16346
rect 4904 16294 4906 16346
rect 4744 16292 4768 16294
rect 4824 16292 4848 16294
rect 4904 16292 4928 16294
rect 4688 16272 4984 16292
rect 4620 16108 4672 16114
rect 4540 16068 4620 16096
rect 4540 15638 4568 16068
rect 4620 16050 4672 16056
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3528 14482 3556 15302
rect 4080 14958 4108 15438
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4448 14618 4476 14826
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 4540 13938 4568 15574
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4632 15094 4660 15506
rect 4688 15260 4984 15280
rect 4744 15258 4768 15260
rect 4824 15258 4848 15260
rect 4904 15258 4928 15260
rect 4766 15206 4768 15258
rect 4830 15206 4842 15258
rect 4904 15206 4906 15258
rect 4744 15204 4768 15206
rect 4824 15204 4848 15206
rect 4904 15204 4928 15206
rect 4688 15184 4984 15204
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4632 14550 4660 15030
rect 5092 14618 5120 15982
rect 5276 15570 5304 17002
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6196 16726 6224 16934
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6182 16552 6238 16561
rect 6288 16538 6316 16934
rect 6380 16658 6408 17274
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6472 16794 6500 17070
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6238 16510 6316 16538
rect 6182 16487 6184 16496
rect 6236 16487 6238 16496
rect 6184 16458 6236 16464
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5828 16114 5856 16390
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5276 14958 5304 15302
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4688 14172 4984 14192
rect 4744 14170 4768 14172
rect 4824 14170 4848 14172
rect 4904 14170 4928 14172
rect 4766 14118 4768 14170
rect 4830 14118 4842 14170
rect 4904 14118 4906 14170
rect 4744 14116 4768 14118
rect 4824 14116 4848 14118
rect 4904 14116 4928 14118
rect 4688 14096 4984 14116
rect 5184 14074 5212 14826
rect 5276 14618 5304 14894
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5368 14346 5396 15982
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5736 14618 5764 15914
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6380 15162 6408 15506
rect 6472 15162 6500 16730
rect 6564 16114 6592 21286
rect 6656 21270 6776 21298
rect 6920 21286 6972 21292
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6656 20602 6684 21082
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6748 20482 6776 21270
rect 6932 20534 6960 21286
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 6656 20454 6776 20482
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6656 16794 6684 20454
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6748 19854 6776 20334
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6748 19514 6776 19654
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6748 18970 6776 19450
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 17338 6868 18838
rect 6932 17762 6960 20470
rect 7208 20398 7236 20878
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7024 19990 7052 20198
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 7024 19378 7052 19926
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7116 18766 7144 19654
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 18222 7144 18702
rect 7208 18698 7236 19110
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6932 17734 7052 17762
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6656 16046 6684 16730
rect 6932 16590 6960 17614
rect 7024 17202 7052 17734
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6932 16130 6960 16526
rect 6840 16102 7052 16130
rect 6840 16046 6868 16102
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6380 14618 6408 15098
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6564 14414 6592 15846
rect 6932 15366 6960 15914
rect 7024 15502 7052 16102
rect 7208 15910 7236 16594
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15638 7236 15846
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 14550 6960 15302
rect 7392 15026 7420 15982
rect 7484 15706 7512 22902
rect 8036 22234 8064 23800
rect 8680 22506 8708 23800
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 8420 22332 8716 22352
rect 8476 22330 8500 22332
rect 8556 22330 8580 22332
rect 8636 22330 8660 22332
rect 8498 22278 8500 22330
rect 8562 22278 8574 22330
rect 8636 22278 8638 22330
rect 8476 22276 8500 22278
rect 8556 22276 8580 22278
rect 8636 22276 8660 22278
rect 8420 22256 8716 22276
rect 7564 22228 7616 22234
rect 7564 22170 7616 22176
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 7576 21690 7604 22170
rect 7840 22024 7892 22030
rect 7892 21984 7972 22012
rect 7840 21966 7892 21972
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7668 21690 7696 21830
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7852 21554 7880 21830
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18154 7604 18702
rect 7668 18630 7696 19246
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7760 17882 7788 21286
rect 7944 20398 7972 21984
rect 8036 21486 8064 22170
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8298 21584 8354 21593
rect 8116 21548 8168 21554
rect 8404 21554 8432 22102
rect 8298 21519 8354 21528
rect 8392 21548 8444 21554
rect 8116 21490 8168 21496
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8128 21078 8156 21490
rect 8312 21350 8340 21519
rect 8392 21490 8444 21496
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7852 19378 7880 19722
rect 8022 19408 8078 19417
rect 7840 19372 7892 19378
rect 8022 19343 8024 19352
rect 7840 19314 7892 19320
rect 8076 19343 8078 19352
rect 8024 19314 8076 19320
rect 8220 19310 8248 21286
rect 8420 21244 8716 21264
rect 8476 21242 8500 21244
rect 8556 21242 8580 21244
rect 8636 21242 8660 21244
rect 8498 21190 8500 21242
rect 8562 21190 8574 21242
rect 8636 21190 8638 21242
rect 8476 21188 8500 21190
rect 8556 21188 8580 21190
rect 8636 21188 8660 21190
rect 8420 21168 8716 21188
rect 9048 21078 9076 21422
rect 9036 21072 9088 21078
rect 9036 21014 9088 21020
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 20398 8432 20742
rect 9232 20466 9260 21014
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 9324 20330 9352 23800
rect 9968 22250 9996 23800
rect 10612 22250 10640 23800
rect 9876 22222 9996 22250
rect 10336 22222 10640 22250
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8420 20156 8716 20176
rect 8476 20154 8500 20156
rect 8556 20154 8580 20156
rect 8636 20154 8660 20156
rect 8498 20102 8500 20154
rect 8562 20102 8574 20154
rect 8636 20102 8638 20154
rect 8476 20100 8500 20102
rect 8556 20100 8580 20102
rect 8636 20100 8660 20102
rect 8420 20080 8716 20100
rect 8864 20058 8892 20198
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8220 18970 8248 19246
rect 8420 19068 8716 19088
rect 8476 19066 8500 19068
rect 8556 19066 8580 19068
rect 8636 19066 8660 19068
rect 8498 19014 8500 19066
rect 8562 19014 8574 19066
rect 8636 19014 8638 19066
rect 8476 19012 8500 19014
rect 8556 19012 8580 19014
rect 8636 19012 8660 19014
rect 8420 18992 8716 19012
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8036 18290 8064 18770
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8772 18222 8800 18634
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8024 18148 8076 18154
rect 8024 18090 8076 18096
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 8036 17338 8064 18090
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8220 17678 8248 18022
rect 8420 17980 8716 18000
rect 8476 17978 8500 17980
rect 8556 17978 8580 17980
rect 8636 17978 8660 17980
rect 8498 17926 8500 17978
rect 8562 17926 8574 17978
rect 8636 17926 8638 17978
rect 8476 17924 8500 17926
rect 8556 17924 8580 17926
rect 8636 17924 8660 17926
rect 8420 17904 8716 17924
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7484 14822 7512 15642
rect 7668 15162 7696 17070
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 8036 14958 8064 16186
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 6564 13938 6592 14350
rect 7024 14074 7052 14758
rect 8128 14550 8156 17478
rect 8588 17338 8616 17750
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8220 15026 8248 16730
rect 8312 16538 8340 17002
rect 8420 16892 8716 16912
rect 8476 16890 8500 16892
rect 8556 16890 8580 16892
rect 8636 16890 8660 16892
rect 8498 16838 8500 16890
rect 8562 16838 8574 16890
rect 8636 16838 8638 16890
rect 8476 16836 8500 16838
rect 8556 16836 8580 16838
rect 8636 16836 8660 16838
rect 8420 16816 8716 16836
rect 8312 16510 8432 16538
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16114 8340 16390
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8312 15638 8340 16050
rect 8404 15978 8432 16510
rect 8772 16130 8800 18158
rect 8864 16726 8892 19858
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9140 19417 9168 19722
rect 9126 19408 9182 19417
rect 9126 19343 9182 19352
rect 9140 18902 9168 19343
rect 9128 18896 9180 18902
rect 9128 18838 9180 18844
rect 9140 18086 9168 18838
rect 9232 18834 9260 19790
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9324 18290 9352 19858
rect 9692 19854 9720 20266
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9784 19786 9812 20946
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18902 9720 19110
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9036 17808 9088 17814
rect 8956 17768 9036 17796
rect 8956 17610 8984 17768
rect 9036 17750 9088 17756
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8956 16590 8984 17002
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8864 16250 8892 16526
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8772 16102 8892 16130
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8420 15804 8716 15824
rect 8476 15802 8500 15804
rect 8556 15802 8580 15804
rect 8636 15802 8660 15804
rect 8498 15750 8500 15802
rect 8562 15750 8574 15802
rect 8636 15750 8638 15802
rect 8476 15748 8500 15750
rect 8556 15748 8580 15750
rect 8636 15748 8660 15750
rect 8420 15728 8716 15748
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8772 15162 8800 15982
rect 8864 15978 8892 16102
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8956 15434 8984 16526
rect 9048 15706 9076 16594
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 9140 15162 9168 17682
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9232 15570 9260 16594
rect 9324 16250 9352 18226
rect 9416 17542 9444 18566
rect 9508 18086 9536 18770
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9416 15570 9444 17478
rect 9508 17338 9536 18022
rect 9600 17882 9628 18702
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9692 15706 9720 17682
rect 9784 17338 9812 19722
rect 9876 19718 9904 22222
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10048 21480 10100 21486
rect 10046 21448 10048 21457
rect 10100 21448 10102 21457
rect 10046 21383 10102 21392
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 20262 10088 21286
rect 10152 21146 10180 22034
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10244 20058 10272 21966
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9876 17134 9904 19178
rect 9968 18970 9996 19790
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9968 18222 9996 18906
rect 10048 18760 10100 18766
rect 10100 18720 10180 18748
rect 10048 18702 10100 18708
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 10060 17882 10088 18226
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9784 16590 9812 17070
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9784 15434 9812 16526
rect 9876 16114 9904 16934
rect 10060 16114 10088 17478
rect 10152 17066 10180 18720
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10336 17082 10364 22222
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10428 20398 10456 21286
rect 10520 21010 10548 21422
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10612 20398 10640 22102
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10704 20754 10732 21354
rect 11072 21350 11100 21966
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11072 21146 11100 21286
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 10704 20726 10916 20754
rect 10704 20602 10732 20726
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10600 20392 10652 20398
rect 10796 20380 10824 20538
rect 10888 20466 10916 20726
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10600 20334 10652 20340
rect 10704 20352 10824 20380
rect 10704 19514 10732 20352
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10796 19514 10824 20198
rect 11164 19854 11192 21286
rect 11256 19854 11284 23800
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11610 21040 11666 21049
rect 11808 21010 11836 21626
rect 11900 21146 11928 23800
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11992 21570 12020 21966
rect 12152 21788 12448 21808
rect 12208 21786 12232 21788
rect 12288 21786 12312 21788
rect 12368 21786 12392 21788
rect 12230 21734 12232 21786
rect 12294 21734 12306 21786
rect 12368 21734 12370 21786
rect 12208 21732 12232 21734
rect 12288 21732 12312 21734
rect 12368 21732 12392 21734
rect 12152 21712 12448 21732
rect 12072 21616 12124 21622
rect 11992 21564 12072 21570
rect 11992 21558 12124 21564
rect 12544 21570 12572 23800
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12636 21690 12664 22034
rect 12900 21956 12952 21962
rect 12900 21898 12952 21904
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12912 21593 12940 21898
rect 12898 21584 12954 21593
rect 11992 21542 12112 21558
rect 12544 21542 12756 21570
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11610 20975 11666 20984
rect 11796 21004 11848 21010
rect 11624 20874 11652 20975
rect 11796 20946 11848 20952
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 11164 19310 11192 19790
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10796 18426 10824 18702
rect 10980 18426 11008 19178
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10704 17134 10732 18294
rect 11164 18222 11192 19110
rect 11256 18290 11284 19654
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10980 17338 11008 17614
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10692 17128 10744 17134
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 10244 16114 10272 17070
rect 10336 17054 10456 17082
rect 10692 17070 10744 17076
rect 11072 17066 11100 17614
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10336 15910 10364 16934
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15706 10364 15846
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10428 15586 10456 17054
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16794 11100 17002
rect 11256 16794 11284 17070
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10336 15558 10456 15586
rect 11072 15570 11100 15982
rect 11060 15564 11112 15570
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 8420 14716 8716 14736
rect 8476 14714 8500 14716
rect 8556 14714 8580 14716
rect 8636 14714 8660 14716
rect 8498 14662 8500 14714
rect 8562 14662 8574 14714
rect 8636 14662 8638 14714
rect 8476 14660 8500 14662
rect 8556 14660 8580 14662
rect 8636 14660 8660 14662
rect 8420 14640 8716 14660
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3528 13530 3556 13738
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12374 3372 13262
rect 3436 12714 3464 13398
rect 3620 13258 3648 13874
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13530 4108 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3988 12986 4016 13262
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12442 3464 12650
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3160 3670 3188 12038
rect 3988 11694 4016 12922
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4080 12646 4108 12854
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12306 4108 12582
rect 4448 12374 4476 13330
rect 4540 13190 4568 13874
rect 5552 13818 5580 13874
rect 5460 13790 5580 13818
rect 6274 13832 6330 13841
rect 6092 13796 6144 13802
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4688 13084 4984 13104
rect 4744 13082 4768 13084
rect 4824 13082 4848 13084
rect 4904 13082 4928 13084
rect 4766 13030 4768 13082
rect 4830 13030 4842 13082
rect 4904 13030 4906 13082
rect 4744 13028 4768 13030
rect 4824 13028 4848 13030
rect 4904 13028 4928 13030
rect 4688 13008 4984 13028
rect 5092 12986 5120 13330
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5276 12782 5304 13670
rect 5460 13462 5488 13790
rect 6274 13767 6276 13776
rect 6092 13738 6144 13744
rect 6328 13767 6330 13776
rect 6276 13738 6328 13744
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 6104 13394 6132 13738
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13394 6224 13670
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6104 12986 6132 13330
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5276 12442 5304 12718
rect 6288 12442 6316 13738
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13190 6408 13670
rect 6748 13462 6776 13942
rect 7392 13870 7420 14418
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13870 8708 14214
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 6840 13530 6868 13806
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 7392 13326 7420 13806
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8420 13628 8716 13648
rect 8476 13626 8500 13628
rect 8556 13626 8580 13628
rect 8636 13626 8660 13628
rect 8498 13574 8500 13626
rect 8562 13574 8574 13626
rect 8636 13574 8638 13626
rect 8476 13572 8500 13574
rect 8556 13572 8580 13574
rect 8636 13572 8660 13574
rect 8420 13552 8716 13572
rect 8772 13462 8800 13670
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6380 12374 6408 13126
rect 7392 12782 7420 13262
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12782 8800 13126
rect 8956 12918 8984 13262
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4448 11898 4476 12310
rect 6920 12232 6972 12238
rect 7024 12220 7052 12582
rect 8312 12374 8340 12582
rect 8420 12540 8716 12560
rect 8476 12538 8500 12540
rect 8556 12538 8580 12540
rect 8636 12538 8660 12540
rect 8498 12486 8500 12538
rect 8562 12486 8574 12538
rect 8636 12486 8638 12538
rect 8476 12484 8500 12486
rect 8556 12484 8580 12486
rect 8636 12484 8660 12486
rect 8420 12464 8716 12484
rect 9048 12442 9076 14894
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14618 9444 14758
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9692 14414 9720 14894
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 13938 9444 14214
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 6972 12192 7052 12220
rect 6920 12174 6972 12180
rect 4688 11996 4984 12016
rect 4744 11994 4768 11996
rect 4824 11994 4848 11996
rect 4904 11994 4928 11996
rect 4766 11942 4768 11994
rect 4830 11942 4842 11994
rect 4904 11942 4906 11994
rect 4744 11940 4768 11942
rect 4824 11940 4848 11942
rect 4904 11940 4928 11942
rect 4688 11920 4984 11940
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 6932 11694 6960 12174
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11218 6960 11630
rect 8220 11626 8248 12242
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8220 11354 8248 11562
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11286 8340 12106
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8420 11452 8716 11472
rect 8476 11450 8500 11452
rect 8556 11450 8580 11452
rect 8636 11450 8660 11452
rect 8498 11398 8500 11450
rect 8562 11398 8574 11450
rect 8636 11398 8638 11450
rect 8476 11396 8500 11398
rect 8556 11396 8580 11398
rect 8636 11396 8660 11398
rect 8420 11376 8716 11396
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 4688 10908 4984 10928
rect 4744 10906 4768 10908
rect 4824 10906 4848 10908
rect 4904 10906 4928 10908
rect 4766 10854 4768 10906
rect 4830 10854 4842 10906
rect 4904 10854 4906 10906
rect 4744 10852 4768 10854
rect 4824 10852 4848 10854
rect 4904 10852 4928 10854
rect 4688 10832 4984 10852
rect 6932 10674 6960 11154
rect 8680 10810 8708 11154
rect 8772 11150 8800 11834
rect 9048 11218 9076 12378
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 8312 10198 8340 10746
rect 8772 10606 8800 11086
rect 9140 11082 9168 12922
rect 9416 12918 9444 13874
rect 9692 13870 9720 14350
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9416 12238 9444 12854
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9692 11694 9720 13670
rect 9784 12986 9812 14418
rect 9876 13258 9904 14758
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9784 12170 9812 12650
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 9876 11778 9904 12582
rect 9784 11750 9904 11778
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8420 10364 8716 10384
rect 8476 10362 8500 10364
rect 8556 10362 8580 10364
rect 8636 10362 8660 10364
rect 8498 10310 8500 10362
rect 8562 10310 8574 10362
rect 8636 10310 8638 10362
rect 8476 10308 8500 10310
rect 8556 10308 8580 10310
rect 8636 10308 8660 10310
rect 8420 10288 8716 10308
rect 9324 10266 9352 11562
rect 9784 11150 9812 11750
rect 9968 11642 9996 13806
rect 10060 12442 10088 15506
rect 10336 14482 10364 15558
rect 11060 15506 11112 15512
rect 10508 15496 10560 15502
rect 10428 15456 10508 15484
rect 10428 14890 10456 15456
rect 10508 15438 10560 15444
rect 11072 15162 11100 15506
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10428 14618 10456 14826
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10152 13530 10180 13942
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 13326 10272 13874
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12850 10272 13262
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10152 12306 10180 12378
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10152 11762 10180 12242
rect 10336 11898 10364 13942
rect 10520 13841 10548 15098
rect 11348 14958 11376 20742
rect 12152 20700 12448 20720
rect 12208 20698 12232 20700
rect 12288 20698 12312 20700
rect 12368 20698 12392 20700
rect 12230 20646 12232 20698
rect 12294 20646 12306 20698
rect 12368 20646 12370 20698
rect 12208 20644 12232 20646
rect 12288 20644 12312 20646
rect 12368 20644 12392 20646
rect 12152 20624 12448 20644
rect 11888 20528 11940 20534
rect 12544 20516 12572 21354
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 20516 12664 20742
rect 11888 20470 11940 20476
rect 12452 20488 12664 20516
rect 11900 19961 11928 20470
rect 12452 20398 12480 20488
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 11886 19952 11942 19961
rect 11886 19887 11942 19896
rect 11702 19272 11758 19281
rect 11702 19207 11704 19216
rect 11756 19207 11758 19216
rect 11704 19178 11756 19184
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 18358 11468 19110
rect 11520 18828 11572 18834
rect 11716 18816 11744 19178
rect 11572 18788 11744 18816
rect 11520 18770 11572 18776
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11808 18222 11836 18566
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 16250 11836 16526
rect 11900 16454 11928 19887
rect 12452 19802 12480 20334
rect 12728 20040 12756 21542
rect 12898 21519 12954 21528
rect 13096 21418 13124 22102
rect 13188 22098 13216 23800
rect 13832 22438 13860 23800
rect 14476 23746 14504 23800
rect 14476 23718 14964 23746
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 13096 21146 13124 21354
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13188 20602 13216 21014
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12636 20012 12756 20040
rect 12532 19984 12584 19990
rect 12530 19952 12532 19961
rect 12584 19952 12586 19961
rect 12530 19887 12586 19896
rect 12452 19774 12572 19802
rect 12152 19612 12448 19632
rect 12208 19610 12232 19612
rect 12288 19610 12312 19612
rect 12368 19610 12392 19612
rect 12230 19558 12232 19610
rect 12294 19558 12306 19610
rect 12368 19558 12370 19610
rect 12208 19556 12232 19558
rect 12288 19556 12312 19558
rect 12368 19556 12392 19558
rect 12152 19536 12448 19556
rect 12440 19440 12492 19446
rect 12438 19408 12440 19417
rect 12492 19408 12494 19417
rect 12438 19343 12494 19352
rect 12544 19310 12572 19774
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18902 12572 19246
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12152 18524 12448 18544
rect 12208 18522 12232 18524
rect 12288 18522 12312 18524
rect 12368 18522 12392 18524
rect 12230 18470 12232 18522
rect 12294 18470 12306 18522
rect 12368 18470 12370 18522
rect 12208 18468 12232 18470
rect 12288 18468 12312 18470
rect 12368 18468 12392 18470
rect 12152 18448 12448 18468
rect 12544 18086 12572 18838
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12084 17338 12112 17750
rect 12440 17672 12492 17678
rect 12438 17640 12440 17649
rect 12492 17640 12494 17649
rect 12438 17575 12494 17584
rect 12152 17436 12448 17456
rect 12208 17434 12232 17436
rect 12288 17434 12312 17436
rect 12368 17434 12392 17436
rect 12230 17382 12232 17434
rect 12294 17382 12306 17434
rect 12368 17382 12370 17434
rect 12208 17380 12232 17382
rect 12288 17380 12312 17382
rect 12368 17380 12392 17382
rect 12152 17360 12448 17380
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12544 17066 12572 18022
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 15570 11928 16050
rect 11992 15978 12020 16526
rect 12152 16348 12448 16368
rect 12208 16346 12232 16348
rect 12288 16346 12312 16348
rect 12368 16346 12392 16348
rect 12230 16294 12232 16346
rect 12294 16294 12306 16346
rect 12368 16294 12370 16346
rect 12208 16292 12232 16294
rect 12288 16292 12312 16294
rect 12368 16292 12392 16294
rect 12152 16272 12448 16292
rect 12072 16040 12124 16046
rect 12532 16040 12584 16046
rect 12072 15982 12124 15988
rect 12452 16000 12532 16028
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11992 15706 12020 15914
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 12084 15366 12112 15982
rect 12452 15502 12480 16000
rect 12532 15982 12584 15988
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 12072 15360 12124 15366
rect 12452 15348 12480 15438
rect 12452 15320 12572 15348
rect 12072 15302 12124 15308
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10888 13938 10916 14418
rect 11348 13954 11376 14894
rect 11440 14482 11468 15302
rect 12152 15260 12448 15280
rect 12208 15258 12232 15260
rect 12288 15258 12312 15260
rect 12368 15258 12392 15260
rect 12230 15206 12232 15258
rect 12294 15206 12306 15258
rect 12368 15206 12370 15258
rect 12208 15204 12232 15206
rect 12288 15204 12312 15206
rect 12368 15204 12392 15206
rect 12152 15184 12448 15204
rect 12544 15162 12572 15320
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12636 15094 12664 20012
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19242 12756 19858
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12728 18630 12756 19178
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12728 17134 12756 17274
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16522 12756 16934
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12728 15706 12756 16458
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14482 12020 14826
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 10876 13932 10928 13938
rect 11348 13926 11468 13954
rect 10876 13874 10928 13880
rect 11440 13870 11468 13926
rect 11336 13864 11388 13870
rect 10506 13832 10562 13841
rect 11336 13806 11388 13812
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 10506 13767 10562 13776
rect 10692 13796 10744 13802
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9876 11614 9996 11642
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 4688 9820 4984 9840
rect 4744 9818 4768 9820
rect 4824 9818 4848 9820
rect 4904 9818 4928 9820
rect 4766 9766 4768 9818
rect 4830 9766 4842 9818
rect 4904 9766 4906 9818
rect 4744 9764 4768 9766
rect 4824 9764 4848 9766
rect 4904 9764 4928 9766
rect 4688 9744 4984 9764
rect 8420 9276 8716 9296
rect 8476 9274 8500 9276
rect 8556 9274 8580 9276
rect 8636 9274 8660 9276
rect 8498 9222 8500 9274
rect 8562 9222 8574 9274
rect 8636 9222 8638 9274
rect 8476 9220 8500 9222
rect 8556 9220 8580 9222
rect 8636 9220 8660 9222
rect 8420 9200 8716 9220
rect 9600 9042 9628 10066
rect 9692 9518 9720 11018
rect 9876 10266 9904 11614
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 10606 9996 11494
rect 10152 11354 10180 11698
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10060 11014 10088 11290
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10266 9996 10542
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10060 10062 10088 10950
rect 10152 10606 10180 11290
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10428 10266 10456 13670
rect 10520 13394 10548 13767
rect 10692 13738 10744 13744
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10704 13326 10732 13738
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13530 10916 13670
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12646 10640 13126
rect 10704 12782 10732 13262
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10704 12442 10732 12718
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10704 10810 10732 11154
rect 10980 11150 11008 12922
rect 11348 11354 11376 13806
rect 11808 12850 11836 14010
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12986 11928 13330
rect 11992 13258 12020 14418
rect 12152 14172 12448 14192
rect 12208 14170 12232 14172
rect 12288 14170 12312 14172
rect 12368 14170 12392 14172
rect 12230 14118 12232 14170
rect 12294 14118 12306 14170
rect 12368 14118 12370 14170
rect 12208 14116 12232 14118
rect 12288 14116 12312 14118
rect 12368 14116 12392 14118
rect 12152 14096 12448 14116
rect 12636 13938 12664 14758
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12728 14278 12756 14554
rect 12820 14482 12848 19790
rect 13004 18970 13032 19790
rect 13096 19514 13124 20538
rect 13372 19922 13400 21966
rect 13740 21690 13768 22034
rect 13820 21888 13872 21894
rect 14004 21888 14056 21894
rect 13872 21836 13952 21842
rect 13820 21830 13952 21836
rect 14004 21830 14056 21836
rect 13832 21814 13952 21830
rect 13924 21690 13952 21814
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13740 21078 13768 21626
rect 14016 21486 14044 21830
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13924 20806 13952 21422
rect 14200 21418 14228 22102
rect 14844 22098 14872 22374
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14936 22030 14964 23718
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14200 21146 14228 21354
rect 14476 21350 14504 21966
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13556 20058 13584 20334
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13740 19922 13768 20538
rect 14384 20398 14412 20742
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14200 20058 14228 20334
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13372 19825 13400 19858
rect 13358 19816 13414 19825
rect 13358 19751 13414 19760
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 13084 18760 13136 18766
rect 13136 18720 13308 18748
rect 13084 18702 13136 18708
rect 13280 18222 13308 18720
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12912 17882 12940 18022
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 13280 17542 13308 18158
rect 13372 17649 13400 19751
rect 13832 19514 13860 19994
rect 13912 19848 13964 19854
rect 13910 19816 13912 19825
rect 13964 19816 13966 19825
rect 13910 19751 13966 19760
rect 14384 19514 14412 20334
rect 14476 20312 14504 21286
rect 14556 20324 14608 20330
rect 14476 20284 14556 20312
rect 14556 20266 14608 20272
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14568 19786 14596 19994
rect 14752 19854 14780 21830
rect 14936 21690 14964 21830
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 15120 21078 15148 23800
rect 15764 23746 15792 23800
rect 17052 23746 17080 23800
rect 15488 23718 15792 23746
rect 16960 23718 17080 23746
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15108 21072 15160 21078
rect 14922 21040 14978 21049
rect 15108 21014 15160 21020
rect 14922 20975 14978 20984
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14752 19378 14780 19790
rect 14936 19553 14964 20975
rect 15120 20058 15148 21014
rect 15212 20942 15240 21898
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14922 19544 14978 19553
rect 14922 19479 14978 19488
rect 15016 19508 15068 19514
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18902 14044 19110
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14292 18834 14320 19246
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14384 18222 14412 19314
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18970 14504 19110
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14556 18828 14608 18834
rect 14556 18770 14608 18776
rect 14568 18426 14596 18770
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14016 17882 14044 18090
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14108 17882 14136 18022
rect 14476 17882 14504 18022
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13358 17640 13414 17649
rect 13358 17575 13414 17584
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17134 13308 17478
rect 13832 17338 13860 17682
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13556 16658 13584 17070
rect 14476 17066 14504 17818
rect 14648 17672 14700 17678
rect 14646 17640 14648 17649
rect 14700 17640 14702 17649
rect 14646 17575 14702 17584
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13268 14952 13320 14958
rect 13320 14912 13400 14940
rect 13268 14894 13320 14900
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 13372 14414 13400 14912
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12898 13832 12954 13841
rect 12624 13796 12676 13802
rect 12898 13767 12900 13776
rect 12624 13738 12676 13744
rect 12952 13767 12954 13776
rect 12900 13738 12952 13744
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13462 12480 13670
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12348 13320 12400 13326
rect 12084 13268 12348 13274
rect 12084 13262 12400 13268
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12084 13246 12388 13262
rect 12532 13252 12584 13258
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 11898 11560 12242
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11532 11354 11560 11834
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10704 10198 10732 10746
rect 11072 10606 11100 10950
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11072 10266 11100 10542
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 11716 9654 11744 12718
rect 12084 12714 12112 13246
rect 12532 13194 12584 13200
rect 12152 13084 12448 13104
rect 12208 13082 12232 13084
rect 12288 13082 12312 13084
rect 12368 13082 12392 13084
rect 12230 13030 12232 13082
rect 12294 13030 12306 13082
rect 12368 13030 12370 13082
rect 12208 13028 12232 13030
rect 12288 13028 12312 13030
rect 12368 13028 12392 13030
rect 12152 13008 12448 13028
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 12084 12442 12112 12650
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12152 11996 12448 12016
rect 12208 11994 12232 11996
rect 12288 11994 12312 11996
rect 12368 11994 12392 11996
rect 12230 11942 12232 11994
rect 12294 11942 12306 11994
rect 12368 11942 12370 11994
rect 12208 11940 12232 11942
rect 12288 11940 12312 11942
rect 12368 11940 12392 11942
rect 12152 11920 12448 11940
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 11354 11836 11562
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11808 10810 11836 11290
rect 12544 11150 12572 13194
rect 12636 12986 12664 13738
rect 13372 13734 13400 14350
rect 13464 14074 13492 15438
rect 13832 15434 13860 15846
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 14958 13860 15370
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13462 13400 13670
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 13004 12850 13032 13330
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12238 13032 12786
rect 13924 12646 13952 15302
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 12850 14044 14214
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12636 11898 12664 12174
rect 14108 11898 14136 16662
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16114 14228 16594
rect 14936 16250 14964 19479
rect 15016 19450 15068 19456
rect 15028 18222 15056 19450
rect 15106 18728 15162 18737
rect 15212 18698 15240 19994
rect 15304 19446 15332 22034
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15396 20602 15424 21286
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15488 19922 15516 23718
rect 15884 22332 16180 22352
rect 15940 22330 15964 22332
rect 16020 22330 16044 22332
rect 16100 22330 16124 22332
rect 15962 22278 15964 22330
rect 16026 22278 16038 22330
rect 16100 22278 16102 22330
rect 15940 22276 15964 22278
rect 16020 22276 16044 22278
rect 16100 22276 16124 22278
rect 15884 22256 16180 22276
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15580 20602 15608 20946
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15672 20466 15700 21830
rect 15750 21584 15806 21593
rect 15750 21519 15806 21528
rect 15764 21350 15792 21519
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15884 21244 16180 21264
rect 15940 21242 15964 21244
rect 16020 21242 16044 21244
rect 16100 21242 16124 21244
rect 15962 21190 15964 21242
rect 16026 21190 16038 21242
rect 16100 21190 16102 21242
rect 15940 21188 15964 21190
rect 16020 21188 16044 21190
rect 16100 21188 16124 21190
rect 15884 21168 16180 21188
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15672 20040 15700 20402
rect 15884 20156 16180 20176
rect 15940 20154 15964 20156
rect 16020 20154 16044 20156
rect 16100 20154 16124 20156
rect 15962 20102 15964 20154
rect 16026 20102 16038 20154
rect 16100 20102 16102 20154
rect 15940 20100 15964 20102
rect 16020 20100 16044 20102
rect 16100 20100 16124 20102
rect 15884 20080 16180 20100
rect 16224 20058 16252 21422
rect 16212 20052 16264 20058
rect 15672 20012 15884 20040
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15106 18663 15162 18672
rect 15200 18692 15252 18698
rect 15120 18630 15148 18663
rect 15200 18634 15252 18640
rect 15108 18624 15160 18630
rect 15108 18566 15160 18572
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 15028 17882 15056 18158
rect 15120 18068 15148 18566
rect 15304 18426 15332 19110
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15120 18040 15240 18068
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 16726 15148 17682
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 15212 16454 15240 18040
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15304 17134 15332 17682
rect 15396 17649 15424 19314
rect 15672 19009 15700 19858
rect 15856 19854 15884 20012
rect 16212 19994 16264 20000
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16316 19786 16344 21830
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16592 20398 16620 21286
rect 16868 20534 16896 21286
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16500 19922 16528 20198
rect 16578 20088 16634 20097
rect 16578 20023 16634 20032
rect 16592 19990 16620 20023
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16592 19854 16620 19926
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 19446 15884 19654
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 15658 19000 15714 19009
rect 15568 18964 15620 18970
rect 15658 18935 15714 18944
rect 15568 18906 15620 18912
rect 15580 18850 15608 18906
rect 15476 18828 15528 18834
rect 15580 18822 15700 18850
rect 15476 18770 15528 18776
rect 15488 17814 15516 18770
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 15382 17640 15438 17649
rect 15382 17575 15438 17584
rect 15488 17338 15516 17750
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16590 15332 17070
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15706 14228 15846
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14568 15162 14596 16050
rect 15212 15910 15240 16390
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15304 15706 15332 15982
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14476 14074 14504 14826
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13530 14596 14486
rect 14752 14278 14780 14758
rect 15120 14550 15148 14758
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13938 14780 14214
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14372 13388 14424 13394
rect 14372 13330 14424 13336
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14384 12986 14412 13330
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 11898 14320 12242
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11150 12940 11630
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12152 10908 12448 10928
rect 12208 10906 12232 10908
rect 12288 10906 12312 10908
rect 12368 10906 12392 10908
rect 12230 10854 12232 10906
rect 12294 10854 12306 10906
rect 12368 10854 12370 10906
rect 12208 10852 12232 10854
rect 12288 10852 12312 10854
rect 12368 10852 12392 10854
rect 12152 10832 12448 10852
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 12808 10600 12860 10606
rect 12912 10588 12940 11086
rect 12860 10560 12940 10588
rect 12808 10542 12860 10548
rect 12912 10062 12940 10560
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 4688 8732 4984 8752
rect 4744 8730 4768 8732
rect 4824 8730 4848 8732
rect 4904 8730 4928 8732
rect 4766 8678 4768 8730
rect 4830 8678 4842 8730
rect 4904 8678 4906 8730
rect 4744 8676 4768 8678
rect 4824 8676 4848 8678
rect 4904 8676 4928 8678
rect 4688 8656 4984 8676
rect 9600 8634 9628 8978
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7760 7954 7788 8366
rect 8420 8188 8716 8208
rect 8476 8186 8500 8188
rect 8556 8186 8580 8188
rect 8636 8186 8660 8188
rect 8498 8134 8500 8186
rect 8562 8134 8574 8186
rect 8636 8134 8638 8186
rect 8476 8132 8500 8134
rect 8556 8132 8580 8134
rect 8636 8132 8660 8134
rect 8420 8112 8716 8132
rect 9600 8090 9628 8570
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 4688 7644 4984 7664
rect 4744 7642 4768 7644
rect 4824 7642 4848 7644
rect 4904 7642 4928 7644
rect 4766 7590 4768 7642
rect 4830 7590 4842 7642
rect 4904 7590 4906 7642
rect 4744 7588 4768 7590
rect 4824 7588 4848 7590
rect 4904 7588 4928 7590
rect 4688 7568 4984 7588
rect 8220 7002 8248 7890
rect 9324 7410 9352 8026
rect 9600 7954 9628 8026
rect 9784 7954 9812 9590
rect 12084 9586 12112 9862
rect 12152 9820 12448 9840
rect 12208 9818 12232 9820
rect 12288 9818 12312 9820
rect 12368 9818 12392 9820
rect 12230 9766 12232 9818
rect 12294 9766 12306 9818
rect 12368 9766 12370 9818
rect 12208 9764 12232 9766
rect 12288 9764 12312 9766
rect 12368 9764 12392 9766
rect 12152 9744 12448 9764
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 9178 10916 9386
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8634 10548 8978
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10888 8430 10916 9114
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8430 11100 8774
rect 11532 8634 11560 8978
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 8430 11652 9318
rect 11702 8528 11758 8537
rect 12084 8514 12112 9522
rect 12912 9500 12940 9998
rect 12992 9512 13044 9518
rect 12912 9472 12992 9500
rect 12912 9042 12940 9472
rect 12992 9454 13044 9460
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12152 8732 12448 8752
rect 12208 8730 12232 8732
rect 12288 8730 12312 8732
rect 12368 8730 12392 8732
rect 12230 8678 12232 8730
rect 12294 8678 12306 8730
rect 12368 8678 12370 8730
rect 12208 8676 12232 8678
rect 12288 8676 12312 8678
rect 12368 8676 12392 8678
rect 12152 8656 12448 8676
rect 12636 8634 12664 8978
rect 13188 8838 13216 9386
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 9110 13584 9318
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 11992 8498 12112 8514
rect 11702 8463 11758 8472
rect 11980 8492 12112 8498
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11072 8022 11100 8366
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10888 7546 10916 7890
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7750 11008 7822
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8420 7100 8716 7120
rect 8476 7098 8500 7100
rect 8556 7098 8580 7100
rect 8636 7098 8660 7100
rect 8498 7046 8500 7098
rect 8562 7046 8574 7098
rect 8636 7046 8638 7098
rect 8476 7044 8500 7046
rect 8556 7044 8580 7046
rect 8636 7044 8660 7046
rect 8420 7024 8716 7044
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 9324 6866 9352 7346
rect 10888 6934 10916 7482
rect 10980 7342 11008 7686
rect 11164 7342 11192 7686
rect 11256 7410 11284 8298
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11716 7274 11744 8463
rect 12032 8486 12112 8492
rect 11980 8434 12032 8440
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 8090 12020 8230
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11808 7546 11836 7958
rect 12084 7886 12112 8486
rect 12162 8528 12218 8537
rect 12162 8463 12164 8472
rect 12216 8463 12218 8472
rect 12164 8434 12216 8440
rect 12636 7954 12664 8570
rect 13004 7954 13032 8774
rect 13188 8090 13216 8774
rect 13832 8362 13860 9454
rect 14016 8838 14044 11222
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14108 10810 14136 11154
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14200 9994 14228 11562
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 11082 14320 11154
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 10198 14320 11018
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10674 14412 10950
rect 14476 10810 14504 13330
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14844 12714 14872 13194
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14660 12442 14688 12650
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 15028 12374 15056 14010
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15304 13394 15332 13738
rect 15396 13394 15424 14962
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 12442 15148 12582
rect 15580 12458 15608 18634
rect 15672 18154 15700 18822
rect 15764 18748 15792 19314
rect 15884 19068 16180 19088
rect 15940 19066 15964 19068
rect 16020 19066 16044 19068
rect 16100 19066 16124 19068
rect 15962 19014 15964 19066
rect 16026 19014 16038 19066
rect 16100 19014 16102 19066
rect 15940 19012 15964 19014
rect 16020 19012 16044 19014
rect 16100 19012 16124 19014
rect 15884 18992 16180 19012
rect 15936 18760 15988 18766
rect 15764 18720 15936 18748
rect 15936 18702 15988 18708
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15884 17980 16180 18000
rect 15940 17978 15964 17980
rect 16020 17978 16044 17980
rect 16100 17978 16124 17980
rect 15962 17926 15964 17978
rect 16026 17926 16038 17978
rect 16100 17926 16102 17978
rect 15940 17924 15964 17926
rect 16020 17924 16044 17926
rect 16100 17924 16124 17926
rect 15884 17904 16180 17924
rect 15884 16892 16180 16912
rect 15940 16890 15964 16892
rect 16020 16890 16044 16892
rect 16100 16890 16124 16892
rect 15962 16838 15964 16890
rect 16026 16838 16038 16890
rect 16100 16838 16102 16890
rect 15940 16836 15964 16838
rect 16020 16836 16044 16838
rect 16100 16836 16124 16838
rect 15884 16816 16180 16836
rect 16224 16726 16252 19314
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16396 19304 16448 19310
rect 16960 19281 16988 23718
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17052 19990 17080 21286
rect 17144 20602 17172 21286
rect 17328 21146 17356 21490
rect 17420 21457 17448 21830
rect 17696 21690 17724 23800
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17406 21448 17462 21457
rect 17406 21383 17462 21392
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17236 20466 17264 21014
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 17420 19854 17448 20742
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17512 20097 17540 20334
rect 17498 20088 17554 20097
rect 17498 20023 17554 20032
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 16946 19272 17002 19281
rect 16448 19252 16528 19258
rect 16396 19246 16528 19252
rect 16316 18986 16344 19246
rect 16408 19230 16528 19246
rect 16316 18958 16436 18986
rect 16302 18864 16358 18873
rect 16302 18799 16358 18808
rect 16316 18766 16344 18799
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16408 18426 16436 18958
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16500 18306 16528 19230
rect 16580 19236 16632 19242
rect 16946 19207 17002 19216
rect 16580 19178 16632 19184
rect 16592 18970 16620 19178
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16856 18760 16908 18766
rect 16854 18728 16856 18737
rect 16908 18728 16910 18737
rect 16854 18663 16910 18672
rect 16408 18278 16528 18306
rect 16408 18222 16436 18278
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 17746 16436 18158
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16684 17882 16712 18022
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 17052 17610 17080 19110
rect 17144 18766 17172 19654
rect 17604 19446 17632 19790
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 17882 17172 18702
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16114 17080 16390
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 15672 15162 15700 16050
rect 15884 15804 16180 15824
rect 15940 15802 15964 15804
rect 16020 15802 16044 15804
rect 16100 15802 16124 15804
rect 15962 15750 15964 15802
rect 16026 15750 16038 15802
rect 16100 15750 16102 15802
rect 15940 15748 15964 15750
rect 16020 15748 16044 15750
rect 16100 15748 16124 15750
rect 15884 15728 16180 15748
rect 17052 15638 17080 16050
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15672 14618 15700 14826
rect 15884 14716 16180 14736
rect 15940 14714 15964 14716
rect 16020 14714 16044 14716
rect 16100 14714 16124 14716
rect 15962 14662 15964 14714
rect 16026 14662 16038 14714
rect 16100 14662 16102 14714
rect 15940 14660 15964 14662
rect 16020 14660 16044 14662
rect 16100 14660 16124 14662
rect 15884 14640 16180 14660
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 16224 14414 16252 15030
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 12866 15700 14282
rect 15764 12986 15792 14350
rect 15884 13628 16180 13648
rect 15940 13626 15964 13628
rect 16020 13626 16044 13628
rect 16100 13626 16124 13628
rect 15962 13574 15964 13626
rect 16026 13574 16038 13626
rect 16100 13574 16102 13626
rect 15940 13572 15964 13574
rect 16020 13572 16044 13574
rect 16100 13572 16124 13574
rect 15884 13552 16180 13572
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15672 12838 15792 12866
rect 15856 12850 15884 13330
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 15571 12442 15608 12458
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15396 11830 15424 12106
rect 15488 11898 15516 12106
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14568 10606 14596 11494
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14660 10130 14688 10950
rect 14936 10674 14964 11562
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15120 10606 15148 11154
rect 15212 11150 15240 11698
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15014 10160 15070 10169
rect 14648 10124 14700 10130
rect 15014 10095 15070 10104
rect 14648 10066 14700 10072
rect 15028 10062 15056 10095
rect 15120 10062 15148 10542
rect 15396 10282 15424 11766
rect 15580 11694 15608 12038
rect 15672 11898 15700 12174
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15764 11626 15792 12838
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15884 12540 16180 12560
rect 15940 12538 15964 12540
rect 16020 12538 16044 12540
rect 16100 12538 16124 12540
rect 15962 12486 15964 12538
rect 16026 12486 16038 12538
rect 16100 12486 16102 12538
rect 15940 12484 15964 12486
rect 16020 12484 16044 12486
rect 16100 12484 16124 12486
rect 15884 12464 16180 12484
rect 16224 12442 16252 13126
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11694 16160 12174
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15884 11452 16180 11472
rect 15940 11450 15964 11452
rect 16020 11450 16044 11452
rect 16100 11450 16124 11452
rect 15962 11398 15964 11450
rect 16026 11398 16038 11450
rect 16100 11398 16102 11450
rect 15940 11396 15964 11398
rect 16020 11396 16044 11398
rect 16100 11396 16124 11398
rect 15884 11376 16180 11396
rect 16224 10538 16252 11494
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 15884 10364 16180 10384
rect 15940 10362 15964 10364
rect 16020 10362 16044 10364
rect 16100 10362 16124 10364
rect 15962 10310 15964 10362
rect 16026 10310 16038 10362
rect 16100 10310 16102 10362
rect 15940 10308 15964 10310
rect 16020 10308 16044 10310
rect 16100 10308 16124 10310
rect 15884 10288 16180 10308
rect 15396 10254 15516 10282
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14922 9072 14978 9081
rect 15120 9042 15148 9998
rect 15396 9654 15424 10066
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15488 9450 15516 10254
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 14922 9007 14924 9016
rect 14976 9007 14978 9016
rect 15108 9036 15160 9042
rect 14924 8978 14976 8984
rect 15108 8978 15160 8984
rect 15120 8945 15148 8978
rect 15200 8968 15252 8974
rect 15106 8936 15162 8945
rect 14464 8900 14516 8906
rect 15396 8922 15424 9318
rect 15252 8916 15424 8922
rect 15200 8910 15424 8916
rect 15212 8894 15424 8910
rect 15106 8871 15162 8880
rect 14464 8842 14516 8848
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 4688 6556 4984 6576
rect 4744 6554 4768 6556
rect 4824 6554 4848 6556
rect 4904 6554 4928 6556
rect 4766 6502 4768 6554
rect 4830 6502 4842 6554
rect 4904 6502 4906 6554
rect 4744 6500 4768 6502
rect 4824 6500 4848 6502
rect 4904 6500 4928 6502
rect 4688 6480 4984 6500
rect 9324 6458 9352 6802
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8420 6012 8716 6032
rect 8476 6010 8500 6012
rect 8556 6010 8580 6012
rect 8636 6010 8660 6012
rect 8498 5958 8500 6010
rect 8562 5958 8574 6010
rect 8636 5958 8638 6010
rect 8476 5956 8500 5958
rect 8556 5956 8580 5958
rect 8636 5956 8660 5958
rect 8420 5936 8716 5956
rect 9324 5778 9352 6394
rect 10336 6254 10364 6598
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 11072 5846 11100 6394
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 4688 5468 4984 5488
rect 4744 5466 4768 5468
rect 4824 5466 4848 5468
rect 4904 5466 4928 5468
rect 4766 5414 4768 5466
rect 4830 5414 4842 5466
rect 4904 5414 4906 5466
rect 4744 5412 4768 5414
rect 4824 5412 4848 5414
rect 4904 5412 4928 5414
rect 4688 5392 4984 5412
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 8420 4924 8716 4944
rect 8476 4922 8500 4924
rect 8556 4922 8580 4924
rect 8636 4922 8660 4924
rect 8498 4870 8500 4922
rect 8562 4870 8574 4922
rect 8636 4870 8638 4922
rect 8476 4868 8500 4870
rect 8556 4868 8580 4870
rect 8636 4868 8660 4870
rect 8420 4848 8716 4868
rect 11164 4758 11192 4966
rect 11256 4826 11284 6598
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5914 11376 6122
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11348 5234 11376 5850
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11440 4622 11468 7210
rect 12084 6934 12112 7822
rect 12152 7644 12448 7664
rect 12208 7642 12232 7644
rect 12288 7642 12312 7644
rect 12368 7642 12392 7644
rect 12230 7590 12232 7642
rect 12294 7590 12306 7642
rect 12368 7590 12370 7642
rect 12208 7588 12232 7590
rect 12288 7588 12312 7590
rect 12368 7588 12392 7590
rect 12152 7568 12448 7588
rect 13096 7410 13124 7822
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 6934 12664 7210
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11532 6458 11560 6802
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5846 11836 6054
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11808 5098 11836 5782
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11992 4554 12020 6802
rect 12152 6556 12448 6576
rect 12208 6554 12232 6556
rect 12288 6554 12312 6556
rect 12368 6554 12392 6556
rect 12230 6502 12232 6554
rect 12294 6502 12306 6554
rect 12368 6502 12370 6554
rect 12208 6500 12232 6502
rect 12288 6500 12312 6502
rect 12368 6500 12392 6502
rect 12152 6480 12448 6500
rect 12544 6458 12572 6870
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12728 5846 12756 6802
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 5914 12848 6734
rect 12912 6662 12940 7142
rect 13280 7002 13308 7278
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 13004 6458 13032 6734
rect 13832 6662 13860 8298
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7342 14044 7686
rect 14108 7546 14136 7890
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 6866 14044 7142
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12152 5468 12448 5488
rect 12208 5466 12232 5468
rect 12288 5466 12312 5468
rect 12368 5466 12392 5468
rect 12230 5414 12232 5466
rect 12294 5414 12306 5466
rect 12368 5414 12370 5466
rect 12208 5412 12232 5414
rect 12288 5412 12312 5414
rect 12368 5412 12392 5414
rect 12152 5392 12448 5412
rect 12820 5098 12848 5850
rect 12912 5778 12940 6054
rect 13004 5778 13032 6394
rect 13832 6254 13860 6598
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5914 14044 6122
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12912 5030 12940 5714
rect 13004 5166 13032 5714
rect 13740 5370 13768 5782
rect 14200 5370 14228 6190
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14292 5166 14320 8774
rect 14476 8430 14504 8842
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14648 8628 14700 8634
rect 14568 8588 14648 8616
rect 14568 8498 14596 8588
rect 14648 8570 14700 8576
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14648 8424 14700 8430
rect 14700 8372 14780 8378
rect 14648 8366 14780 8372
rect 14660 8350 14780 8366
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14384 8090 14412 8230
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14476 7478 14504 7890
rect 14660 7818 14688 8230
rect 14752 7993 14780 8350
rect 15120 8294 15148 8774
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14922 8120 14978 8129
rect 14922 8055 14978 8064
rect 14936 8022 14964 8055
rect 14924 8016 14976 8022
rect 14738 7984 14794 7993
rect 14924 7958 14976 7964
rect 14738 7919 14794 7928
rect 15396 7886 15424 8894
rect 15580 8634 15608 10066
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 9081 15700 9318
rect 15884 9276 16180 9296
rect 15940 9274 15964 9276
rect 16020 9274 16044 9276
rect 16100 9274 16124 9276
rect 15962 9222 15964 9274
rect 16026 9222 16038 9274
rect 16100 9222 16102 9274
rect 15940 9220 15964 9222
rect 16020 9220 16044 9222
rect 16100 9220 16124 9222
rect 15884 9200 16180 9220
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15658 9072 15714 9081
rect 15658 9007 15714 9016
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15764 8537 15792 9114
rect 15750 8528 15806 8537
rect 15750 8463 15806 8472
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 8129 15608 8366
rect 15884 8188 16180 8208
rect 15940 8186 15964 8188
rect 16020 8186 16044 8188
rect 16100 8186 16124 8188
rect 15962 8134 15964 8186
rect 16026 8134 16038 8186
rect 16100 8134 16102 8186
rect 15940 8132 15964 8134
rect 16020 8132 16044 8134
rect 16100 8132 16124 8134
rect 15566 8120 15622 8129
rect 15884 8112 16180 8132
rect 15566 8055 15622 8064
rect 16026 7984 16082 7993
rect 16026 7919 16028 7928
rect 16080 7919 16082 7928
rect 16028 7890 16080 7896
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7562 14596 7686
rect 14568 7534 14780 7562
rect 14752 7478 14780 7534
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14476 7206 14504 7414
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 7002 14780 7142
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14384 5914 14412 6938
rect 15120 6730 15148 7278
rect 15304 7206 15332 7754
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14752 5914 14780 6122
rect 15304 5914 15332 7142
rect 15488 6458 15516 7210
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15580 5846 15608 6598
rect 15672 5914 15700 7822
rect 15884 7100 16180 7120
rect 15940 7098 15964 7100
rect 16020 7098 16044 7100
rect 16100 7098 16124 7100
rect 15962 7046 15964 7098
rect 16026 7046 16038 7098
rect 16100 7046 16102 7098
rect 15940 7044 15964 7046
rect 16020 7044 16044 7046
rect 16100 7044 16124 7046
rect 15884 7024 16180 7044
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15856 6458 15884 6802
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15884 6012 16180 6032
rect 15940 6010 15964 6012
rect 16020 6010 16044 6012
rect 16100 6010 16124 6012
rect 15962 5958 15964 6010
rect 16026 5958 16038 6010
rect 16100 5958 16102 6010
rect 15940 5956 15964 5958
rect 16020 5956 16044 5958
rect 16100 5956 16124 5958
rect 15884 5936 16180 5956
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 16316 5098 16344 14962
rect 16408 14482 16436 15506
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 15026 16712 15302
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16776 14958 16804 15438
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16408 13802 16436 14418
rect 16500 13870 16528 14758
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16592 13530 16620 14418
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16408 11762 16436 12786
rect 16592 12782 16620 13466
rect 16868 12986 16896 14758
rect 17052 14618 17080 15302
rect 17144 14890 17172 15846
rect 17236 15570 17264 16594
rect 17328 16250 17356 18770
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17236 14906 17264 15506
rect 17604 15366 17632 16594
rect 17696 15978 17724 20470
rect 17880 20262 17908 21898
rect 18064 21554 18092 22102
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18248 21486 18276 21830
rect 18340 21486 18368 23800
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18064 20466 18092 20878
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19990 17908 20198
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17972 19310 18000 19654
rect 18064 19514 18092 19926
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17868 17672 17920 17678
rect 17972 17660 18000 19246
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18064 17746 18092 18226
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17920 17632 18000 17660
rect 17868 17614 17920 17620
rect 18064 17202 18092 17682
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16726 18092 17138
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 18064 15570 18092 15982
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17132 14884 17184 14890
rect 17236 14878 17356 14906
rect 17132 14826 17184 14832
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 13818 17080 14214
rect 17052 13790 17172 13818
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13546 17080 13670
rect 16960 13530 17080 13546
rect 16948 13524 17080 13530
rect 17000 13518 17080 13524
rect 16948 13466 17000 13472
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 17052 12646 17080 13518
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17144 12374 17172 13790
rect 17236 12918 17264 14758
rect 17328 14346 17356 14878
rect 17696 14362 17724 15302
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17604 14334 17724 14362
rect 17604 13870 17632 14334
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17328 12442 17356 13670
rect 17604 12986 17632 13806
rect 17696 13462 17724 14214
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17696 12714 17724 13398
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16500 11898 16528 12242
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16408 11218 16436 11562
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10810 16436 11154
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 9994 16436 10474
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 9042 16436 9318
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16500 8974 16528 10542
rect 16684 10130 16712 12310
rect 17788 12238 17816 13942
rect 17880 12918 17908 14214
rect 17972 14074 18000 15030
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14074 18092 14894
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17972 12782 18000 13126
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11694 17172 12038
rect 17972 11830 18000 12174
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16868 10470 16896 11494
rect 16960 11354 16988 11494
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16960 10538 16988 11290
rect 17972 11218 18000 11630
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16856 10464 16908 10470
rect 17052 10418 17080 10474
rect 16856 10406 16908 10412
rect 16960 10390 17080 10418
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16868 9518 16896 9930
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16488 8968 16540 8974
rect 16486 8936 16488 8945
rect 16540 8936 16542 8945
rect 16486 8871 16542 8880
rect 16776 8838 16804 9046
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16684 8634 16712 8774
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16408 8090 16436 8298
rect 16488 8288 16540 8294
rect 16592 8276 16620 8502
rect 16868 8498 16896 9454
rect 16960 9450 16988 10390
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 17052 8566 17080 9998
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16540 8248 16620 8276
rect 16764 8288 16816 8294
rect 16488 8230 16540 8236
rect 16764 8230 16816 8236
rect 16500 8090 16528 8230
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16408 7868 16436 8026
rect 16776 7954 16804 8230
rect 17420 7993 17448 9998
rect 17972 9722 18000 11154
rect 18064 10606 18092 12038
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17972 9518 18000 9658
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17512 8566 17540 9318
rect 17604 8634 17632 9318
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17604 8090 17632 8434
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17406 7984 17462 7993
rect 16764 7948 16816 7954
rect 17406 7919 17462 7928
rect 16764 7890 16816 7896
rect 16488 7880 16540 7886
rect 16408 7840 16488 7868
rect 16488 7822 16540 7828
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16408 5710 16436 7482
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16500 6730 16528 7210
rect 16592 6866 16620 7278
rect 16684 7206 16712 7346
rect 16776 7342 16804 7890
rect 17420 7886 17448 7919
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 17420 6866 17448 7346
rect 17880 7342 17908 8978
rect 17972 8498 18000 9046
rect 18064 8838 18092 9590
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 7546 18000 8434
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 7954 18092 8230
rect 18156 8022 18184 19450
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 17814 18460 18566
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18248 12238 18276 14418
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18340 12186 18368 13806
rect 18432 12594 18460 17750
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18524 14482 18552 15506
rect 18616 15094 18644 21490
rect 18984 19514 19012 23800
rect 19628 22930 19656 23800
rect 19352 22902 19656 22930
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19076 19922 19104 20470
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19154 19544 19210 19553
rect 18972 19508 19024 19514
rect 19154 19479 19156 19488
rect 18972 19450 19024 19456
rect 19208 19479 19210 19488
rect 19156 19450 19208 19456
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 18834 19012 19246
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18984 18426 19012 18770
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 19076 16794 19104 17002
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18708 15026 18736 16662
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18524 14226 18552 14418
rect 18604 14272 18656 14278
rect 18524 14220 18604 14226
rect 18524 14214 18656 14220
rect 18524 14198 18644 14214
rect 18524 13802 18552 14198
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18524 13530 18552 13738
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18524 13190 18552 13466
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12714 18552 13126
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18432 12566 18552 12594
rect 18340 12158 18460 12186
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18248 9926 18276 9998
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18248 9330 18276 9658
rect 18340 9518 18368 11018
rect 18432 10169 18460 12158
rect 18418 10160 18474 10169
rect 18418 10095 18474 10104
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18432 9330 18460 9386
rect 18248 9302 18460 9330
rect 18248 8974 18276 9302
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8498 18276 8910
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18432 7954 18460 8230
rect 18524 8090 18552 12566
rect 18800 12238 18828 14826
rect 19260 13530 19288 21354
rect 19352 19417 19380 22902
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19444 20602 19472 22034
rect 19616 21788 19912 21808
rect 19672 21786 19696 21788
rect 19752 21786 19776 21788
rect 19832 21786 19856 21788
rect 19694 21734 19696 21786
rect 19758 21734 19770 21786
rect 19832 21734 19834 21786
rect 19672 21732 19696 21734
rect 19752 21732 19776 21734
rect 19832 21732 19856 21734
rect 19616 21712 19912 21732
rect 20272 21622 20300 23800
rect 20260 21616 20312 21622
rect 20260 21558 20312 21564
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19536 20398 19564 20742
rect 19616 20700 19912 20720
rect 19672 20698 19696 20700
rect 19752 20698 19776 20700
rect 19832 20698 19856 20700
rect 19694 20646 19696 20698
rect 19758 20646 19770 20698
rect 19832 20646 19834 20698
rect 19672 20644 19696 20646
rect 19752 20644 19776 20646
rect 19832 20644 19856 20646
rect 19616 20624 19912 20644
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19338 19408 19394 19417
rect 19338 19343 19394 19352
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19352 17610 19380 19178
rect 19444 17882 19472 19790
rect 19616 19612 19912 19632
rect 19672 19610 19696 19612
rect 19752 19610 19776 19612
rect 19832 19610 19856 19612
rect 19694 19558 19696 19610
rect 19758 19558 19770 19610
rect 19832 19558 19834 19610
rect 19672 19556 19696 19558
rect 19752 19556 19776 19558
rect 19832 19556 19856 19558
rect 19616 19536 19912 19556
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19536 18154 19564 19110
rect 19996 18970 20024 20198
rect 20916 19990 20944 23800
rect 21560 21010 21588 23800
rect 21836 21622 21864 24239
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 21914 23624 21970 23633
rect 21914 23559 21970 23568
rect 21928 21690 21956 23559
rect 22006 22944 22062 22953
rect 22006 22879 22062 22888
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 22020 21146 22048 22879
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 22204 20330 22232 23800
rect 22848 23746 22876 23800
rect 22848 23718 22968 23746
rect 22466 21584 22522 21593
rect 22466 21519 22522 21528
rect 22480 20602 22508 21519
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 22112 19938 22140 20198
rect 22388 20074 22416 20402
rect 22466 20224 22522 20233
rect 22466 20159 22522 20168
rect 22296 20058 22416 20074
rect 22480 20058 22508 20159
rect 22284 20052 22416 20058
rect 22336 20046 22416 20052
rect 22468 20052 22520 20058
rect 22284 19994 22336 20000
rect 22468 19994 22520 20000
rect 22376 19984 22428 19990
rect 22112 19922 22324 19938
rect 22376 19926 22428 19932
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 22112 19916 22336 19922
rect 22112 19910 22284 19916
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19616 18524 19912 18544
rect 19672 18522 19696 18524
rect 19752 18522 19776 18524
rect 19832 18522 19856 18524
rect 19694 18470 19696 18522
rect 19758 18470 19770 18522
rect 19832 18470 19834 18522
rect 19672 18468 19696 18470
rect 19752 18468 19776 18470
rect 19832 18468 19856 18470
rect 19616 18448 19912 18468
rect 19996 18426 20024 18770
rect 20088 18426 20116 19858
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20364 18970 20392 19178
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20364 18222 20392 18906
rect 20456 18358 20484 19654
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18766 20852 19246
rect 21008 18834 21036 19654
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18902 21128 19110
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21178 18864 21234 18873
rect 20996 18828 21048 18834
rect 21178 18799 21234 18808
rect 20996 18770 21048 18776
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20640 18290 20668 18362
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19536 17882 19564 18090
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19444 17338 19472 17682
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 19616 17436 19912 17456
rect 19672 17434 19696 17436
rect 19752 17434 19776 17436
rect 19832 17434 19856 17436
rect 19694 17382 19696 17434
rect 19758 17382 19770 17434
rect 19832 17382 19834 17434
rect 19672 17380 19696 17382
rect 19752 17380 19776 17382
rect 19832 17380 19856 17382
rect 19616 17360 19912 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 20180 17202 20208 17614
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16726 19748 16934
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 15978 19380 16526
rect 19444 16250 19472 16594
rect 20180 16590 20208 17138
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 19616 16348 19912 16368
rect 19672 16346 19696 16348
rect 19752 16346 19776 16348
rect 19832 16346 19856 16348
rect 19694 16294 19696 16346
rect 19758 16294 19770 16346
rect 19832 16294 19834 16346
rect 19672 16292 19696 16294
rect 19752 16292 19776 16294
rect 19832 16292 19856 16294
rect 19616 16272 19912 16292
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 20180 16114 20208 16526
rect 20272 16522 20300 17682
rect 20640 17678 20668 18226
rect 20824 18154 20852 18702
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 21192 17814 21220 18799
rect 21180 17808 21232 17814
rect 21180 17750 21232 17756
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20456 17134 20484 17478
rect 21376 17338 21404 19858
rect 21916 19780 21968 19786
rect 21916 19722 21968 19728
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18222 21680 19110
rect 21928 18222 21956 19722
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21468 17678 21496 18158
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20258 16280 20314 16289
rect 20258 16215 20314 16224
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19352 15706 19380 15914
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19904 15638 19932 15846
rect 19892 15632 19944 15638
rect 19338 15600 19394 15609
rect 19892 15574 19944 15580
rect 19996 15570 20024 15846
rect 19338 15535 19394 15544
rect 19984 15564 20036 15570
rect 19352 15366 19380 15535
rect 19984 15506 20036 15512
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19616 15260 19912 15280
rect 19672 15258 19696 15260
rect 19752 15258 19776 15260
rect 19832 15258 19856 15260
rect 19694 15206 19696 15258
rect 19758 15206 19770 15258
rect 19832 15206 19834 15258
rect 19672 15204 19696 15206
rect 19752 15204 19776 15206
rect 19832 15204 19856 15206
rect 19616 15184 19912 15204
rect 19996 15162 20024 15506
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 19352 14929 19380 15098
rect 20180 15026 20208 16050
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19338 14920 19394 14929
rect 19338 14855 19394 14864
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19352 14550 19380 14758
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19352 14385 19380 14486
rect 19444 14482 19472 14758
rect 19812 14618 19840 14826
rect 20272 14618 20300 16215
rect 20916 16114 20944 16390
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19338 14376 19394 14385
rect 19338 14311 19394 14320
rect 19444 14074 19472 14418
rect 19616 14172 19912 14192
rect 19672 14170 19696 14172
rect 19752 14170 19776 14172
rect 19832 14170 19856 14172
rect 19694 14118 19696 14170
rect 19758 14118 19770 14170
rect 19832 14118 19834 14170
rect 19672 14116 19696 14118
rect 19752 14116 19776 14118
rect 19832 14116 19856 14118
rect 19616 14096 19912 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 20272 13938 20300 14554
rect 20364 14278 20392 15982
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20456 15570 20484 15846
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20824 15162 20852 15846
rect 21008 15706 21036 16934
rect 21468 16658 21496 17614
rect 21652 17066 21680 18158
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21548 17060 21600 17066
rect 21548 17002 21600 17008
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21192 16250 21220 16594
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21560 16096 21588 17002
rect 21744 16726 21772 17818
rect 21836 17814 21864 18022
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21836 17134 21864 17750
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21928 16454 21956 18158
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21640 16108 21692 16114
rect 21560 16068 21640 16096
rect 21640 16050 21692 16056
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 21376 14958 21404 15438
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21376 14414 21404 14894
rect 21560 14482 21588 15846
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19616 13796 19668 13802
rect 19536 13756 19616 13784
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18708 11082 18736 11562
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 10470 18736 11018
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18616 10130 18644 10406
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 9042 18644 9454
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18708 8922 18736 10406
rect 18616 8894 18736 8922
rect 18616 8616 18644 8894
rect 18696 8628 18748 8634
rect 18616 8588 18696 8616
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7954 18644 8588
rect 18696 8570 18748 8576
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 18064 7206 18092 7890
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16500 5778 16528 6666
rect 17604 6322 17632 7142
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5098 16436 5646
rect 17236 5370 17264 5714
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 15884 4924 16180 4944
rect 15940 4922 15964 4924
rect 16020 4922 16044 4924
rect 16100 4922 16124 4924
rect 15962 4870 15964 4922
rect 16026 4870 16038 4922
rect 16100 4870 16102 4922
rect 15940 4868 15964 4870
rect 16020 4868 16044 4870
rect 16100 4868 16124 4870
rect 15884 4848 16180 4868
rect 16408 4706 16436 5034
rect 17788 5012 17816 5510
rect 17880 5166 17908 5510
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17868 5024 17920 5030
rect 17788 4984 17868 5012
rect 17788 4758 17816 4984
rect 17868 4966 17920 4972
rect 17776 4752 17828 4758
rect 16408 4690 16528 4706
rect 17776 4694 17828 4700
rect 16408 4684 16540 4690
rect 16408 4678 16488 4684
rect 16488 4626 16540 4632
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 4688 4380 4984 4400
rect 4744 4378 4768 4380
rect 4824 4378 4848 4380
rect 4904 4378 4928 4380
rect 4766 4326 4768 4378
rect 4830 4326 4842 4378
rect 4904 4326 4906 4378
rect 4744 4324 4768 4326
rect 4824 4324 4848 4326
rect 4904 4324 4928 4326
rect 4688 4304 4984 4324
rect 12152 4380 12448 4400
rect 12208 4378 12232 4380
rect 12288 4378 12312 4380
rect 12368 4378 12392 4380
rect 12230 4326 12232 4378
rect 12294 4326 12306 4378
rect 12368 4326 12370 4378
rect 12208 4324 12232 4326
rect 12288 4324 12312 4326
rect 12368 4324 12392 4326
rect 12152 4304 12448 4324
rect 16500 4010 16528 4626
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4078 17816 4422
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 8420 3836 8716 3856
rect 8476 3834 8500 3836
rect 8556 3834 8580 3836
rect 8636 3834 8660 3836
rect 8498 3782 8500 3834
rect 8562 3782 8574 3834
rect 8636 3782 8638 3834
rect 8476 3780 8500 3782
rect 8556 3780 8580 3782
rect 8636 3780 8660 3782
rect 8420 3760 8716 3780
rect 15884 3836 16180 3856
rect 15940 3834 15964 3836
rect 16020 3834 16044 3836
rect 16100 3834 16124 3836
rect 15962 3782 15964 3834
rect 16026 3782 16038 3834
rect 16100 3782 16102 3834
rect 15940 3780 15964 3782
rect 16020 3780 16044 3782
rect 16100 3780 16124 3782
rect 15884 3760 16180 3780
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2332 3194 2360 3538
rect 16500 3534 16528 3946
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 3670 18000 3878
rect 18064 3738 18092 7142
rect 18156 7002 18184 7210
rect 18616 7002 18644 7890
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18156 6322 18184 6938
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18248 6254 18276 6734
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18248 4826 18276 5714
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5370 18368 5646
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18248 3942 18276 4626
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 4688 3292 4984 3312
rect 4744 3290 4768 3292
rect 4824 3290 4848 3292
rect 4904 3290 4928 3292
rect 4766 3238 4768 3290
rect 4830 3238 4842 3290
rect 4904 3238 4906 3290
rect 4744 3236 4768 3238
rect 4824 3236 4848 3238
rect 4904 3236 4928 3238
rect 4688 3216 4984 3236
rect 12152 3292 12448 3312
rect 12208 3290 12232 3292
rect 12288 3290 12312 3292
rect 12368 3290 12392 3292
rect 12230 3238 12232 3290
rect 12294 3238 12306 3290
rect 12368 3238 12370 3290
rect 12208 3236 12232 3238
rect 12288 3236 12312 3238
rect 12368 3236 12392 3238
rect 12152 3216 12448 3236
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 2044 3120 2096 3126
rect 1950 3088 2006 3097
rect 2044 3062 2096 3068
rect 1950 3023 1952 3032
rect 2004 3023 2006 3032
rect 1952 2994 2004 3000
rect 2056 800 2084 3062
rect 2516 2990 2544 3130
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 4688 2204 4984 2224
rect 4744 2202 4768 2204
rect 4824 2202 4848 2204
rect 4904 2202 4928 2204
rect 4766 2150 4768 2202
rect 4830 2150 4842 2202
rect 4904 2150 4906 2202
rect 4744 2148 4768 2150
rect 4824 2148 4848 2150
rect 4904 2148 4928 2150
rect 4688 2128 4984 2148
rect 6104 800 6132 2926
rect 8420 2748 8716 2768
rect 8476 2746 8500 2748
rect 8556 2746 8580 2748
rect 8636 2746 8660 2748
rect 8498 2694 8500 2746
rect 8562 2694 8574 2746
rect 8636 2694 8638 2746
rect 8476 2692 8500 2694
rect 8556 2692 8580 2694
rect 8636 2692 8660 2694
rect 8420 2672 8716 2692
rect 10244 800 10272 3130
rect 16500 2990 16528 3470
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 17788 2922 17816 3334
rect 17880 3194 17908 3538
rect 17960 3528 18012 3534
rect 18012 3476 18092 3482
rect 17960 3470 18092 3476
rect 17972 3454 18092 3470
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17880 2990 17908 3130
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 18064 2854 18092 3454
rect 18892 3126 18920 13466
rect 19536 13190 19564 13756
rect 19616 13738 19668 13744
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19536 12782 19564 13126
rect 19616 13084 19912 13104
rect 19672 13082 19696 13084
rect 19752 13082 19776 13084
rect 19832 13082 19856 13084
rect 19694 13030 19696 13082
rect 19758 13030 19770 13082
rect 19832 13030 19834 13082
rect 19672 13028 19696 13030
rect 19752 13028 19776 13030
rect 19832 13028 19856 13030
rect 19616 13008 19912 13028
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 10606 19012 12038
rect 19260 11762 19288 12242
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19352 11694 19380 12106
rect 19444 11898 19472 12242
rect 19628 12238 19656 12582
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19430 11656 19486 11665
rect 19430 11591 19486 11600
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11286 19104 11494
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19076 10674 19104 11222
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 19352 10538 19380 11222
rect 19444 11014 19472 11591
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19444 10282 19472 10610
rect 19536 10606 19564 12174
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19616 11996 19912 12016
rect 19672 11994 19696 11996
rect 19752 11994 19776 11996
rect 19832 11994 19856 11996
rect 19694 11942 19696 11994
rect 19758 11942 19770 11994
rect 19832 11942 19834 11994
rect 19672 11940 19696 11942
rect 19752 11940 19776 11942
rect 19832 11940 19856 11942
rect 19616 11920 19912 11940
rect 19996 11762 20024 12038
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 20088 11694 20116 13806
rect 20260 13728 20312 13734
rect 20364 13716 20392 14214
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20312 13688 20392 13716
rect 20260 13670 20312 13676
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20180 12850 20208 13126
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20272 11694 20300 13670
rect 20456 13462 20484 14010
rect 20548 13938 20576 14214
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 13530 20576 13874
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20626 13560 20682 13569
rect 20536 13524 20588 13530
rect 20626 13495 20682 13504
rect 20536 13466 20588 13472
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 12986 20392 13330
rect 20640 13002 20668 13495
rect 20732 13394 20760 13806
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20548 12974 20668 13002
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 11218 19932 11494
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19904 11098 19932 11154
rect 19904 11070 20024 11098
rect 19616 10908 19912 10928
rect 19672 10906 19696 10908
rect 19752 10906 19776 10908
rect 19832 10906 19856 10908
rect 19694 10854 19696 10906
rect 19758 10854 19770 10906
rect 19832 10854 19834 10906
rect 19672 10852 19696 10854
rect 19752 10852 19776 10854
rect 19832 10852 19856 10854
rect 19616 10832 19912 10852
rect 19996 10674 20024 11070
rect 20088 10810 20116 11630
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19444 10254 19564 10282
rect 20088 10266 20116 10542
rect 18972 10192 19024 10198
rect 18970 10160 18972 10169
rect 19432 10192 19484 10198
rect 19024 10160 19026 10169
rect 19432 10134 19484 10140
rect 18970 10095 19026 10104
rect 19444 9654 19472 10134
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19352 9110 19380 9318
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19246 8936 19302 8945
rect 19246 8871 19302 8880
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19168 7002 19196 8026
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19260 6730 19288 8871
rect 19338 8392 19394 8401
rect 19338 8327 19394 8336
rect 19352 8294 19380 8327
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19352 7886 19380 8026
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19444 7342 19472 9318
rect 19536 9217 19564 10254
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20180 10062 20208 10950
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 19616 9820 19912 9840
rect 19672 9818 19696 9820
rect 19752 9818 19776 9820
rect 19832 9818 19856 9820
rect 19694 9766 19696 9818
rect 19758 9766 19770 9818
rect 19832 9766 19834 9818
rect 19672 9764 19696 9766
rect 19752 9764 19776 9766
rect 19832 9764 19856 9766
rect 19616 9744 19912 9764
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19522 9208 19578 9217
rect 19812 9178 19840 9318
rect 19522 9143 19578 9152
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19536 8634 19564 8978
rect 19616 8968 19668 8974
rect 19614 8936 19616 8945
rect 19668 8936 19670 8945
rect 19614 8871 19670 8880
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19616 8732 19912 8752
rect 19672 8730 19696 8732
rect 19752 8730 19776 8732
rect 19832 8730 19856 8732
rect 19694 8678 19696 8730
rect 19758 8678 19770 8730
rect 19832 8678 19834 8730
rect 19672 8676 19696 8678
rect 19752 8676 19776 8678
rect 19832 8676 19856 8678
rect 19616 8656 19912 8676
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 7041 19380 7142
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19432 6928 19484 6934
rect 19430 6896 19432 6905
rect 19484 6896 19486 6905
rect 19430 6831 19486 6840
rect 19536 6798 19564 8570
rect 19800 8560 19852 8566
rect 19852 8520 19932 8548
rect 19800 8502 19852 8508
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19720 8294 19748 8434
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19708 8288 19760 8294
rect 19812 8265 19840 8298
rect 19904 8294 19932 8520
rect 19892 8288 19944 8294
rect 19708 8230 19760 8236
rect 19798 8256 19854 8265
rect 19892 8230 19944 8236
rect 19798 8191 19854 8200
rect 19996 7954 20024 8842
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19616 7644 19912 7664
rect 19672 7642 19696 7644
rect 19752 7642 19776 7644
rect 19832 7642 19856 7644
rect 19694 7590 19696 7642
rect 19758 7590 19770 7642
rect 19832 7590 19834 7642
rect 19672 7588 19696 7590
rect 19752 7588 19776 7590
rect 19832 7588 19856 7590
rect 19616 7568 19912 7588
rect 19616 7472 19668 7478
rect 19614 7440 19616 7449
rect 19668 7440 19670 7449
rect 20088 7426 20116 9930
rect 20180 9450 20208 9998
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 20272 9330 20300 11018
rect 19996 7410 20116 7426
rect 19614 7375 19670 7384
rect 19984 7404 20116 7410
rect 20036 7398 20116 7404
rect 20180 9302 20300 9330
rect 19984 7346 20036 7352
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19168 6322 19196 6598
rect 19444 6390 19472 6734
rect 19628 6644 19656 7278
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19996 6866 20024 7142
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19536 6616 19656 6644
rect 19432 6384 19484 6390
rect 19338 6352 19394 6361
rect 19156 6316 19208 6322
rect 19432 6326 19484 6332
rect 19338 6287 19340 6296
rect 19156 6258 19208 6264
rect 19392 6287 19394 6296
rect 19340 6258 19392 6264
rect 19536 6254 19564 6616
rect 19616 6556 19912 6576
rect 19672 6554 19696 6556
rect 19752 6554 19776 6556
rect 19832 6554 19856 6556
rect 19694 6502 19696 6554
rect 19758 6502 19770 6554
rect 19832 6502 19834 6554
rect 19672 6500 19696 6502
rect 19752 6500 19776 6502
rect 19832 6500 19856 6502
rect 19616 6480 19912 6500
rect 19798 6352 19854 6361
rect 19798 6287 19854 6296
rect 19812 6254 19840 6287
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19531 6248 19583 6254
rect 19531 6190 19583 6196
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19340 6112 19392 6118
rect 19338 6080 19340 6089
rect 19392 6080 19394 6089
rect 19338 6015 19394 6024
rect 19444 5953 19472 6190
rect 19430 5944 19486 5953
rect 19536 5914 19564 6190
rect 19430 5879 19486 5888
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19260 5030 19288 5510
rect 19432 5364 19484 5370
rect 19536 5352 19564 5714
rect 20180 5681 20208 9302
rect 20364 9194 20392 12922
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20456 12714 20484 12786
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20548 12322 20576 12974
rect 20824 12782 20852 13126
rect 20916 12986 20944 13262
rect 20904 12980 20956 12986
rect 21180 12980 21232 12986
rect 20904 12922 20956 12928
rect 21100 12940 21180 12968
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20456 11898 20484 12310
rect 20548 12294 20668 12322
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20548 11082 20576 12174
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20640 9994 20668 12294
rect 20916 12238 20944 12922
rect 20996 12708 21048 12714
rect 20996 12650 21048 12656
rect 21008 12374 21036 12650
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20732 11354 20760 11698
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20916 10130 20944 10542
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20732 9450 20760 10066
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9518 20852 9998
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20272 9166 20392 9194
rect 20272 7970 20300 9166
rect 20732 9042 20760 9386
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20364 8090 20392 8978
rect 20442 8936 20498 8945
rect 21100 8922 21128 12940
rect 21180 12922 21232 12928
rect 21914 12880 21970 12889
rect 21914 12815 21970 12824
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21836 12374 21864 12582
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21652 11286 21680 11562
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21376 10810 21404 11222
rect 21456 11212 21508 11218
rect 21456 11154 21508 11160
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21468 10606 21496 11154
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21652 10538 21680 11086
rect 21730 10976 21786 10985
rect 21730 10911 21786 10920
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21652 10266 21680 10474
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21180 10124 21232 10130
rect 21180 10066 21232 10072
rect 21192 9722 21220 10066
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21560 9450 21588 9862
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21100 8894 21220 8922
rect 20442 8871 20498 8880
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20272 7942 20392 7970
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20166 5672 20222 5681
rect 20166 5607 20222 5616
rect 19616 5468 19912 5488
rect 19672 5466 19696 5468
rect 19752 5466 19776 5468
rect 19832 5466 19856 5468
rect 19694 5414 19696 5466
rect 19758 5414 19770 5466
rect 19832 5414 19834 5466
rect 19672 5412 19696 5414
rect 19752 5412 19776 5414
rect 19832 5412 19856 5414
rect 19616 5392 19912 5412
rect 19484 5324 19564 5352
rect 19432 5306 19484 5312
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19260 4622 19288 4966
rect 19352 4758 19380 5170
rect 19524 5092 19576 5098
rect 19524 5034 19576 5040
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19168 3194 19196 4558
rect 19444 3738 19472 4626
rect 19536 4486 19564 5034
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19616 4380 19912 4400
rect 19672 4378 19696 4380
rect 19752 4378 19776 4380
rect 19832 4378 19856 4380
rect 19694 4326 19696 4378
rect 19758 4326 19770 4378
rect 19832 4326 19834 4378
rect 19672 4324 19696 4326
rect 19752 4324 19776 4326
rect 19832 4324 19856 4326
rect 19616 4304 19912 4324
rect 19996 4282 20024 4558
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19996 4078 20024 4218
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 15884 2748 16180 2768
rect 15940 2746 15964 2748
rect 16020 2746 16044 2748
rect 16100 2746 16124 2748
rect 15962 2694 15964 2746
rect 16026 2694 16038 2746
rect 16100 2694 16102 2746
rect 15940 2692 15964 2694
rect 16020 2692 16044 2694
rect 16100 2692 16124 2694
rect 15884 2672 16180 2692
rect 18064 2514 18092 2790
rect 19352 2582 19380 3402
rect 19536 2650 19564 3946
rect 19812 3738 19840 3946
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19616 3292 19912 3312
rect 19672 3290 19696 3292
rect 19752 3290 19776 3292
rect 19832 3290 19856 3292
rect 19694 3238 19696 3290
rect 19758 3238 19770 3290
rect 19832 3238 19834 3290
rect 19672 3236 19696 3238
rect 19752 3236 19776 3238
rect 19832 3236 19856 3238
rect 19616 3216 19912 3236
rect 20088 2650 20116 4966
rect 20180 4826 20208 4966
rect 20272 4826 20300 6734
rect 20364 6474 20392 7942
rect 20456 6780 20484 8871
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 20548 8498 21036 8514
rect 20536 8492 21036 8498
rect 20588 8486 21036 8492
rect 20536 8434 20588 8440
rect 21008 8430 21036 8486
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 20732 7818 20760 8366
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 7546 20760 7754
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20536 7336 20588 7342
rect 20588 7284 20760 7290
rect 20536 7278 20760 7284
rect 20548 7274 20760 7278
rect 20548 7268 20772 7274
rect 20548 7262 20720 7268
rect 20720 7210 20772 7216
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 6792 20588 6798
rect 20456 6752 20536 6780
rect 20456 6662 20484 6752
rect 20536 6734 20588 6740
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20364 6446 20484 6474
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20364 5914 20392 6190
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20180 3942 20208 4626
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 2990 20208 3878
rect 20272 3738 20300 4558
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20272 2922 20300 3674
rect 20364 3602 20392 5238
rect 20456 4321 20484 6446
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5953 20576 6258
rect 20534 5944 20590 5953
rect 20640 5914 20668 6802
rect 20732 6390 20760 7210
rect 20916 7002 20944 7822
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20916 6254 20944 6802
rect 21008 6662 21036 8366
rect 21100 8294 21128 8774
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7342 21128 7822
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20534 5879 20590 5888
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20732 5794 20760 6122
rect 20916 5914 20944 6190
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20640 5778 20760 5794
rect 20628 5772 20760 5778
rect 20680 5766 20760 5772
rect 20628 5714 20680 5720
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20442 4312 20498 4321
rect 20442 4247 20498 4256
rect 20548 3738 20576 5646
rect 21008 4758 21036 6054
rect 21100 5370 21128 6802
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 21192 5001 21220 8894
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21468 7546 21496 7890
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21744 7290 21772 10911
rect 21928 9178 21956 12815
rect 22020 11830 22048 13330
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21928 8616 21956 9114
rect 22008 8628 22060 8634
rect 21928 8588 22008 8616
rect 22008 8570 22060 8576
rect 21824 8288 21876 8294
rect 21822 8256 21824 8265
rect 21876 8256 21878 8265
rect 21822 8191 21878 8200
rect 21652 7262 21772 7290
rect 22112 7274 22140 19910
rect 22284 19858 22336 19864
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22296 19394 22324 19654
rect 22204 19366 22324 19394
rect 22204 17270 22232 19366
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22296 18970 22324 19178
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22388 18698 22416 19926
rect 22572 19802 22600 21286
rect 22834 20904 22890 20913
rect 22834 20839 22890 20848
rect 22744 20324 22796 20330
rect 22744 20266 22796 20272
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 19922 22692 20198
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22572 19774 22692 19802
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22480 18578 22508 18702
rect 22388 18550 22508 18578
rect 22388 18426 22416 18550
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22388 17202 22416 18362
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22480 17202 22508 18090
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22388 17082 22416 17138
rect 22388 17054 22600 17082
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16250 22416 16934
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22480 16114 22508 16730
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 13938 22232 15846
rect 22296 15162 22324 16050
rect 22572 15706 22600 17054
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 15586 22692 19774
rect 22756 19446 22784 20266
rect 22848 20058 22876 20839
rect 22940 20466 22968 23718
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 22834 19544 22890 19553
rect 22834 19479 22836 19488
rect 22888 19479 22890 19488
rect 22836 19450 22888 19456
rect 22744 19440 22796 19446
rect 22744 19382 22796 19388
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 17134 22784 18566
rect 22836 17536 22888 17542
rect 22836 17478 22888 17484
rect 22744 17128 22796 17134
rect 22744 17070 22796 17076
rect 22572 15558 22692 15586
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22388 14958 22416 15302
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22388 14770 22416 14894
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22296 13870 22324 14758
rect 22388 14742 22508 14770
rect 22480 13870 22508 14742
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22572 13530 22600 15558
rect 22848 14958 22876 17478
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22940 16114 22968 16390
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22940 15638 22968 16050
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22940 14482 22968 14758
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22664 13462 22692 14214
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22652 13456 22704 13462
rect 22652 13398 22704 13404
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12850 22508 13126
rect 22664 12850 22692 13398
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22756 12782 22784 13670
rect 22940 13326 22968 14418
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22664 11762 22692 12038
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22388 10810 22416 11698
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22388 10062 22416 10746
rect 22480 10130 22508 11290
rect 22664 11286 22692 11698
rect 22756 11694 22784 12582
rect 23032 12442 23060 19110
rect 23124 18329 23152 19654
rect 23110 18320 23166 18329
rect 23110 18255 23166 18264
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17678 23152 18158
rect 23112 17672 23164 17678
rect 23110 17640 23112 17649
rect 23164 17640 23166 17649
rect 23110 17575 23166 17584
rect 23110 16960 23166 16969
rect 23110 16895 23166 16904
rect 23124 16794 23152 16895
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23124 15570 23152 16730
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23124 13462 23152 13942
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23124 12646 23152 13398
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23216 12458 23244 20742
rect 23308 12986 23336 21422
rect 23492 20534 23520 23800
rect 23570 22264 23626 22273
rect 23570 22199 23626 22208
rect 23584 22098 23612 22199
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 24136 21962 24164 23800
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23400 19310 23428 19858
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23124 12430 23244 12458
rect 23018 12336 23074 12345
rect 22928 12300 22980 12306
rect 23018 12271 23074 12280
rect 22928 12242 22980 12248
rect 22940 11762 22968 12242
rect 22928 11756 22980 11762
rect 22928 11698 22980 11704
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22652 11280 22704 11286
rect 22652 11222 22704 11228
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 10266 22876 10406
rect 22926 10296 22982 10305
rect 22836 10260 22888 10266
rect 22926 10231 22982 10240
rect 22836 10202 22888 10208
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22940 9654 22968 10231
rect 22652 9648 22704 9654
rect 22928 9648 22980 9654
rect 22652 9590 22704 9596
rect 22742 9616 22798 9625
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22296 8498 22324 8774
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22284 8492 22336 8498
rect 22204 8452 22284 8480
rect 22100 7268 22152 7274
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21284 5914 21312 6598
rect 21652 6186 21680 7262
rect 22100 7210 22152 7216
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21916 6928 21968 6934
rect 21916 6870 21968 6876
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6254 21864 6734
rect 21928 6662 21956 6870
rect 22020 6866 22048 7142
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 22204 6798 22232 8452
rect 22284 8434 22336 8440
rect 22282 7440 22338 7449
rect 22282 7375 22284 7384
rect 22336 7375 22338 7384
rect 22284 7346 22336 7352
rect 22282 6896 22338 6905
rect 22388 6866 22416 8502
rect 22480 8498 22508 8978
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22480 8378 22508 8434
rect 22480 8350 22600 8378
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22480 8022 22508 8230
rect 22572 8090 22600 8350
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22282 6831 22338 6840
rect 22376 6860 22428 6866
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21468 5710 21496 5850
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5166 21404 5510
rect 21468 5302 21496 5646
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21178 4992 21234 5001
rect 21178 4927 21234 4936
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 21376 4690 21404 5102
rect 21652 4826 21680 6122
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21376 4146 21404 4626
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20916 4010 20944 4082
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20536 3732 20588 3738
rect 20536 3674 20588 3680
rect 20916 3602 20944 3946
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20916 2990 20944 3538
rect 21008 3194 21036 3538
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 20272 2446 20300 2858
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20732 2650 20760 2790
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20916 2514 20944 2926
rect 21008 2582 21036 3130
rect 20996 2576 21048 2582
rect 20996 2518 21048 2524
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 12152 2204 12448 2224
rect 12208 2202 12232 2204
rect 12288 2202 12312 2204
rect 12368 2202 12392 2204
rect 12230 2150 12232 2202
rect 12294 2150 12306 2202
rect 12368 2150 12370 2202
rect 12208 2148 12232 2150
rect 12288 2148 12312 2150
rect 12368 2148 12392 2150
rect 12152 2128 12448 2148
rect 19616 2204 19912 2224
rect 19672 2202 19696 2204
rect 19752 2202 19776 2204
rect 19832 2202 19856 2204
rect 19694 2150 19696 2202
rect 19758 2150 19770 2202
rect 19832 2150 19834 2202
rect 19672 2148 19696 2150
rect 19752 2148 19776 2150
rect 19832 2148 19856 2150
rect 19616 2128 19912 2148
rect 2042 0 2098 800
rect 6090 0 6146 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18418 0 18474 800
rect 21928 377 21956 6598
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 3670 22048 6054
rect 22112 5846 22140 6666
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 22204 5370 22232 6598
rect 22296 6254 22324 6831
rect 22376 6802 22428 6808
rect 22466 6352 22522 6361
rect 22466 6287 22468 6296
rect 22520 6287 22522 6296
rect 22468 6258 22520 6264
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22296 5370 22324 6190
rect 22572 5914 22600 7142
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22664 5794 22692 9590
rect 22742 9551 22798 9560
rect 22848 9608 22928 9636
rect 22756 6866 22784 9551
rect 22848 7342 22876 9608
rect 22928 9590 22980 9596
rect 23032 9586 23060 12271
rect 23124 9926 23152 12430
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23124 9761 23152 9862
rect 23110 9752 23166 9761
rect 23110 9687 23166 9696
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 22926 8256 22982 8265
rect 22926 8191 22982 8200
rect 22940 8022 22968 8191
rect 22928 8016 22980 8022
rect 22928 7958 22980 7964
rect 23032 7954 23060 9318
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23032 7585 23060 7890
rect 23018 7576 23074 7585
rect 23018 7511 23074 7520
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 23032 7041 23060 7511
rect 23018 7032 23074 7041
rect 23018 6967 23074 6976
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22572 5766 22692 5794
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22008 3664 22060 3670
rect 22008 3606 22060 3612
rect 22204 3398 22232 3674
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22020 2582 22048 3334
rect 22296 3194 22324 5102
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22388 3466 22416 4966
rect 22572 3641 22600 5766
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22558 3632 22614 3641
rect 22558 3567 22614 3576
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22664 2990 22692 5034
rect 22756 4758 22784 6802
rect 22928 6180 22980 6186
rect 22928 6122 22980 6128
rect 22940 5778 22968 6122
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5370 22968 5714
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22928 5092 22980 5098
rect 22928 5034 22980 5040
rect 22940 4826 22968 5034
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22744 4752 22796 4758
rect 22744 4694 22796 4700
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22848 4282 22876 4626
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22756 3602 22784 3946
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22664 2514 22692 2790
rect 22756 2650 22784 3538
rect 22848 2990 22876 4218
rect 23032 4146 23060 6967
rect 23216 6934 23244 12310
rect 23386 9752 23442 9761
rect 23386 9687 23442 9696
rect 23204 6928 23256 6934
rect 23204 6870 23256 6876
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22940 3058 22968 3470
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 23032 2854 23060 4082
rect 23400 2961 23428 9687
rect 23480 7268 23532 7274
rect 23480 7210 23532 7216
rect 23386 2952 23442 2961
rect 23386 2887 23442 2896
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22744 2644 22796 2650
rect 22744 2586 22796 2592
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22480 800 22508 2382
rect 23492 921 23520 7210
rect 23584 6089 23612 20198
rect 23676 9586 23704 20946
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23676 9110 23704 9386
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23570 6080 23626 6089
rect 23570 6015 23626 6024
rect 23584 2281 23612 6015
rect 23570 2272 23626 2281
rect 23570 2207 23626 2216
rect 23676 1601 23704 9046
rect 23662 1592 23718 1601
rect 23662 1527 23718 1536
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 21914 368 21970 377
rect 21914 303 21970 312
rect 22466 0 22522 800
<< via2 >>
rect 21822 24248 21878 24304
rect 2318 21548 2374 21584
rect 2318 21528 2320 21548
rect 2320 21528 2372 21548
rect 2372 21528 2374 21548
rect 4688 21786 4744 21788
rect 4768 21786 4824 21788
rect 4848 21786 4904 21788
rect 4928 21786 4984 21788
rect 4688 21734 4714 21786
rect 4714 21734 4744 21786
rect 4768 21734 4778 21786
rect 4778 21734 4824 21786
rect 4848 21734 4894 21786
rect 4894 21734 4904 21786
rect 4928 21734 4958 21786
rect 4958 21734 4984 21786
rect 4688 21732 4744 21734
rect 4768 21732 4824 21734
rect 4848 21732 4904 21734
rect 4928 21732 4984 21734
rect 1582 20460 1638 20496
rect 1582 20440 1584 20460
rect 1584 20440 1636 20460
rect 1636 20440 1638 20460
rect 2686 16496 2742 16552
rect 4688 20698 4744 20700
rect 4768 20698 4824 20700
rect 4848 20698 4904 20700
rect 4928 20698 4984 20700
rect 4688 20646 4714 20698
rect 4714 20646 4744 20698
rect 4768 20646 4778 20698
rect 4778 20646 4824 20698
rect 4848 20646 4894 20698
rect 4894 20646 4904 20698
rect 4928 20646 4958 20698
rect 4958 20646 4984 20698
rect 4688 20644 4744 20646
rect 4768 20644 4824 20646
rect 4848 20644 4904 20646
rect 4928 20644 4984 20646
rect 4618 20440 4674 20496
rect 4986 20440 5042 20496
rect 4688 19610 4744 19612
rect 4768 19610 4824 19612
rect 4848 19610 4904 19612
rect 4928 19610 4984 19612
rect 4688 19558 4714 19610
rect 4714 19558 4744 19610
rect 4768 19558 4778 19610
rect 4778 19558 4824 19610
rect 4848 19558 4894 19610
rect 4894 19558 4904 19610
rect 4928 19558 4958 19610
rect 4958 19558 4984 19610
rect 4688 19556 4744 19558
rect 4768 19556 4824 19558
rect 4848 19556 4904 19558
rect 4928 19556 4984 19558
rect 4688 18522 4744 18524
rect 4768 18522 4824 18524
rect 4848 18522 4904 18524
rect 4928 18522 4984 18524
rect 4688 18470 4714 18522
rect 4714 18470 4744 18522
rect 4768 18470 4778 18522
rect 4778 18470 4824 18522
rect 4848 18470 4894 18522
rect 4894 18470 4904 18522
rect 4928 18470 4958 18522
rect 4958 18470 4984 18522
rect 4688 18468 4744 18470
rect 4768 18468 4824 18470
rect 4848 18468 4904 18470
rect 4928 18468 4984 18470
rect 5998 20440 6054 20496
rect 4688 17434 4744 17436
rect 4768 17434 4824 17436
rect 4848 17434 4904 17436
rect 4928 17434 4984 17436
rect 4688 17382 4714 17434
rect 4714 17382 4744 17434
rect 4768 17382 4778 17434
rect 4778 17382 4824 17434
rect 4848 17382 4894 17434
rect 4894 17382 4904 17434
rect 4928 17382 4958 17434
rect 4958 17382 4984 17434
rect 4688 17380 4744 17382
rect 4768 17380 4824 17382
rect 4848 17380 4904 17382
rect 4928 17380 4984 17382
rect 2870 15272 2926 15328
rect 2686 13796 2742 13832
rect 2686 13776 2688 13796
rect 2688 13776 2740 13796
rect 2740 13776 2742 13796
rect 1398 9152 1454 9208
rect 4688 16346 4744 16348
rect 4768 16346 4824 16348
rect 4848 16346 4904 16348
rect 4928 16346 4984 16348
rect 4688 16294 4714 16346
rect 4714 16294 4744 16346
rect 4768 16294 4778 16346
rect 4778 16294 4824 16346
rect 4848 16294 4894 16346
rect 4894 16294 4904 16346
rect 4928 16294 4958 16346
rect 4958 16294 4984 16346
rect 4688 16292 4744 16294
rect 4768 16292 4824 16294
rect 4848 16292 4904 16294
rect 4928 16292 4984 16294
rect 4688 15258 4744 15260
rect 4768 15258 4824 15260
rect 4848 15258 4904 15260
rect 4928 15258 4984 15260
rect 4688 15206 4714 15258
rect 4714 15206 4744 15258
rect 4768 15206 4778 15258
rect 4778 15206 4824 15258
rect 4848 15206 4894 15258
rect 4894 15206 4904 15258
rect 4928 15206 4958 15258
rect 4958 15206 4984 15258
rect 4688 15204 4744 15206
rect 4768 15204 4824 15206
rect 4848 15204 4904 15206
rect 4928 15204 4984 15206
rect 6182 16516 6238 16552
rect 6182 16496 6184 16516
rect 6184 16496 6236 16516
rect 6236 16496 6238 16516
rect 4688 14170 4744 14172
rect 4768 14170 4824 14172
rect 4848 14170 4904 14172
rect 4928 14170 4984 14172
rect 4688 14118 4714 14170
rect 4714 14118 4744 14170
rect 4768 14118 4778 14170
rect 4778 14118 4824 14170
rect 4848 14118 4894 14170
rect 4894 14118 4904 14170
rect 4928 14118 4958 14170
rect 4958 14118 4984 14170
rect 4688 14116 4744 14118
rect 4768 14116 4824 14118
rect 4848 14116 4904 14118
rect 4928 14116 4984 14118
rect 8420 22330 8476 22332
rect 8500 22330 8556 22332
rect 8580 22330 8636 22332
rect 8660 22330 8716 22332
rect 8420 22278 8446 22330
rect 8446 22278 8476 22330
rect 8500 22278 8510 22330
rect 8510 22278 8556 22330
rect 8580 22278 8626 22330
rect 8626 22278 8636 22330
rect 8660 22278 8690 22330
rect 8690 22278 8716 22330
rect 8420 22276 8476 22278
rect 8500 22276 8556 22278
rect 8580 22276 8636 22278
rect 8660 22276 8716 22278
rect 8298 21528 8354 21584
rect 8022 19372 8078 19408
rect 8022 19352 8024 19372
rect 8024 19352 8076 19372
rect 8076 19352 8078 19372
rect 8420 21242 8476 21244
rect 8500 21242 8556 21244
rect 8580 21242 8636 21244
rect 8660 21242 8716 21244
rect 8420 21190 8446 21242
rect 8446 21190 8476 21242
rect 8500 21190 8510 21242
rect 8510 21190 8556 21242
rect 8580 21190 8626 21242
rect 8626 21190 8636 21242
rect 8660 21190 8690 21242
rect 8690 21190 8716 21242
rect 8420 21188 8476 21190
rect 8500 21188 8556 21190
rect 8580 21188 8636 21190
rect 8660 21188 8716 21190
rect 8420 20154 8476 20156
rect 8500 20154 8556 20156
rect 8580 20154 8636 20156
rect 8660 20154 8716 20156
rect 8420 20102 8446 20154
rect 8446 20102 8476 20154
rect 8500 20102 8510 20154
rect 8510 20102 8556 20154
rect 8580 20102 8626 20154
rect 8626 20102 8636 20154
rect 8660 20102 8690 20154
rect 8690 20102 8716 20154
rect 8420 20100 8476 20102
rect 8500 20100 8556 20102
rect 8580 20100 8636 20102
rect 8660 20100 8716 20102
rect 8420 19066 8476 19068
rect 8500 19066 8556 19068
rect 8580 19066 8636 19068
rect 8660 19066 8716 19068
rect 8420 19014 8446 19066
rect 8446 19014 8476 19066
rect 8500 19014 8510 19066
rect 8510 19014 8556 19066
rect 8580 19014 8626 19066
rect 8626 19014 8636 19066
rect 8660 19014 8690 19066
rect 8690 19014 8716 19066
rect 8420 19012 8476 19014
rect 8500 19012 8556 19014
rect 8580 19012 8636 19014
rect 8660 19012 8716 19014
rect 8420 17978 8476 17980
rect 8500 17978 8556 17980
rect 8580 17978 8636 17980
rect 8660 17978 8716 17980
rect 8420 17926 8446 17978
rect 8446 17926 8476 17978
rect 8500 17926 8510 17978
rect 8510 17926 8556 17978
rect 8580 17926 8626 17978
rect 8626 17926 8636 17978
rect 8660 17926 8690 17978
rect 8690 17926 8716 17978
rect 8420 17924 8476 17926
rect 8500 17924 8556 17926
rect 8580 17924 8636 17926
rect 8660 17924 8716 17926
rect 8420 16890 8476 16892
rect 8500 16890 8556 16892
rect 8580 16890 8636 16892
rect 8660 16890 8716 16892
rect 8420 16838 8446 16890
rect 8446 16838 8476 16890
rect 8500 16838 8510 16890
rect 8510 16838 8556 16890
rect 8580 16838 8626 16890
rect 8626 16838 8636 16890
rect 8660 16838 8690 16890
rect 8690 16838 8716 16890
rect 8420 16836 8476 16838
rect 8500 16836 8556 16838
rect 8580 16836 8636 16838
rect 8660 16836 8716 16838
rect 9126 19352 9182 19408
rect 8420 15802 8476 15804
rect 8500 15802 8556 15804
rect 8580 15802 8636 15804
rect 8660 15802 8716 15804
rect 8420 15750 8446 15802
rect 8446 15750 8476 15802
rect 8500 15750 8510 15802
rect 8510 15750 8556 15802
rect 8580 15750 8626 15802
rect 8626 15750 8636 15802
rect 8660 15750 8690 15802
rect 8690 15750 8716 15802
rect 8420 15748 8476 15750
rect 8500 15748 8556 15750
rect 8580 15748 8636 15750
rect 8660 15748 8716 15750
rect 10046 21428 10048 21448
rect 10048 21428 10100 21448
rect 10100 21428 10102 21448
rect 10046 21392 10102 21428
rect 11610 20984 11666 21040
rect 12152 21786 12208 21788
rect 12232 21786 12288 21788
rect 12312 21786 12368 21788
rect 12392 21786 12448 21788
rect 12152 21734 12178 21786
rect 12178 21734 12208 21786
rect 12232 21734 12242 21786
rect 12242 21734 12288 21786
rect 12312 21734 12358 21786
rect 12358 21734 12368 21786
rect 12392 21734 12422 21786
rect 12422 21734 12448 21786
rect 12152 21732 12208 21734
rect 12232 21732 12288 21734
rect 12312 21732 12368 21734
rect 12392 21732 12448 21734
rect 8420 14714 8476 14716
rect 8500 14714 8556 14716
rect 8580 14714 8636 14716
rect 8660 14714 8716 14716
rect 8420 14662 8446 14714
rect 8446 14662 8476 14714
rect 8500 14662 8510 14714
rect 8510 14662 8556 14714
rect 8580 14662 8626 14714
rect 8626 14662 8636 14714
rect 8660 14662 8690 14714
rect 8690 14662 8716 14714
rect 8420 14660 8476 14662
rect 8500 14660 8556 14662
rect 8580 14660 8636 14662
rect 8660 14660 8716 14662
rect 4688 13082 4744 13084
rect 4768 13082 4824 13084
rect 4848 13082 4904 13084
rect 4928 13082 4984 13084
rect 4688 13030 4714 13082
rect 4714 13030 4744 13082
rect 4768 13030 4778 13082
rect 4778 13030 4824 13082
rect 4848 13030 4894 13082
rect 4894 13030 4904 13082
rect 4928 13030 4958 13082
rect 4958 13030 4984 13082
rect 4688 13028 4744 13030
rect 4768 13028 4824 13030
rect 4848 13028 4904 13030
rect 4928 13028 4984 13030
rect 6274 13796 6330 13832
rect 6274 13776 6276 13796
rect 6276 13776 6328 13796
rect 6328 13776 6330 13796
rect 8420 13626 8476 13628
rect 8500 13626 8556 13628
rect 8580 13626 8636 13628
rect 8660 13626 8716 13628
rect 8420 13574 8446 13626
rect 8446 13574 8476 13626
rect 8500 13574 8510 13626
rect 8510 13574 8556 13626
rect 8580 13574 8626 13626
rect 8626 13574 8636 13626
rect 8660 13574 8690 13626
rect 8690 13574 8716 13626
rect 8420 13572 8476 13574
rect 8500 13572 8556 13574
rect 8580 13572 8636 13574
rect 8660 13572 8716 13574
rect 8420 12538 8476 12540
rect 8500 12538 8556 12540
rect 8580 12538 8636 12540
rect 8660 12538 8716 12540
rect 8420 12486 8446 12538
rect 8446 12486 8476 12538
rect 8500 12486 8510 12538
rect 8510 12486 8556 12538
rect 8580 12486 8626 12538
rect 8626 12486 8636 12538
rect 8660 12486 8690 12538
rect 8690 12486 8716 12538
rect 8420 12484 8476 12486
rect 8500 12484 8556 12486
rect 8580 12484 8636 12486
rect 8660 12484 8716 12486
rect 4688 11994 4744 11996
rect 4768 11994 4824 11996
rect 4848 11994 4904 11996
rect 4928 11994 4984 11996
rect 4688 11942 4714 11994
rect 4714 11942 4744 11994
rect 4768 11942 4778 11994
rect 4778 11942 4824 11994
rect 4848 11942 4894 11994
rect 4894 11942 4904 11994
rect 4928 11942 4958 11994
rect 4958 11942 4984 11994
rect 4688 11940 4744 11942
rect 4768 11940 4824 11942
rect 4848 11940 4904 11942
rect 4928 11940 4984 11942
rect 8420 11450 8476 11452
rect 8500 11450 8556 11452
rect 8580 11450 8636 11452
rect 8660 11450 8716 11452
rect 8420 11398 8446 11450
rect 8446 11398 8476 11450
rect 8500 11398 8510 11450
rect 8510 11398 8556 11450
rect 8580 11398 8626 11450
rect 8626 11398 8636 11450
rect 8660 11398 8690 11450
rect 8690 11398 8716 11450
rect 8420 11396 8476 11398
rect 8500 11396 8556 11398
rect 8580 11396 8636 11398
rect 8660 11396 8716 11398
rect 4688 10906 4744 10908
rect 4768 10906 4824 10908
rect 4848 10906 4904 10908
rect 4928 10906 4984 10908
rect 4688 10854 4714 10906
rect 4714 10854 4744 10906
rect 4768 10854 4778 10906
rect 4778 10854 4824 10906
rect 4848 10854 4894 10906
rect 4894 10854 4904 10906
rect 4928 10854 4958 10906
rect 4958 10854 4984 10906
rect 4688 10852 4744 10854
rect 4768 10852 4824 10854
rect 4848 10852 4904 10854
rect 4928 10852 4984 10854
rect 8420 10362 8476 10364
rect 8500 10362 8556 10364
rect 8580 10362 8636 10364
rect 8660 10362 8716 10364
rect 8420 10310 8446 10362
rect 8446 10310 8476 10362
rect 8500 10310 8510 10362
rect 8510 10310 8556 10362
rect 8580 10310 8626 10362
rect 8626 10310 8636 10362
rect 8660 10310 8690 10362
rect 8690 10310 8716 10362
rect 8420 10308 8476 10310
rect 8500 10308 8556 10310
rect 8580 10308 8636 10310
rect 8660 10308 8716 10310
rect 12152 20698 12208 20700
rect 12232 20698 12288 20700
rect 12312 20698 12368 20700
rect 12392 20698 12448 20700
rect 12152 20646 12178 20698
rect 12178 20646 12208 20698
rect 12232 20646 12242 20698
rect 12242 20646 12288 20698
rect 12312 20646 12358 20698
rect 12358 20646 12368 20698
rect 12392 20646 12422 20698
rect 12422 20646 12448 20698
rect 12152 20644 12208 20646
rect 12232 20644 12288 20646
rect 12312 20644 12368 20646
rect 12392 20644 12448 20646
rect 11886 19896 11942 19952
rect 11702 19236 11758 19272
rect 11702 19216 11704 19236
rect 11704 19216 11756 19236
rect 11756 19216 11758 19236
rect 12898 21528 12954 21584
rect 12530 19932 12532 19952
rect 12532 19932 12584 19952
rect 12584 19932 12586 19952
rect 12530 19896 12586 19932
rect 12152 19610 12208 19612
rect 12232 19610 12288 19612
rect 12312 19610 12368 19612
rect 12392 19610 12448 19612
rect 12152 19558 12178 19610
rect 12178 19558 12208 19610
rect 12232 19558 12242 19610
rect 12242 19558 12288 19610
rect 12312 19558 12358 19610
rect 12358 19558 12368 19610
rect 12392 19558 12422 19610
rect 12422 19558 12448 19610
rect 12152 19556 12208 19558
rect 12232 19556 12288 19558
rect 12312 19556 12368 19558
rect 12392 19556 12448 19558
rect 12438 19388 12440 19408
rect 12440 19388 12492 19408
rect 12492 19388 12494 19408
rect 12438 19352 12494 19388
rect 12152 18522 12208 18524
rect 12232 18522 12288 18524
rect 12312 18522 12368 18524
rect 12392 18522 12448 18524
rect 12152 18470 12178 18522
rect 12178 18470 12208 18522
rect 12232 18470 12242 18522
rect 12242 18470 12288 18522
rect 12312 18470 12358 18522
rect 12358 18470 12368 18522
rect 12392 18470 12422 18522
rect 12422 18470 12448 18522
rect 12152 18468 12208 18470
rect 12232 18468 12288 18470
rect 12312 18468 12368 18470
rect 12392 18468 12448 18470
rect 12438 17620 12440 17640
rect 12440 17620 12492 17640
rect 12492 17620 12494 17640
rect 12438 17584 12494 17620
rect 12152 17434 12208 17436
rect 12232 17434 12288 17436
rect 12312 17434 12368 17436
rect 12392 17434 12448 17436
rect 12152 17382 12178 17434
rect 12178 17382 12208 17434
rect 12232 17382 12242 17434
rect 12242 17382 12288 17434
rect 12312 17382 12358 17434
rect 12358 17382 12368 17434
rect 12392 17382 12422 17434
rect 12422 17382 12448 17434
rect 12152 17380 12208 17382
rect 12232 17380 12288 17382
rect 12312 17380 12368 17382
rect 12392 17380 12448 17382
rect 12152 16346 12208 16348
rect 12232 16346 12288 16348
rect 12312 16346 12368 16348
rect 12392 16346 12448 16348
rect 12152 16294 12178 16346
rect 12178 16294 12208 16346
rect 12232 16294 12242 16346
rect 12242 16294 12288 16346
rect 12312 16294 12358 16346
rect 12358 16294 12368 16346
rect 12392 16294 12422 16346
rect 12422 16294 12448 16346
rect 12152 16292 12208 16294
rect 12232 16292 12288 16294
rect 12312 16292 12368 16294
rect 12392 16292 12448 16294
rect 12152 15258 12208 15260
rect 12232 15258 12288 15260
rect 12312 15258 12368 15260
rect 12392 15258 12448 15260
rect 12152 15206 12178 15258
rect 12178 15206 12208 15258
rect 12232 15206 12242 15258
rect 12242 15206 12288 15258
rect 12312 15206 12358 15258
rect 12358 15206 12368 15258
rect 12392 15206 12422 15258
rect 12422 15206 12448 15258
rect 12152 15204 12208 15206
rect 12232 15204 12288 15206
rect 12312 15204 12368 15206
rect 12392 15204 12448 15206
rect 10506 13776 10562 13832
rect 4688 9818 4744 9820
rect 4768 9818 4824 9820
rect 4848 9818 4904 9820
rect 4928 9818 4984 9820
rect 4688 9766 4714 9818
rect 4714 9766 4744 9818
rect 4768 9766 4778 9818
rect 4778 9766 4824 9818
rect 4848 9766 4894 9818
rect 4894 9766 4904 9818
rect 4928 9766 4958 9818
rect 4958 9766 4984 9818
rect 4688 9764 4744 9766
rect 4768 9764 4824 9766
rect 4848 9764 4904 9766
rect 4928 9764 4984 9766
rect 8420 9274 8476 9276
rect 8500 9274 8556 9276
rect 8580 9274 8636 9276
rect 8660 9274 8716 9276
rect 8420 9222 8446 9274
rect 8446 9222 8476 9274
rect 8500 9222 8510 9274
rect 8510 9222 8556 9274
rect 8580 9222 8626 9274
rect 8626 9222 8636 9274
rect 8660 9222 8690 9274
rect 8690 9222 8716 9274
rect 8420 9220 8476 9222
rect 8500 9220 8556 9222
rect 8580 9220 8636 9222
rect 8660 9220 8716 9222
rect 12152 14170 12208 14172
rect 12232 14170 12288 14172
rect 12312 14170 12368 14172
rect 12392 14170 12448 14172
rect 12152 14118 12178 14170
rect 12178 14118 12208 14170
rect 12232 14118 12242 14170
rect 12242 14118 12288 14170
rect 12312 14118 12358 14170
rect 12358 14118 12368 14170
rect 12392 14118 12422 14170
rect 12422 14118 12448 14170
rect 12152 14116 12208 14118
rect 12232 14116 12288 14118
rect 12312 14116 12368 14118
rect 12392 14116 12448 14118
rect 13358 19760 13414 19816
rect 13910 19796 13912 19816
rect 13912 19796 13964 19816
rect 13964 19796 13966 19816
rect 13910 19760 13966 19796
rect 14922 20984 14978 21040
rect 14922 19488 14978 19544
rect 13358 17584 13414 17640
rect 14646 17620 14648 17640
rect 14648 17620 14700 17640
rect 14700 17620 14702 17640
rect 14646 17584 14702 17620
rect 12898 13796 12954 13832
rect 12898 13776 12900 13796
rect 12900 13776 12952 13796
rect 12952 13776 12954 13796
rect 12152 13082 12208 13084
rect 12232 13082 12288 13084
rect 12312 13082 12368 13084
rect 12392 13082 12448 13084
rect 12152 13030 12178 13082
rect 12178 13030 12208 13082
rect 12232 13030 12242 13082
rect 12242 13030 12288 13082
rect 12312 13030 12358 13082
rect 12358 13030 12368 13082
rect 12392 13030 12422 13082
rect 12422 13030 12448 13082
rect 12152 13028 12208 13030
rect 12232 13028 12288 13030
rect 12312 13028 12368 13030
rect 12392 13028 12448 13030
rect 12152 11994 12208 11996
rect 12232 11994 12288 11996
rect 12312 11994 12368 11996
rect 12392 11994 12448 11996
rect 12152 11942 12178 11994
rect 12178 11942 12208 11994
rect 12232 11942 12242 11994
rect 12242 11942 12288 11994
rect 12312 11942 12358 11994
rect 12358 11942 12368 11994
rect 12392 11942 12422 11994
rect 12422 11942 12448 11994
rect 12152 11940 12208 11942
rect 12232 11940 12288 11942
rect 12312 11940 12368 11942
rect 12392 11940 12448 11942
rect 15106 18672 15162 18728
rect 15884 22330 15940 22332
rect 15964 22330 16020 22332
rect 16044 22330 16100 22332
rect 16124 22330 16180 22332
rect 15884 22278 15910 22330
rect 15910 22278 15940 22330
rect 15964 22278 15974 22330
rect 15974 22278 16020 22330
rect 16044 22278 16090 22330
rect 16090 22278 16100 22330
rect 16124 22278 16154 22330
rect 16154 22278 16180 22330
rect 15884 22276 15940 22278
rect 15964 22276 16020 22278
rect 16044 22276 16100 22278
rect 16124 22276 16180 22278
rect 15750 21528 15806 21584
rect 15884 21242 15940 21244
rect 15964 21242 16020 21244
rect 16044 21242 16100 21244
rect 16124 21242 16180 21244
rect 15884 21190 15910 21242
rect 15910 21190 15940 21242
rect 15964 21190 15974 21242
rect 15974 21190 16020 21242
rect 16044 21190 16090 21242
rect 16090 21190 16100 21242
rect 16124 21190 16154 21242
rect 16154 21190 16180 21242
rect 15884 21188 15940 21190
rect 15964 21188 16020 21190
rect 16044 21188 16100 21190
rect 16124 21188 16180 21190
rect 15884 20154 15940 20156
rect 15964 20154 16020 20156
rect 16044 20154 16100 20156
rect 16124 20154 16180 20156
rect 15884 20102 15910 20154
rect 15910 20102 15940 20154
rect 15964 20102 15974 20154
rect 15974 20102 16020 20154
rect 16044 20102 16090 20154
rect 16090 20102 16100 20154
rect 16124 20102 16154 20154
rect 16154 20102 16180 20154
rect 15884 20100 15940 20102
rect 15964 20100 16020 20102
rect 16044 20100 16100 20102
rect 16124 20100 16180 20102
rect 16578 20032 16634 20088
rect 15658 18944 15714 19000
rect 15382 17584 15438 17640
rect 12152 10906 12208 10908
rect 12232 10906 12288 10908
rect 12312 10906 12368 10908
rect 12392 10906 12448 10908
rect 12152 10854 12178 10906
rect 12178 10854 12208 10906
rect 12232 10854 12242 10906
rect 12242 10854 12288 10906
rect 12312 10854 12358 10906
rect 12358 10854 12368 10906
rect 12392 10854 12422 10906
rect 12422 10854 12448 10906
rect 12152 10852 12208 10854
rect 12232 10852 12288 10854
rect 12312 10852 12368 10854
rect 12392 10852 12448 10854
rect 4688 8730 4744 8732
rect 4768 8730 4824 8732
rect 4848 8730 4904 8732
rect 4928 8730 4984 8732
rect 4688 8678 4714 8730
rect 4714 8678 4744 8730
rect 4768 8678 4778 8730
rect 4778 8678 4824 8730
rect 4848 8678 4894 8730
rect 4894 8678 4904 8730
rect 4928 8678 4958 8730
rect 4958 8678 4984 8730
rect 4688 8676 4744 8678
rect 4768 8676 4824 8678
rect 4848 8676 4904 8678
rect 4928 8676 4984 8678
rect 8420 8186 8476 8188
rect 8500 8186 8556 8188
rect 8580 8186 8636 8188
rect 8660 8186 8716 8188
rect 8420 8134 8446 8186
rect 8446 8134 8476 8186
rect 8500 8134 8510 8186
rect 8510 8134 8556 8186
rect 8580 8134 8626 8186
rect 8626 8134 8636 8186
rect 8660 8134 8690 8186
rect 8690 8134 8716 8186
rect 8420 8132 8476 8134
rect 8500 8132 8556 8134
rect 8580 8132 8636 8134
rect 8660 8132 8716 8134
rect 4688 7642 4744 7644
rect 4768 7642 4824 7644
rect 4848 7642 4904 7644
rect 4928 7642 4984 7644
rect 4688 7590 4714 7642
rect 4714 7590 4744 7642
rect 4768 7590 4778 7642
rect 4778 7590 4824 7642
rect 4848 7590 4894 7642
rect 4894 7590 4904 7642
rect 4928 7590 4958 7642
rect 4958 7590 4984 7642
rect 4688 7588 4744 7590
rect 4768 7588 4824 7590
rect 4848 7588 4904 7590
rect 4928 7588 4984 7590
rect 12152 9818 12208 9820
rect 12232 9818 12288 9820
rect 12312 9818 12368 9820
rect 12392 9818 12448 9820
rect 12152 9766 12178 9818
rect 12178 9766 12208 9818
rect 12232 9766 12242 9818
rect 12242 9766 12288 9818
rect 12312 9766 12358 9818
rect 12358 9766 12368 9818
rect 12392 9766 12422 9818
rect 12422 9766 12448 9818
rect 12152 9764 12208 9766
rect 12232 9764 12288 9766
rect 12312 9764 12368 9766
rect 12392 9764 12448 9766
rect 11702 8472 11758 8528
rect 12152 8730 12208 8732
rect 12232 8730 12288 8732
rect 12312 8730 12368 8732
rect 12392 8730 12448 8732
rect 12152 8678 12178 8730
rect 12178 8678 12208 8730
rect 12232 8678 12242 8730
rect 12242 8678 12288 8730
rect 12312 8678 12358 8730
rect 12358 8678 12368 8730
rect 12392 8678 12422 8730
rect 12422 8678 12448 8730
rect 12152 8676 12208 8678
rect 12232 8676 12288 8678
rect 12312 8676 12368 8678
rect 12392 8676 12448 8678
rect 8420 7098 8476 7100
rect 8500 7098 8556 7100
rect 8580 7098 8636 7100
rect 8660 7098 8716 7100
rect 8420 7046 8446 7098
rect 8446 7046 8476 7098
rect 8500 7046 8510 7098
rect 8510 7046 8556 7098
rect 8580 7046 8626 7098
rect 8626 7046 8636 7098
rect 8660 7046 8690 7098
rect 8690 7046 8716 7098
rect 8420 7044 8476 7046
rect 8500 7044 8556 7046
rect 8580 7044 8636 7046
rect 8660 7044 8716 7046
rect 12162 8492 12218 8528
rect 12162 8472 12164 8492
rect 12164 8472 12216 8492
rect 12216 8472 12218 8492
rect 15884 19066 15940 19068
rect 15964 19066 16020 19068
rect 16044 19066 16100 19068
rect 16124 19066 16180 19068
rect 15884 19014 15910 19066
rect 15910 19014 15940 19066
rect 15964 19014 15974 19066
rect 15974 19014 16020 19066
rect 16044 19014 16090 19066
rect 16090 19014 16100 19066
rect 16124 19014 16154 19066
rect 16154 19014 16180 19066
rect 15884 19012 15940 19014
rect 15964 19012 16020 19014
rect 16044 19012 16100 19014
rect 16124 19012 16180 19014
rect 15884 17978 15940 17980
rect 15964 17978 16020 17980
rect 16044 17978 16100 17980
rect 16124 17978 16180 17980
rect 15884 17926 15910 17978
rect 15910 17926 15940 17978
rect 15964 17926 15974 17978
rect 15974 17926 16020 17978
rect 16044 17926 16090 17978
rect 16090 17926 16100 17978
rect 16124 17926 16154 17978
rect 16154 17926 16180 17978
rect 15884 17924 15940 17926
rect 15964 17924 16020 17926
rect 16044 17924 16100 17926
rect 16124 17924 16180 17926
rect 15884 16890 15940 16892
rect 15964 16890 16020 16892
rect 16044 16890 16100 16892
rect 16124 16890 16180 16892
rect 15884 16838 15910 16890
rect 15910 16838 15940 16890
rect 15964 16838 15974 16890
rect 15974 16838 16020 16890
rect 16044 16838 16090 16890
rect 16090 16838 16100 16890
rect 16124 16838 16154 16890
rect 16154 16838 16180 16890
rect 15884 16836 15940 16838
rect 15964 16836 16020 16838
rect 16044 16836 16100 16838
rect 16124 16836 16180 16838
rect 17406 21392 17462 21448
rect 17498 20032 17554 20088
rect 16302 18808 16358 18864
rect 16946 19216 17002 19272
rect 16854 18708 16856 18728
rect 16856 18708 16908 18728
rect 16908 18708 16910 18728
rect 16854 18672 16910 18708
rect 15884 15802 15940 15804
rect 15964 15802 16020 15804
rect 16044 15802 16100 15804
rect 16124 15802 16180 15804
rect 15884 15750 15910 15802
rect 15910 15750 15940 15802
rect 15964 15750 15974 15802
rect 15974 15750 16020 15802
rect 16044 15750 16090 15802
rect 16090 15750 16100 15802
rect 16124 15750 16154 15802
rect 16154 15750 16180 15802
rect 15884 15748 15940 15750
rect 15964 15748 16020 15750
rect 16044 15748 16100 15750
rect 16124 15748 16180 15750
rect 15884 14714 15940 14716
rect 15964 14714 16020 14716
rect 16044 14714 16100 14716
rect 16124 14714 16180 14716
rect 15884 14662 15910 14714
rect 15910 14662 15940 14714
rect 15964 14662 15974 14714
rect 15974 14662 16020 14714
rect 16044 14662 16090 14714
rect 16090 14662 16100 14714
rect 16124 14662 16154 14714
rect 16154 14662 16180 14714
rect 15884 14660 15940 14662
rect 15964 14660 16020 14662
rect 16044 14660 16100 14662
rect 16124 14660 16180 14662
rect 15884 13626 15940 13628
rect 15964 13626 16020 13628
rect 16044 13626 16100 13628
rect 16124 13626 16180 13628
rect 15884 13574 15910 13626
rect 15910 13574 15940 13626
rect 15964 13574 15974 13626
rect 15974 13574 16020 13626
rect 16044 13574 16090 13626
rect 16090 13574 16100 13626
rect 16124 13574 16154 13626
rect 16154 13574 16180 13626
rect 15884 13572 15940 13574
rect 15964 13572 16020 13574
rect 16044 13572 16100 13574
rect 16124 13572 16180 13574
rect 15014 10104 15070 10160
rect 15884 12538 15940 12540
rect 15964 12538 16020 12540
rect 16044 12538 16100 12540
rect 16124 12538 16180 12540
rect 15884 12486 15910 12538
rect 15910 12486 15940 12538
rect 15964 12486 15974 12538
rect 15974 12486 16020 12538
rect 16044 12486 16090 12538
rect 16090 12486 16100 12538
rect 16124 12486 16154 12538
rect 16154 12486 16180 12538
rect 15884 12484 15940 12486
rect 15964 12484 16020 12486
rect 16044 12484 16100 12486
rect 16124 12484 16180 12486
rect 15884 11450 15940 11452
rect 15964 11450 16020 11452
rect 16044 11450 16100 11452
rect 16124 11450 16180 11452
rect 15884 11398 15910 11450
rect 15910 11398 15940 11450
rect 15964 11398 15974 11450
rect 15974 11398 16020 11450
rect 16044 11398 16090 11450
rect 16090 11398 16100 11450
rect 16124 11398 16154 11450
rect 16154 11398 16180 11450
rect 15884 11396 15940 11398
rect 15964 11396 16020 11398
rect 16044 11396 16100 11398
rect 16124 11396 16180 11398
rect 15884 10362 15940 10364
rect 15964 10362 16020 10364
rect 16044 10362 16100 10364
rect 16124 10362 16180 10364
rect 15884 10310 15910 10362
rect 15910 10310 15940 10362
rect 15964 10310 15974 10362
rect 15974 10310 16020 10362
rect 16044 10310 16090 10362
rect 16090 10310 16100 10362
rect 16124 10310 16154 10362
rect 16154 10310 16180 10362
rect 15884 10308 15940 10310
rect 15964 10308 16020 10310
rect 16044 10308 16100 10310
rect 16124 10308 16180 10310
rect 14922 9036 14978 9072
rect 14922 9016 14924 9036
rect 14924 9016 14976 9036
rect 14976 9016 14978 9036
rect 15106 8880 15162 8936
rect 4688 6554 4744 6556
rect 4768 6554 4824 6556
rect 4848 6554 4904 6556
rect 4928 6554 4984 6556
rect 4688 6502 4714 6554
rect 4714 6502 4744 6554
rect 4768 6502 4778 6554
rect 4778 6502 4824 6554
rect 4848 6502 4894 6554
rect 4894 6502 4904 6554
rect 4928 6502 4958 6554
rect 4958 6502 4984 6554
rect 4688 6500 4744 6502
rect 4768 6500 4824 6502
rect 4848 6500 4904 6502
rect 4928 6500 4984 6502
rect 8420 6010 8476 6012
rect 8500 6010 8556 6012
rect 8580 6010 8636 6012
rect 8660 6010 8716 6012
rect 8420 5958 8446 6010
rect 8446 5958 8476 6010
rect 8500 5958 8510 6010
rect 8510 5958 8556 6010
rect 8580 5958 8626 6010
rect 8626 5958 8636 6010
rect 8660 5958 8690 6010
rect 8690 5958 8716 6010
rect 8420 5956 8476 5958
rect 8500 5956 8556 5958
rect 8580 5956 8636 5958
rect 8660 5956 8716 5958
rect 4688 5466 4744 5468
rect 4768 5466 4824 5468
rect 4848 5466 4904 5468
rect 4928 5466 4984 5468
rect 4688 5414 4714 5466
rect 4714 5414 4744 5466
rect 4768 5414 4778 5466
rect 4778 5414 4824 5466
rect 4848 5414 4894 5466
rect 4894 5414 4904 5466
rect 4928 5414 4958 5466
rect 4958 5414 4984 5466
rect 4688 5412 4744 5414
rect 4768 5412 4824 5414
rect 4848 5412 4904 5414
rect 4928 5412 4984 5414
rect 8420 4922 8476 4924
rect 8500 4922 8556 4924
rect 8580 4922 8636 4924
rect 8660 4922 8716 4924
rect 8420 4870 8446 4922
rect 8446 4870 8476 4922
rect 8500 4870 8510 4922
rect 8510 4870 8556 4922
rect 8580 4870 8626 4922
rect 8626 4870 8636 4922
rect 8660 4870 8690 4922
rect 8690 4870 8716 4922
rect 8420 4868 8476 4870
rect 8500 4868 8556 4870
rect 8580 4868 8636 4870
rect 8660 4868 8716 4870
rect 12152 7642 12208 7644
rect 12232 7642 12288 7644
rect 12312 7642 12368 7644
rect 12392 7642 12448 7644
rect 12152 7590 12178 7642
rect 12178 7590 12208 7642
rect 12232 7590 12242 7642
rect 12242 7590 12288 7642
rect 12312 7590 12358 7642
rect 12358 7590 12368 7642
rect 12392 7590 12422 7642
rect 12422 7590 12448 7642
rect 12152 7588 12208 7590
rect 12232 7588 12288 7590
rect 12312 7588 12368 7590
rect 12392 7588 12448 7590
rect 12152 6554 12208 6556
rect 12232 6554 12288 6556
rect 12312 6554 12368 6556
rect 12392 6554 12448 6556
rect 12152 6502 12178 6554
rect 12178 6502 12208 6554
rect 12232 6502 12242 6554
rect 12242 6502 12288 6554
rect 12312 6502 12358 6554
rect 12358 6502 12368 6554
rect 12392 6502 12422 6554
rect 12422 6502 12448 6554
rect 12152 6500 12208 6502
rect 12232 6500 12288 6502
rect 12312 6500 12368 6502
rect 12392 6500 12448 6502
rect 12152 5466 12208 5468
rect 12232 5466 12288 5468
rect 12312 5466 12368 5468
rect 12392 5466 12448 5468
rect 12152 5414 12178 5466
rect 12178 5414 12208 5466
rect 12232 5414 12242 5466
rect 12242 5414 12288 5466
rect 12312 5414 12358 5466
rect 12358 5414 12368 5466
rect 12392 5414 12422 5466
rect 12422 5414 12448 5466
rect 12152 5412 12208 5414
rect 12232 5412 12288 5414
rect 12312 5412 12368 5414
rect 12392 5412 12448 5414
rect 14922 8064 14978 8120
rect 14738 7928 14794 7984
rect 15884 9274 15940 9276
rect 15964 9274 16020 9276
rect 16044 9274 16100 9276
rect 16124 9274 16180 9276
rect 15884 9222 15910 9274
rect 15910 9222 15940 9274
rect 15964 9222 15974 9274
rect 15974 9222 16020 9274
rect 16044 9222 16090 9274
rect 16090 9222 16100 9274
rect 16124 9222 16154 9274
rect 16154 9222 16180 9274
rect 15884 9220 15940 9222
rect 15964 9220 16020 9222
rect 16044 9220 16100 9222
rect 16124 9220 16180 9222
rect 15658 9016 15714 9072
rect 15750 8472 15806 8528
rect 15884 8186 15940 8188
rect 15964 8186 16020 8188
rect 16044 8186 16100 8188
rect 16124 8186 16180 8188
rect 15884 8134 15910 8186
rect 15910 8134 15940 8186
rect 15964 8134 15974 8186
rect 15974 8134 16020 8186
rect 16044 8134 16090 8186
rect 16090 8134 16100 8186
rect 16124 8134 16154 8186
rect 16154 8134 16180 8186
rect 15884 8132 15940 8134
rect 15964 8132 16020 8134
rect 16044 8132 16100 8134
rect 16124 8132 16180 8134
rect 15566 8064 15622 8120
rect 16026 7948 16082 7984
rect 16026 7928 16028 7948
rect 16028 7928 16080 7948
rect 16080 7928 16082 7948
rect 15884 7098 15940 7100
rect 15964 7098 16020 7100
rect 16044 7098 16100 7100
rect 16124 7098 16180 7100
rect 15884 7046 15910 7098
rect 15910 7046 15940 7098
rect 15964 7046 15974 7098
rect 15974 7046 16020 7098
rect 16044 7046 16090 7098
rect 16090 7046 16100 7098
rect 16124 7046 16154 7098
rect 16154 7046 16180 7098
rect 15884 7044 15940 7046
rect 15964 7044 16020 7046
rect 16044 7044 16100 7046
rect 16124 7044 16180 7046
rect 15884 6010 15940 6012
rect 15964 6010 16020 6012
rect 16044 6010 16100 6012
rect 16124 6010 16180 6012
rect 15884 5958 15910 6010
rect 15910 5958 15940 6010
rect 15964 5958 15974 6010
rect 15974 5958 16020 6010
rect 16044 5958 16090 6010
rect 16090 5958 16100 6010
rect 16124 5958 16154 6010
rect 16154 5958 16180 6010
rect 15884 5956 15940 5958
rect 15964 5956 16020 5958
rect 16044 5956 16100 5958
rect 16124 5956 16180 5958
rect 16486 8916 16488 8936
rect 16488 8916 16540 8936
rect 16540 8916 16542 8936
rect 16486 8880 16542 8916
rect 17406 7928 17462 7984
rect 19154 19508 19210 19544
rect 19154 19488 19156 19508
rect 19156 19488 19208 19508
rect 19208 19488 19210 19508
rect 18418 10104 18474 10160
rect 19616 21786 19672 21788
rect 19696 21786 19752 21788
rect 19776 21786 19832 21788
rect 19856 21786 19912 21788
rect 19616 21734 19642 21786
rect 19642 21734 19672 21786
rect 19696 21734 19706 21786
rect 19706 21734 19752 21786
rect 19776 21734 19822 21786
rect 19822 21734 19832 21786
rect 19856 21734 19886 21786
rect 19886 21734 19912 21786
rect 19616 21732 19672 21734
rect 19696 21732 19752 21734
rect 19776 21732 19832 21734
rect 19856 21732 19912 21734
rect 19616 20698 19672 20700
rect 19696 20698 19752 20700
rect 19776 20698 19832 20700
rect 19856 20698 19912 20700
rect 19616 20646 19642 20698
rect 19642 20646 19672 20698
rect 19696 20646 19706 20698
rect 19706 20646 19752 20698
rect 19776 20646 19822 20698
rect 19822 20646 19832 20698
rect 19856 20646 19886 20698
rect 19886 20646 19912 20698
rect 19616 20644 19672 20646
rect 19696 20644 19752 20646
rect 19776 20644 19832 20646
rect 19856 20644 19912 20646
rect 19338 19352 19394 19408
rect 19616 19610 19672 19612
rect 19696 19610 19752 19612
rect 19776 19610 19832 19612
rect 19856 19610 19912 19612
rect 19616 19558 19642 19610
rect 19642 19558 19672 19610
rect 19696 19558 19706 19610
rect 19706 19558 19752 19610
rect 19776 19558 19822 19610
rect 19822 19558 19832 19610
rect 19856 19558 19886 19610
rect 19886 19558 19912 19610
rect 19616 19556 19672 19558
rect 19696 19556 19752 19558
rect 19776 19556 19832 19558
rect 19856 19556 19912 19558
rect 21914 23568 21970 23624
rect 22006 22888 22062 22944
rect 22466 21528 22522 21584
rect 22466 20168 22522 20224
rect 19616 18522 19672 18524
rect 19696 18522 19752 18524
rect 19776 18522 19832 18524
rect 19856 18522 19912 18524
rect 19616 18470 19642 18522
rect 19642 18470 19672 18522
rect 19696 18470 19706 18522
rect 19706 18470 19752 18522
rect 19776 18470 19822 18522
rect 19822 18470 19832 18522
rect 19856 18470 19886 18522
rect 19886 18470 19912 18522
rect 19616 18468 19672 18470
rect 19696 18468 19752 18470
rect 19776 18468 19832 18470
rect 19856 18468 19912 18470
rect 21178 18808 21234 18864
rect 19616 17434 19672 17436
rect 19696 17434 19752 17436
rect 19776 17434 19832 17436
rect 19856 17434 19912 17436
rect 19616 17382 19642 17434
rect 19642 17382 19672 17434
rect 19696 17382 19706 17434
rect 19706 17382 19752 17434
rect 19776 17382 19822 17434
rect 19822 17382 19832 17434
rect 19856 17382 19886 17434
rect 19886 17382 19912 17434
rect 19616 17380 19672 17382
rect 19696 17380 19752 17382
rect 19776 17380 19832 17382
rect 19856 17380 19912 17382
rect 19616 16346 19672 16348
rect 19696 16346 19752 16348
rect 19776 16346 19832 16348
rect 19856 16346 19912 16348
rect 19616 16294 19642 16346
rect 19642 16294 19672 16346
rect 19696 16294 19706 16346
rect 19706 16294 19752 16346
rect 19776 16294 19822 16346
rect 19822 16294 19832 16346
rect 19856 16294 19886 16346
rect 19886 16294 19912 16346
rect 19616 16292 19672 16294
rect 19696 16292 19752 16294
rect 19776 16292 19832 16294
rect 19856 16292 19912 16294
rect 20258 16224 20314 16280
rect 19338 15544 19394 15600
rect 19616 15258 19672 15260
rect 19696 15258 19752 15260
rect 19776 15258 19832 15260
rect 19856 15258 19912 15260
rect 19616 15206 19642 15258
rect 19642 15206 19672 15258
rect 19696 15206 19706 15258
rect 19706 15206 19752 15258
rect 19776 15206 19822 15258
rect 19822 15206 19832 15258
rect 19856 15206 19886 15258
rect 19886 15206 19912 15258
rect 19616 15204 19672 15206
rect 19696 15204 19752 15206
rect 19776 15204 19832 15206
rect 19856 15204 19912 15206
rect 19338 14864 19394 14920
rect 19338 14320 19394 14376
rect 19616 14170 19672 14172
rect 19696 14170 19752 14172
rect 19776 14170 19832 14172
rect 19856 14170 19912 14172
rect 19616 14118 19642 14170
rect 19642 14118 19672 14170
rect 19696 14118 19706 14170
rect 19706 14118 19752 14170
rect 19776 14118 19822 14170
rect 19822 14118 19832 14170
rect 19856 14118 19886 14170
rect 19886 14118 19912 14170
rect 19616 14116 19672 14118
rect 19696 14116 19752 14118
rect 19776 14116 19832 14118
rect 19856 14116 19912 14118
rect 15884 4922 15940 4924
rect 15964 4922 16020 4924
rect 16044 4922 16100 4924
rect 16124 4922 16180 4924
rect 15884 4870 15910 4922
rect 15910 4870 15940 4922
rect 15964 4870 15974 4922
rect 15974 4870 16020 4922
rect 16044 4870 16090 4922
rect 16090 4870 16100 4922
rect 16124 4870 16154 4922
rect 16154 4870 16180 4922
rect 15884 4868 15940 4870
rect 15964 4868 16020 4870
rect 16044 4868 16100 4870
rect 16124 4868 16180 4870
rect 4688 4378 4744 4380
rect 4768 4378 4824 4380
rect 4848 4378 4904 4380
rect 4928 4378 4984 4380
rect 4688 4326 4714 4378
rect 4714 4326 4744 4378
rect 4768 4326 4778 4378
rect 4778 4326 4824 4378
rect 4848 4326 4894 4378
rect 4894 4326 4904 4378
rect 4928 4326 4958 4378
rect 4958 4326 4984 4378
rect 4688 4324 4744 4326
rect 4768 4324 4824 4326
rect 4848 4324 4904 4326
rect 4928 4324 4984 4326
rect 12152 4378 12208 4380
rect 12232 4378 12288 4380
rect 12312 4378 12368 4380
rect 12392 4378 12448 4380
rect 12152 4326 12178 4378
rect 12178 4326 12208 4378
rect 12232 4326 12242 4378
rect 12242 4326 12288 4378
rect 12312 4326 12358 4378
rect 12358 4326 12368 4378
rect 12392 4326 12422 4378
rect 12422 4326 12448 4378
rect 12152 4324 12208 4326
rect 12232 4324 12288 4326
rect 12312 4324 12368 4326
rect 12392 4324 12448 4326
rect 8420 3834 8476 3836
rect 8500 3834 8556 3836
rect 8580 3834 8636 3836
rect 8660 3834 8716 3836
rect 8420 3782 8446 3834
rect 8446 3782 8476 3834
rect 8500 3782 8510 3834
rect 8510 3782 8556 3834
rect 8580 3782 8626 3834
rect 8626 3782 8636 3834
rect 8660 3782 8690 3834
rect 8690 3782 8716 3834
rect 8420 3780 8476 3782
rect 8500 3780 8556 3782
rect 8580 3780 8636 3782
rect 8660 3780 8716 3782
rect 15884 3834 15940 3836
rect 15964 3834 16020 3836
rect 16044 3834 16100 3836
rect 16124 3834 16180 3836
rect 15884 3782 15910 3834
rect 15910 3782 15940 3834
rect 15964 3782 15974 3834
rect 15974 3782 16020 3834
rect 16044 3782 16090 3834
rect 16090 3782 16100 3834
rect 16124 3782 16154 3834
rect 16154 3782 16180 3834
rect 15884 3780 15940 3782
rect 15964 3780 16020 3782
rect 16044 3780 16100 3782
rect 16124 3780 16180 3782
rect 4688 3290 4744 3292
rect 4768 3290 4824 3292
rect 4848 3290 4904 3292
rect 4928 3290 4984 3292
rect 4688 3238 4714 3290
rect 4714 3238 4744 3290
rect 4768 3238 4778 3290
rect 4778 3238 4824 3290
rect 4848 3238 4894 3290
rect 4894 3238 4904 3290
rect 4928 3238 4958 3290
rect 4958 3238 4984 3290
rect 4688 3236 4744 3238
rect 4768 3236 4824 3238
rect 4848 3236 4904 3238
rect 4928 3236 4984 3238
rect 12152 3290 12208 3292
rect 12232 3290 12288 3292
rect 12312 3290 12368 3292
rect 12392 3290 12448 3292
rect 12152 3238 12178 3290
rect 12178 3238 12208 3290
rect 12232 3238 12242 3290
rect 12242 3238 12288 3290
rect 12312 3238 12358 3290
rect 12358 3238 12368 3290
rect 12392 3238 12422 3290
rect 12422 3238 12448 3290
rect 12152 3236 12208 3238
rect 12232 3236 12288 3238
rect 12312 3236 12368 3238
rect 12392 3236 12448 3238
rect 1950 3052 2006 3088
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 4688 2202 4744 2204
rect 4768 2202 4824 2204
rect 4848 2202 4904 2204
rect 4928 2202 4984 2204
rect 4688 2150 4714 2202
rect 4714 2150 4744 2202
rect 4768 2150 4778 2202
rect 4778 2150 4824 2202
rect 4848 2150 4894 2202
rect 4894 2150 4904 2202
rect 4928 2150 4958 2202
rect 4958 2150 4984 2202
rect 4688 2148 4744 2150
rect 4768 2148 4824 2150
rect 4848 2148 4904 2150
rect 4928 2148 4984 2150
rect 8420 2746 8476 2748
rect 8500 2746 8556 2748
rect 8580 2746 8636 2748
rect 8660 2746 8716 2748
rect 8420 2694 8446 2746
rect 8446 2694 8476 2746
rect 8500 2694 8510 2746
rect 8510 2694 8556 2746
rect 8580 2694 8626 2746
rect 8626 2694 8636 2746
rect 8660 2694 8690 2746
rect 8690 2694 8716 2746
rect 8420 2692 8476 2694
rect 8500 2692 8556 2694
rect 8580 2692 8636 2694
rect 8660 2692 8716 2694
rect 19616 13082 19672 13084
rect 19696 13082 19752 13084
rect 19776 13082 19832 13084
rect 19856 13082 19912 13084
rect 19616 13030 19642 13082
rect 19642 13030 19672 13082
rect 19696 13030 19706 13082
rect 19706 13030 19752 13082
rect 19776 13030 19822 13082
rect 19822 13030 19832 13082
rect 19856 13030 19886 13082
rect 19886 13030 19912 13082
rect 19616 13028 19672 13030
rect 19696 13028 19752 13030
rect 19776 13028 19832 13030
rect 19856 13028 19912 13030
rect 19430 11600 19486 11656
rect 19616 11994 19672 11996
rect 19696 11994 19752 11996
rect 19776 11994 19832 11996
rect 19856 11994 19912 11996
rect 19616 11942 19642 11994
rect 19642 11942 19672 11994
rect 19696 11942 19706 11994
rect 19706 11942 19752 11994
rect 19776 11942 19822 11994
rect 19822 11942 19832 11994
rect 19856 11942 19886 11994
rect 19886 11942 19912 11994
rect 19616 11940 19672 11942
rect 19696 11940 19752 11942
rect 19776 11940 19832 11942
rect 19856 11940 19912 11942
rect 20626 13504 20682 13560
rect 19616 10906 19672 10908
rect 19696 10906 19752 10908
rect 19776 10906 19832 10908
rect 19856 10906 19912 10908
rect 19616 10854 19642 10906
rect 19642 10854 19672 10906
rect 19696 10854 19706 10906
rect 19706 10854 19752 10906
rect 19776 10854 19822 10906
rect 19822 10854 19832 10906
rect 19856 10854 19886 10906
rect 19886 10854 19912 10906
rect 19616 10852 19672 10854
rect 19696 10852 19752 10854
rect 19776 10852 19832 10854
rect 19856 10852 19912 10854
rect 18970 10140 18972 10160
rect 18972 10140 19024 10160
rect 19024 10140 19026 10160
rect 18970 10104 19026 10140
rect 19246 8880 19302 8936
rect 19338 8336 19394 8392
rect 19616 9818 19672 9820
rect 19696 9818 19752 9820
rect 19776 9818 19832 9820
rect 19856 9818 19912 9820
rect 19616 9766 19642 9818
rect 19642 9766 19672 9818
rect 19696 9766 19706 9818
rect 19706 9766 19752 9818
rect 19776 9766 19822 9818
rect 19822 9766 19832 9818
rect 19856 9766 19886 9818
rect 19886 9766 19912 9818
rect 19616 9764 19672 9766
rect 19696 9764 19752 9766
rect 19776 9764 19832 9766
rect 19856 9764 19912 9766
rect 19522 9152 19578 9208
rect 19614 8916 19616 8936
rect 19616 8916 19668 8936
rect 19668 8916 19670 8936
rect 19614 8880 19670 8916
rect 19616 8730 19672 8732
rect 19696 8730 19752 8732
rect 19776 8730 19832 8732
rect 19856 8730 19912 8732
rect 19616 8678 19642 8730
rect 19642 8678 19672 8730
rect 19696 8678 19706 8730
rect 19706 8678 19752 8730
rect 19776 8678 19822 8730
rect 19822 8678 19832 8730
rect 19856 8678 19886 8730
rect 19886 8678 19912 8730
rect 19616 8676 19672 8678
rect 19696 8676 19752 8678
rect 19776 8676 19832 8678
rect 19856 8676 19912 8678
rect 19338 6976 19394 7032
rect 19430 6876 19432 6896
rect 19432 6876 19484 6896
rect 19484 6876 19486 6896
rect 19430 6840 19486 6876
rect 19798 8200 19854 8256
rect 19616 7642 19672 7644
rect 19696 7642 19752 7644
rect 19776 7642 19832 7644
rect 19856 7642 19912 7644
rect 19616 7590 19642 7642
rect 19642 7590 19672 7642
rect 19696 7590 19706 7642
rect 19706 7590 19752 7642
rect 19776 7590 19822 7642
rect 19822 7590 19832 7642
rect 19856 7590 19886 7642
rect 19886 7590 19912 7642
rect 19616 7588 19672 7590
rect 19696 7588 19752 7590
rect 19776 7588 19832 7590
rect 19856 7588 19912 7590
rect 19614 7420 19616 7440
rect 19616 7420 19668 7440
rect 19668 7420 19670 7440
rect 19614 7384 19670 7420
rect 19338 6316 19394 6352
rect 19338 6296 19340 6316
rect 19340 6296 19392 6316
rect 19392 6296 19394 6316
rect 19616 6554 19672 6556
rect 19696 6554 19752 6556
rect 19776 6554 19832 6556
rect 19856 6554 19912 6556
rect 19616 6502 19642 6554
rect 19642 6502 19672 6554
rect 19696 6502 19706 6554
rect 19706 6502 19752 6554
rect 19776 6502 19822 6554
rect 19822 6502 19832 6554
rect 19856 6502 19886 6554
rect 19886 6502 19912 6554
rect 19616 6500 19672 6502
rect 19696 6500 19752 6502
rect 19776 6500 19832 6502
rect 19856 6500 19912 6502
rect 19798 6296 19854 6352
rect 19338 6060 19340 6080
rect 19340 6060 19392 6080
rect 19392 6060 19394 6080
rect 19338 6024 19394 6060
rect 19430 5888 19486 5944
rect 20442 8880 20498 8936
rect 21914 12824 21970 12880
rect 21730 10920 21786 10976
rect 20166 5616 20222 5672
rect 19616 5466 19672 5468
rect 19696 5466 19752 5468
rect 19776 5466 19832 5468
rect 19856 5466 19912 5468
rect 19616 5414 19642 5466
rect 19642 5414 19672 5466
rect 19696 5414 19706 5466
rect 19706 5414 19752 5466
rect 19776 5414 19822 5466
rect 19822 5414 19832 5466
rect 19856 5414 19886 5466
rect 19886 5414 19912 5466
rect 19616 5412 19672 5414
rect 19696 5412 19752 5414
rect 19776 5412 19832 5414
rect 19856 5412 19912 5414
rect 19616 4378 19672 4380
rect 19696 4378 19752 4380
rect 19776 4378 19832 4380
rect 19856 4378 19912 4380
rect 19616 4326 19642 4378
rect 19642 4326 19672 4378
rect 19696 4326 19706 4378
rect 19706 4326 19752 4378
rect 19776 4326 19822 4378
rect 19822 4326 19832 4378
rect 19856 4326 19886 4378
rect 19886 4326 19912 4378
rect 19616 4324 19672 4326
rect 19696 4324 19752 4326
rect 19776 4324 19832 4326
rect 19856 4324 19912 4326
rect 15884 2746 15940 2748
rect 15964 2746 16020 2748
rect 16044 2746 16100 2748
rect 16124 2746 16180 2748
rect 15884 2694 15910 2746
rect 15910 2694 15940 2746
rect 15964 2694 15974 2746
rect 15974 2694 16020 2746
rect 16044 2694 16090 2746
rect 16090 2694 16100 2746
rect 16124 2694 16154 2746
rect 16154 2694 16180 2746
rect 15884 2692 15940 2694
rect 15964 2692 16020 2694
rect 16044 2692 16100 2694
rect 16124 2692 16180 2694
rect 19616 3290 19672 3292
rect 19696 3290 19752 3292
rect 19776 3290 19832 3292
rect 19856 3290 19912 3292
rect 19616 3238 19642 3290
rect 19642 3238 19672 3290
rect 19696 3238 19706 3290
rect 19706 3238 19752 3290
rect 19776 3238 19822 3290
rect 19822 3238 19832 3290
rect 19856 3238 19886 3290
rect 19886 3238 19912 3290
rect 19616 3236 19672 3238
rect 19696 3236 19752 3238
rect 19776 3236 19832 3238
rect 19856 3236 19912 3238
rect 20534 5888 20590 5944
rect 20442 4256 20498 4312
rect 21822 8236 21824 8256
rect 21824 8236 21876 8256
rect 21876 8236 21878 8256
rect 21822 8200 21878 8236
rect 22834 20848 22890 20904
rect 22834 19508 22890 19544
rect 22834 19488 22836 19508
rect 22836 19488 22888 19508
rect 22888 19488 22890 19508
rect 23110 18264 23166 18320
rect 23110 17620 23112 17640
rect 23112 17620 23164 17640
rect 23164 17620 23166 17640
rect 23110 17584 23166 17620
rect 23110 16904 23166 16960
rect 23570 22208 23626 22264
rect 23018 12280 23074 12336
rect 22926 10240 22982 10296
rect 22282 7404 22338 7440
rect 22282 7384 22284 7404
rect 22284 7384 22336 7404
rect 22336 7384 22338 7404
rect 22282 6840 22338 6896
rect 21178 4936 21234 4992
rect 12152 2202 12208 2204
rect 12232 2202 12288 2204
rect 12312 2202 12368 2204
rect 12392 2202 12448 2204
rect 12152 2150 12178 2202
rect 12178 2150 12208 2202
rect 12232 2150 12242 2202
rect 12242 2150 12288 2202
rect 12312 2150 12358 2202
rect 12358 2150 12368 2202
rect 12392 2150 12422 2202
rect 12422 2150 12448 2202
rect 12152 2148 12208 2150
rect 12232 2148 12288 2150
rect 12312 2148 12368 2150
rect 12392 2148 12448 2150
rect 19616 2202 19672 2204
rect 19696 2202 19752 2204
rect 19776 2202 19832 2204
rect 19856 2202 19912 2204
rect 19616 2150 19642 2202
rect 19642 2150 19672 2202
rect 19696 2150 19706 2202
rect 19706 2150 19752 2202
rect 19776 2150 19822 2202
rect 19822 2150 19832 2202
rect 19856 2150 19886 2202
rect 19886 2150 19912 2202
rect 19616 2148 19672 2150
rect 19696 2148 19752 2150
rect 19776 2148 19832 2150
rect 19856 2148 19912 2150
rect 22466 6316 22522 6352
rect 22466 6296 22468 6316
rect 22468 6296 22520 6316
rect 22520 6296 22522 6316
rect 22742 9560 22798 9616
rect 23110 9696 23166 9752
rect 22926 8200 22982 8256
rect 23018 7520 23074 7576
rect 23018 6976 23074 7032
rect 22558 3576 22614 3632
rect 23386 9696 23442 9752
rect 23386 2896 23442 2952
rect 23570 6024 23626 6080
rect 23570 2216 23626 2272
rect 23662 1536 23718 1592
rect 23478 856 23534 912
rect 21914 312 21970 368
<< metal3 >>
rect 21817 24306 21883 24309
rect 23800 24306 24600 24336
rect 21817 24304 24600 24306
rect 21817 24248 21822 24304
rect 21878 24248 24600 24304
rect 21817 24246 24600 24248
rect 21817 24243 21883 24246
rect 23800 24216 24600 24246
rect 21909 23626 21975 23629
rect 23800 23626 24600 23656
rect 21909 23624 24600 23626
rect 21909 23568 21914 23624
rect 21970 23568 24600 23624
rect 21909 23566 24600 23568
rect 21909 23563 21975 23566
rect 23800 23536 24600 23566
rect 22001 22946 22067 22949
rect 23800 22946 24600 22976
rect 22001 22944 24600 22946
rect 22001 22888 22006 22944
rect 22062 22888 24600 22944
rect 22001 22886 24600 22888
rect 22001 22883 22067 22886
rect 23800 22856 24600 22886
rect 8408 22336 8728 22337
rect 8408 22272 8416 22336
rect 8480 22272 8496 22336
rect 8560 22272 8576 22336
rect 8640 22272 8656 22336
rect 8720 22272 8728 22336
rect 8408 22271 8728 22272
rect 15872 22336 16192 22337
rect 15872 22272 15880 22336
rect 15944 22272 15960 22336
rect 16024 22272 16040 22336
rect 16104 22272 16120 22336
rect 16184 22272 16192 22336
rect 15872 22271 16192 22272
rect 23565 22266 23631 22269
rect 23800 22266 24600 22296
rect 23565 22264 24600 22266
rect 23565 22208 23570 22264
rect 23626 22208 24600 22264
rect 23565 22206 24600 22208
rect 23565 22203 23631 22206
rect 23800 22176 24600 22206
rect 4676 21792 4996 21793
rect 4676 21728 4684 21792
rect 4748 21728 4764 21792
rect 4828 21728 4844 21792
rect 4908 21728 4924 21792
rect 4988 21728 4996 21792
rect 4676 21727 4996 21728
rect 12140 21792 12460 21793
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 21727 12460 21728
rect 19604 21792 19924 21793
rect 19604 21728 19612 21792
rect 19676 21728 19692 21792
rect 19756 21728 19772 21792
rect 19836 21728 19852 21792
rect 19916 21728 19924 21792
rect 19604 21727 19924 21728
rect 2313 21586 2379 21589
rect 8293 21586 8359 21589
rect 2313 21584 8359 21586
rect 2313 21528 2318 21584
rect 2374 21528 8298 21584
rect 8354 21528 8359 21584
rect 2313 21526 8359 21528
rect 2313 21523 2379 21526
rect 8293 21523 8359 21526
rect 12893 21586 12959 21589
rect 15745 21586 15811 21589
rect 12893 21584 15811 21586
rect 12893 21528 12898 21584
rect 12954 21528 15750 21584
rect 15806 21528 15811 21584
rect 12893 21526 15811 21528
rect 12893 21523 12959 21526
rect 15745 21523 15811 21526
rect 22461 21586 22527 21589
rect 23800 21586 24600 21616
rect 22461 21584 24600 21586
rect 22461 21528 22466 21584
rect 22522 21528 24600 21584
rect 22461 21526 24600 21528
rect 22461 21523 22527 21526
rect 23800 21496 24600 21526
rect 0 21360 800 21480
rect 10041 21450 10107 21453
rect 17401 21450 17467 21453
rect 10041 21448 17467 21450
rect 10041 21392 10046 21448
rect 10102 21392 17406 21448
rect 17462 21392 17467 21448
rect 10041 21390 17467 21392
rect 10041 21387 10107 21390
rect 17401 21387 17467 21390
rect 8408 21248 8728 21249
rect 8408 21184 8416 21248
rect 8480 21184 8496 21248
rect 8560 21184 8576 21248
rect 8640 21184 8656 21248
rect 8720 21184 8728 21248
rect 8408 21183 8728 21184
rect 15872 21248 16192 21249
rect 15872 21184 15880 21248
rect 15944 21184 15960 21248
rect 16024 21184 16040 21248
rect 16104 21184 16120 21248
rect 16184 21184 16192 21248
rect 15872 21183 16192 21184
rect 11605 21042 11671 21045
rect 14917 21042 14983 21045
rect 11605 21040 14983 21042
rect 11605 20984 11610 21040
rect 11666 20984 14922 21040
rect 14978 20984 14983 21040
rect 11605 20982 14983 20984
rect 11605 20979 11671 20982
rect 14917 20979 14983 20982
rect 22829 20906 22895 20909
rect 23800 20906 24600 20936
rect 22829 20904 24600 20906
rect 22829 20848 22834 20904
rect 22890 20848 24600 20904
rect 22829 20846 24600 20848
rect 22829 20843 22895 20846
rect 23800 20816 24600 20846
rect 4676 20704 4996 20705
rect 4676 20640 4684 20704
rect 4748 20640 4764 20704
rect 4828 20640 4844 20704
rect 4908 20640 4924 20704
rect 4988 20640 4996 20704
rect 4676 20639 4996 20640
rect 12140 20704 12460 20705
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 20639 12460 20640
rect 19604 20704 19924 20705
rect 19604 20640 19612 20704
rect 19676 20640 19692 20704
rect 19756 20640 19772 20704
rect 19836 20640 19852 20704
rect 19916 20640 19924 20704
rect 19604 20639 19924 20640
rect 1577 20498 1643 20501
rect 4613 20498 4679 20501
rect 1577 20496 4679 20498
rect 1577 20440 1582 20496
rect 1638 20440 4618 20496
rect 4674 20440 4679 20496
rect 1577 20438 4679 20440
rect 1577 20435 1643 20438
rect 4613 20435 4679 20438
rect 4981 20498 5047 20501
rect 5993 20498 6059 20501
rect 4981 20496 6059 20498
rect 4981 20440 4986 20496
rect 5042 20440 5998 20496
rect 6054 20440 6059 20496
rect 4981 20438 6059 20440
rect 4981 20435 5047 20438
rect 5993 20435 6059 20438
rect 22461 20226 22527 20229
rect 23800 20226 24600 20256
rect 22461 20224 24600 20226
rect 22461 20168 22466 20224
rect 22522 20168 24600 20224
rect 22461 20166 24600 20168
rect 22461 20163 22527 20166
rect 8408 20160 8728 20161
rect 8408 20096 8416 20160
rect 8480 20096 8496 20160
rect 8560 20096 8576 20160
rect 8640 20096 8656 20160
rect 8720 20096 8728 20160
rect 8408 20095 8728 20096
rect 15872 20160 16192 20161
rect 15872 20096 15880 20160
rect 15944 20096 15960 20160
rect 16024 20096 16040 20160
rect 16104 20096 16120 20160
rect 16184 20096 16192 20160
rect 23800 20136 24600 20166
rect 15872 20095 16192 20096
rect 16573 20090 16639 20093
rect 17493 20090 17559 20093
rect 16573 20088 17559 20090
rect 16573 20032 16578 20088
rect 16634 20032 17498 20088
rect 17554 20032 17559 20088
rect 16573 20030 17559 20032
rect 16573 20027 16639 20030
rect 17493 20027 17559 20030
rect 11881 19954 11947 19957
rect 12525 19954 12591 19957
rect 11881 19952 12591 19954
rect 11881 19896 11886 19952
rect 11942 19896 12530 19952
rect 12586 19896 12591 19952
rect 11881 19894 12591 19896
rect 11881 19891 11947 19894
rect 12525 19891 12591 19894
rect 13353 19818 13419 19821
rect 13905 19818 13971 19821
rect 13353 19816 13971 19818
rect 13353 19760 13358 19816
rect 13414 19760 13910 19816
rect 13966 19760 13971 19816
rect 13353 19758 13971 19760
rect 13353 19755 13419 19758
rect 13905 19755 13971 19758
rect 4676 19616 4996 19617
rect 4676 19552 4684 19616
rect 4748 19552 4764 19616
rect 4828 19552 4844 19616
rect 4908 19552 4924 19616
rect 4988 19552 4996 19616
rect 4676 19551 4996 19552
rect 12140 19616 12460 19617
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 19551 12460 19552
rect 19604 19616 19924 19617
rect 19604 19552 19612 19616
rect 19676 19552 19692 19616
rect 19756 19552 19772 19616
rect 19836 19552 19852 19616
rect 19916 19552 19924 19616
rect 19604 19551 19924 19552
rect 14917 19546 14983 19549
rect 19149 19546 19215 19549
rect 14917 19544 19215 19546
rect 14917 19488 14922 19544
rect 14978 19488 19154 19544
rect 19210 19488 19215 19544
rect 14917 19486 19215 19488
rect 14917 19483 14983 19486
rect 19149 19483 19215 19486
rect 22829 19546 22895 19549
rect 23800 19546 24600 19576
rect 22829 19544 24600 19546
rect 22829 19488 22834 19544
rect 22890 19488 24600 19544
rect 22829 19486 24600 19488
rect 22829 19483 22895 19486
rect 23800 19456 24600 19486
rect 8017 19410 8083 19413
rect 9121 19410 9187 19413
rect 8017 19408 9187 19410
rect 8017 19352 8022 19408
rect 8078 19352 9126 19408
rect 9182 19352 9187 19408
rect 8017 19350 9187 19352
rect 8017 19347 8083 19350
rect 9121 19347 9187 19350
rect 12433 19410 12499 19413
rect 19333 19410 19399 19413
rect 12433 19408 19399 19410
rect 12433 19352 12438 19408
rect 12494 19352 19338 19408
rect 19394 19352 19399 19408
rect 12433 19350 19399 19352
rect 12433 19347 12499 19350
rect 19333 19347 19399 19350
rect 11697 19274 11763 19277
rect 16941 19274 17007 19277
rect 11697 19272 17007 19274
rect 11697 19216 11702 19272
rect 11758 19216 16946 19272
rect 17002 19216 17007 19272
rect 11697 19214 17007 19216
rect 11697 19211 11763 19214
rect 16941 19211 17007 19214
rect 8408 19072 8728 19073
rect 8408 19008 8416 19072
rect 8480 19008 8496 19072
rect 8560 19008 8576 19072
rect 8640 19008 8656 19072
rect 8720 19008 8728 19072
rect 8408 19007 8728 19008
rect 15872 19072 16192 19073
rect 15872 19008 15880 19072
rect 15944 19008 15960 19072
rect 16024 19008 16040 19072
rect 16104 19008 16120 19072
rect 16184 19008 16192 19072
rect 15872 19007 16192 19008
rect 15653 19002 15719 19005
rect 15653 19000 15762 19002
rect 15653 18944 15658 19000
rect 15714 18944 15762 19000
rect 15653 18939 15762 18944
rect 15702 18866 15762 18939
rect 16297 18866 16363 18869
rect 15702 18864 16363 18866
rect 15702 18808 16302 18864
rect 16358 18808 16363 18864
rect 15702 18806 16363 18808
rect 16297 18803 16363 18806
rect 21173 18866 21239 18869
rect 23800 18866 24600 18896
rect 21173 18864 24600 18866
rect 21173 18808 21178 18864
rect 21234 18808 24600 18864
rect 21173 18806 24600 18808
rect 21173 18803 21239 18806
rect 23800 18776 24600 18806
rect 15101 18730 15167 18733
rect 16849 18730 16915 18733
rect 15101 18728 16915 18730
rect 15101 18672 15106 18728
rect 15162 18672 16854 18728
rect 16910 18672 16915 18728
rect 15101 18670 16915 18672
rect 15101 18667 15167 18670
rect 16849 18667 16915 18670
rect 4676 18528 4996 18529
rect 4676 18464 4684 18528
rect 4748 18464 4764 18528
rect 4828 18464 4844 18528
rect 4908 18464 4924 18528
rect 4988 18464 4996 18528
rect 4676 18463 4996 18464
rect 12140 18528 12460 18529
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 18463 12460 18464
rect 19604 18528 19924 18529
rect 19604 18464 19612 18528
rect 19676 18464 19692 18528
rect 19756 18464 19772 18528
rect 19836 18464 19852 18528
rect 19916 18464 19924 18528
rect 19604 18463 19924 18464
rect 23105 18322 23171 18325
rect 23800 18322 24600 18352
rect 23105 18320 24600 18322
rect 23105 18264 23110 18320
rect 23166 18264 24600 18320
rect 23105 18262 24600 18264
rect 23105 18259 23171 18262
rect 23800 18232 24600 18262
rect 8408 17984 8728 17985
rect 8408 17920 8416 17984
rect 8480 17920 8496 17984
rect 8560 17920 8576 17984
rect 8640 17920 8656 17984
rect 8720 17920 8728 17984
rect 8408 17919 8728 17920
rect 15872 17984 16192 17985
rect 15872 17920 15880 17984
rect 15944 17920 15960 17984
rect 16024 17920 16040 17984
rect 16104 17920 16120 17984
rect 16184 17920 16192 17984
rect 15872 17919 16192 17920
rect 12433 17642 12499 17645
rect 13353 17642 13419 17645
rect 14641 17642 14707 17645
rect 15377 17642 15443 17645
rect 12433 17640 15443 17642
rect 12433 17584 12438 17640
rect 12494 17584 13358 17640
rect 13414 17584 14646 17640
rect 14702 17584 15382 17640
rect 15438 17584 15443 17640
rect 12433 17582 15443 17584
rect 12433 17579 12499 17582
rect 13353 17579 13419 17582
rect 14641 17579 14707 17582
rect 15377 17579 15443 17582
rect 23105 17642 23171 17645
rect 23800 17642 24600 17672
rect 23105 17640 24600 17642
rect 23105 17584 23110 17640
rect 23166 17584 24600 17640
rect 23105 17582 24600 17584
rect 23105 17579 23171 17582
rect 23800 17552 24600 17582
rect 4676 17440 4996 17441
rect 4676 17376 4684 17440
rect 4748 17376 4764 17440
rect 4828 17376 4844 17440
rect 4908 17376 4924 17440
rect 4988 17376 4996 17440
rect 4676 17375 4996 17376
rect 12140 17440 12460 17441
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 17375 12460 17376
rect 19604 17440 19924 17441
rect 19604 17376 19612 17440
rect 19676 17376 19692 17440
rect 19756 17376 19772 17440
rect 19836 17376 19852 17440
rect 19916 17376 19924 17440
rect 19604 17375 19924 17376
rect 23105 16962 23171 16965
rect 23800 16962 24600 16992
rect 23105 16960 24600 16962
rect 23105 16904 23110 16960
rect 23166 16904 24600 16960
rect 23105 16902 24600 16904
rect 23105 16899 23171 16902
rect 8408 16896 8728 16897
rect 8408 16832 8416 16896
rect 8480 16832 8496 16896
rect 8560 16832 8576 16896
rect 8640 16832 8656 16896
rect 8720 16832 8728 16896
rect 8408 16831 8728 16832
rect 15872 16896 16192 16897
rect 15872 16832 15880 16896
rect 15944 16832 15960 16896
rect 16024 16832 16040 16896
rect 16104 16832 16120 16896
rect 16184 16832 16192 16896
rect 23800 16872 24600 16902
rect 15872 16831 16192 16832
rect 2681 16554 2747 16557
rect 6177 16554 6243 16557
rect 2681 16552 6243 16554
rect 2681 16496 2686 16552
rect 2742 16496 6182 16552
rect 6238 16496 6243 16552
rect 2681 16494 6243 16496
rect 2681 16491 2747 16494
rect 6177 16491 6243 16494
rect 4676 16352 4996 16353
rect 4676 16288 4684 16352
rect 4748 16288 4764 16352
rect 4828 16288 4844 16352
rect 4908 16288 4924 16352
rect 4988 16288 4996 16352
rect 4676 16287 4996 16288
rect 12140 16352 12460 16353
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 16287 12460 16288
rect 19604 16352 19924 16353
rect 19604 16288 19612 16352
rect 19676 16288 19692 16352
rect 19756 16288 19772 16352
rect 19836 16288 19852 16352
rect 19916 16288 19924 16352
rect 19604 16287 19924 16288
rect 20253 16282 20319 16285
rect 23800 16282 24600 16312
rect 20253 16280 24600 16282
rect 20253 16224 20258 16280
rect 20314 16224 24600 16280
rect 20253 16222 24600 16224
rect 20253 16219 20319 16222
rect 23800 16192 24600 16222
rect 8408 15808 8728 15809
rect 8408 15744 8416 15808
rect 8480 15744 8496 15808
rect 8560 15744 8576 15808
rect 8640 15744 8656 15808
rect 8720 15744 8728 15808
rect 8408 15743 8728 15744
rect 15872 15808 16192 15809
rect 15872 15744 15880 15808
rect 15944 15744 15960 15808
rect 16024 15744 16040 15808
rect 16104 15744 16120 15808
rect 16184 15744 16192 15808
rect 15872 15743 16192 15744
rect 19333 15602 19399 15605
rect 23800 15602 24600 15632
rect 19333 15600 24600 15602
rect 19333 15544 19338 15600
rect 19394 15544 24600 15600
rect 19333 15542 24600 15544
rect 19333 15539 19399 15542
rect 23800 15512 24600 15542
rect 0 15330 800 15360
rect 2865 15330 2931 15333
rect 0 15328 2931 15330
rect 0 15272 2870 15328
rect 2926 15272 2931 15328
rect 0 15270 2931 15272
rect 0 15240 800 15270
rect 2865 15267 2931 15270
rect 4676 15264 4996 15265
rect 4676 15200 4684 15264
rect 4748 15200 4764 15264
rect 4828 15200 4844 15264
rect 4908 15200 4924 15264
rect 4988 15200 4996 15264
rect 4676 15199 4996 15200
rect 12140 15264 12460 15265
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 15199 12460 15200
rect 19604 15264 19924 15265
rect 19604 15200 19612 15264
rect 19676 15200 19692 15264
rect 19756 15200 19772 15264
rect 19836 15200 19852 15264
rect 19916 15200 19924 15264
rect 19604 15199 19924 15200
rect 19333 14922 19399 14925
rect 23800 14922 24600 14952
rect 19333 14920 24600 14922
rect 19333 14864 19338 14920
rect 19394 14864 24600 14920
rect 19333 14862 24600 14864
rect 19333 14859 19399 14862
rect 23800 14832 24600 14862
rect 8408 14720 8728 14721
rect 8408 14656 8416 14720
rect 8480 14656 8496 14720
rect 8560 14656 8576 14720
rect 8640 14656 8656 14720
rect 8720 14656 8728 14720
rect 8408 14655 8728 14656
rect 15872 14720 16192 14721
rect 15872 14656 15880 14720
rect 15944 14656 15960 14720
rect 16024 14656 16040 14720
rect 16104 14656 16120 14720
rect 16184 14656 16192 14720
rect 15872 14655 16192 14656
rect 19333 14378 19399 14381
rect 19333 14376 23674 14378
rect 19333 14320 19338 14376
rect 19394 14320 23674 14376
rect 19333 14318 23674 14320
rect 19333 14315 19399 14318
rect 23614 14242 23674 14318
rect 23800 14242 24600 14272
rect 23614 14182 24600 14242
rect 4676 14176 4996 14177
rect 4676 14112 4684 14176
rect 4748 14112 4764 14176
rect 4828 14112 4844 14176
rect 4908 14112 4924 14176
rect 4988 14112 4996 14176
rect 4676 14111 4996 14112
rect 12140 14176 12460 14177
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 14111 12460 14112
rect 19604 14176 19924 14177
rect 19604 14112 19612 14176
rect 19676 14112 19692 14176
rect 19756 14112 19772 14176
rect 19836 14112 19852 14176
rect 19916 14112 19924 14176
rect 23800 14152 24600 14182
rect 19604 14111 19924 14112
rect 2681 13834 2747 13837
rect 6269 13834 6335 13837
rect 2681 13832 6335 13834
rect 2681 13776 2686 13832
rect 2742 13776 6274 13832
rect 6330 13776 6335 13832
rect 2681 13774 6335 13776
rect 2681 13771 2747 13774
rect 6269 13771 6335 13774
rect 10501 13834 10567 13837
rect 12893 13834 12959 13837
rect 10501 13832 12959 13834
rect 10501 13776 10506 13832
rect 10562 13776 12898 13832
rect 12954 13776 12959 13832
rect 10501 13774 12959 13776
rect 10501 13771 10567 13774
rect 12893 13771 12959 13774
rect 8408 13632 8728 13633
rect 8408 13568 8416 13632
rect 8480 13568 8496 13632
rect 8560 13568 8576 13632
rect 8640 13568 8656 13632
rect 8720 13568 8728 13632
rect 8408 13567 8728 13568
rect 15872 13632 16192 13633
rect 15872 13568 15880 13632
rect 15944 13568 15960 13632
rect 16024 13568 16040 13632
rect 16104 13568 16120 13632
rect 16184 13568 16192 13632
rect 15872 13567 16192 13568
rect 20621 13562 20687 13565
rect 23800 13562 24600 13592
rect 20621 13560 24600 13562
rect 20621 13504 20626 13560
rect 20682 13504 24600 13560
rect 20621 13502 24600 13504
rect 20621 13499 20687 13502
rect 23800 13472 24600 13502
rect 4676 13088 4996 13089
rect 4676 13024 4684 13088
rect 4748 13024 4764 13088
rect 4828 13024 4844 13088
rect 4908 13024 4924 13088
rect 4988 13024 4996 13088
rect 4676 13023 4996 13024
rect 12140 13088 12460 13089
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 13023 12460 13024
rect 19604 13088 19924 13089
rect 19604 13024 19612 13088
rect 19676 13024 19692 13088
rect 19756 13024 19772 13088
rect 19836 13024 19852 13088
rect 19916 13024 19924 13088
rect 19604 13023 19924 13024
rect 21909 12882 21975 12885
rect 23800 12882 24600 12912
rect 21909 12880 24600 12882
rect 21909 12824 21914 12880
rect 21970 12824 24600 12880
rect 21909 12822 24600 12824
rect 21909 12819 21975 12822
rect 23800 12792 24600 12822
rect 8408 12544 8728 12545
rect 8408 12480 8416 12544
rect 8480 12480 8496 12544
rect 8560 12480 8576 12544
rect 8640 12480 8656 12544
rect 8720 12480 8728 12544
rect 8408 12479 8728 12480
rect 15872 12544 16192 12545
rect 15872 12480 15880 12544
rect 15944 12480 15960 12544
rect 16024 12480 16040 12544
rect 16104 12480 16120 12544
rect 16184 12480 16192 12544
rect 15872 12479 16192 12480
rect 23013 12338 23079 12341
rect 23800 12338 24600 12368
rect 23013 12336 24600 12338
rect 23013 12280 23018 12336
rect 23074 12280 24600 12336
rect 23013 12278 24600 12280
rect 23013 12275 23079 12278
rect 23800 12248 24600 12278
rect 4676 12000 4996 12001
rect 4676 11936 4684 12000
rect 4748 11936 4764 12000
rect 4828 11936 4844 12000
rect 4908 11936 4924 12000
rect 4988 11936 4996 12000
rect 4676 11935 4996 11936
rect 12140 12000 12460 12001
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 11935 12460 11936
rect 19604 12000 19924 12001
rect 19604 11936 19612 12000
rect 19676 11936 19692 12000
rect 19756 11936 19772 12000
rect 19836 11936 19852 12000
rect 19916 11936 19924 12000
rect 19604 11935 19924 11936
rect 19425 11658 19491 11661
rect 23800 11658 24600 11688
rect 19425 11656 24600 11658
rect 19425 11600 19430 11656
rect 19486 11600 24600 11656
rect 19425 11598 24600 11600
rect 19425 11595 19491 11598
rect 23800 11568 24600 11598
rect 8408 11456 8728 11457
rect 8408 11392 8416 11456
rect 8480 11392 8496 11456
rect 8560 11392 8576 11456
rect 8640 11392 8656 11456
rect 8720 11392 8728 11456
rect 8408 11391 8728 11392
rect 15872 11456 16192 11457
rect 15872 11392 15880 11456
rect 15944 11392 15960 11456
rect 16024 11392 16040 11456
rect 16104 11392 16120 11456
rect 16184 11392 16192 11456
rect 15872 11391 16192 11392
rect 21725 10978 21791 10981
rect 23800 10978 24600 11008
rect 21725 10976 24600 10978
rect 21725 10920 21730 10976
rect 21786 10920 24600 10976
rect 21725 10918 24600 10920
rect 21725 10915 21791 10918
rect 4676 10912 4996 10913
rect 4676 10848 4684 10912
rect 4748 10848 4764 10912
rect 4828 10848 4844 10912
rect 4908 10848 4924 10912
rect 4988 10848 4996 10912
rect 4676 10847 4996 10848
rect 12140 10912 12460 10913
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 10847 12460 10848
rect 19604 10912 19924 10913
rect 19604 10848 19612 10912
rect 19676 10848 19692 10912
rect 19756 10848 19772 10912
rect 19836 10848 19852 10912
rect 19916 10848 19924 10912
rect 23800 10888 24600 10918
rect 19604 10847 19924 10848
rect 8408 10368 8728 10369
rect 8408 10304 8416 10368
rect 8480 10304 8496 10368
rect 8560 10304 8576 10368
rect 8640 10304 8656 10368
rect 8720 10304 8728 10368
rect 8408 10303 8728 10304
rect 15872 10368 16192 10369
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 10303 16192 10304
rect 22921 10298 22987 10301
rect 23800 10298 24600 10328
rect 22921 10296 24600 10298
rect 22921 10240 22926 10296
rect 22982 10240 24600 10296
rect 22921 10238 24600 10240
rect 22921 10235 22987 10238
rect 23800 10208 24600 10238
rect 15009 10162 15075 10165
rect 18413 10162 18479 10165
rect 18965 10162 19031 10165
rect 15009 10160 19031 10162
rect 15009 10104 15014 10160
rect 15070 10104 18418 10160
rect 18474 10104 18970 10160
rect 19026 10104 19031 10160
rect 15009 10102 19031 10104
rect 15009 10099 15075 10102
rect 18413 10099 18479 10102
rect 18965 10099 19031 10102
rect 4676 9824 4996 9825
rect 4676 9760 4684 9824
rect 4748 9760 4764 9824
rect 4828 9760 4844 9824
rect 4908 9760 4924 9824
rect 4988 9760 4996 9824
rect 4676 9759 4996 9760
rect 12140 9824 12460 9825
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 9759 12460 9760
rect 19604 9824 19924 9825
rect 19604 9760 19612 9824
rect 19676 9760 19692 9824
rect 19756 9760 19772 9824
rect 19836 9760 19852 9824
rect 19916 9760 19924 9824
rect 19604 9759 19924 9760
rect 23105 9754 23171 9757
rect 23381 9754 23447 9757
rect 23105 9752 23447 9754
rect 23105 9696 23110 9752
rect 23166 9696 23386 9752
rect 23442 9696 23447 9752
rect 23105 9694 23447 9696
rect 23105 9691 23171 9694
rect 23381 9691 23447 9694
rect 22737 9618 22803 9621
rect 23800 9618 24600 9648
rect 22737 9616 24600 9618
rect 22737 9560 22742 9616
rect 22798 9560 24600 9616
rect 22737 9558 24600 9560
rect 22737 9555 22803 9558
rect 23800 9528 24600 9558
rect 8408 9280 8728 9281
rect 0 9210 800 9240
rect 8408 9216 8416 9280
rect 8480 9216 8496 9280
rect 8560 9216 8576 9280
rect 8640 9216 8656 9280
rect 8720 9216 8728 9280
rect 8408 9215 8728 9216
rect 15872 9280 16192 9281
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 9215 16192 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 19374 9148 19380 9212
rect 19444 9210 19450 9212
rect 19517 9210 19583 9213
rect 19444 9208 19583 9210
rect 19444 9152 19522 9208
rect 19578 9152 19583 9208
rect 19444 9150 19583 9152
rect 19444 9148 19450 9150
rect 19517 9147 19583 9150
rect 14917 9074 14983 9077
rect 15653 9074 15719 9077
rect 14917 9072 15719 9074
rect 14917 9016 14922 9072
rect 14978 9016 15658 9072
rect 15714 9016 15719 9072
rect 14917 9014 15719 9016
rect 14917 9011 14983 9014
rect 15653 9011 15719 9014
rect 15101 8938 15167 8941
rect 16481 8938 16547 8941
rect 15101 8936 16547 8938
rect 15101 8880 15106 8936
rect 15162 8880 16486 8936
rect 16542 8880 16547 8936
rect 15101 8878 16547 8880
rect 15101 8875 15167 8878
rect 16481 8875 16547 8878
rect 19241 8938 19307 8941
rect 19609 8938 19675 8941
rect 19241 8936 19675 8938
rect 19241 8880 19246 8936
rect 19302 8880 19614 8936
rect 19670 8880 19675 8936
rect 19241 8878 19675 8880
rect 19241 8875 19307 8878
rect 19609 8875 19675 8878
rect 20437 8938 20503 8941
rect 23800 8938 24600 8968
rect 20437 8936 24600 8938
rect 20437 8880 20442 8936
rect 20498 8880 24600 8936
rect 20437 8878 24600 8880
rect 20437 8875 20503 8878
rect 23800 8848 24600 8878
rect 4676 8736 4996 8737
rect 4676 8672 4684 8736
rect 4748 8672 4764 8736
rect 4828 8672 4844 8736
rect 4908 8672 4924 8736
rect 4988 8672 4996 8736
rect 4676 8671 4996 8672
rect 12140 8736 12460 8737
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 8671 12460 8672
rect 19604 8736 19924 8737
rect 19604 8672 19612 8736
rect 19676 8672 19692 8736
rect 19756 8672 19772 8736
rect 19836 8672 19852 8736
rect 19916 8672 19924 8736
rect 19604 8671 19924 8672
rect 11697 8530 11763 8533
rect 12157 8530 12223 8533
rect 15745 8530 15811 8533
rect 11697 8528 15811 8530
rect 11697 8472 11702 8528
rect 11758 8472 12162 8528
rect 12218 8472 15750 8528
rect 15806 8472 15811 8528
rect 11697 8470 15811 8472
rect 11697 8467 11763 8470
rect 12157 8467 12223 8470
rect 15745 8467 15811 8470
rect 19333 8396 19399 8397
rect 19333 8392 19380 8396
rect 19444 8394 19450 8396
rect 19333 8336 19338 8392
rect 19333 8332 19380 8336
rect 19444 8334 19490 8394
rect 19444 8332 19450 8334
rect 19333 8331 19399 8332
rect 19793 8258 19859 8261
rect 21817 8258 21883 8261
rect 19793 8256 21883 8258
rect 19793 8200 19798 8256
rect 19854 8200 21822 8256
rect 21878 8200 21883 8256
rect 19793 8198 21883 8200
rect 19793 8195 19859 8198
rect 21817 8195 21883 8198
rect 22921 8258 22987 8261
rect 23800 8258 24600 8288
rect 22921 8256 24600 8258
rect 22921 8200 22926 8256
rect 22982 8200 24600 8256
rect 22921 8198 24600 8200
rect 22921 8195 22987 8198
rect 8408 8192 8728 8193
rect 8408 8128 8416 8192
rect 8480 8128 8496 8192
rect 8560 8128 8576 8192
rect 8640 8128 8656 8192
rect 8720 8128 8728 8192
rect 8408 8127 8728 8128
rect 15872 8192 16192 8193
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 23800 8168 24600 8198
rect 15872 8127 16192 8128
rect 14917 8122 14983 8125
rect 15561 8122 15627 8125
rect 14917 8120 15627 8122
rect 14917 8064 14922 8120
rect 14978 8064 15566 8120
rect 15622 8064 15627 8120
rect 14917 8062 15627 8064
rect 14917 8059 14983 8062
rect 15561 8059 15627 8062
rect 14733 7986 14799 7989
rect 16021 7986 16087 7989
rect 17401 7986 17467 7989
rect 14733 7984 17467 7986
rect 14733 7928 14738 7984
rect 14794 7928 16026 7984
rect 16082 7928 17406 7984
rect 17462 7928 17467 7984
rect 14733 7926 17467 7928
rect 14733 7923 14799 7926
rect 16021 7923 16087 7926
rect 17401 7923 17467 7926
rect 4676 7648 4996 7649
rect 4676 7584 4684 7648
rect 4748 7584 4764 7648
rect 4828 7584 4844 7648
rect 4908 7584 4924 7648
rect 4988 7584 4996 7648
rect 4676 7583 4996 7584
rect 12140 7648 12460 7649
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 7583 12460 7584
rect 19604 7648 19924 7649
rect 19604 7584 19612 7648
rect 19676 7584 19692 7648
rect 19756 7584 19772 7648
rect 19836 7584 19852 7648
rect 19916 7584 19924 7648
rect 19604 7583 19924 7584
rect 23013 7578 23079 7581
rect 23800 7578 24600 7608
rect 23013 7576 24600 7578
rect 23013 7520 23018 7576
rect 23074 7520 24600 7576
rect 23013 7518 24600 7520
rect 23013 7515 23079 7518
rect 23800 7488 24600 7518
rect 19609 7442 19675 7445
rect 22277 7442 22343 7445
rect 19609 7440 22343 7442
rect 19609 7384 19614 7440
rect 19670 7384 22282 7440
rect 22338 7384 22343 7440
rect 19609 7382 22343 7384
rect 19609 7379 19675 7382
rect 22277 7379 22343 7382
rect 8408 7104 8728 7105
rect 8408 7040 8416 7104
rect 8480 7040 8496 7104
rect 8560 7040 8576 7104
rect 8640 7040 8656 7104
rect 8720 7040 8728 7104
rect 8408 7039 8728 7040
rect 15872 7104 16192 7105
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 7039 16192 7040
rect 19333 7034 19399 7037
rect 23013 7034 23079 7037
rect 19333 7032 23079 7034
rect 19333 6976 19338 7032
rect 19394 6976 23018 7032
rect 23074 6976 23079 7032
rect 19333 6974 23079 6976
rect 19333 6971 19399 6974
rect 23013 6971 23079 6974
rect 19425 6898 19491 6901
rect 22277 6898 22343 6901
rect 23800 6898 24600 6928
rect 19425 6896 24600 6898
rect 19425 6840 19430 6896
rect 19486 6840 22282 6896
rect 22338 6840 24600 6896
rect 19425 6838 24600 6840
rect 19425 6835 19491 6838
rect 22277 6835 22343 6838
rect 23800 6808 24600 6838
rect 4676 6560 4996 6561
rect 4676 6496 4684 6560
rect 4748 6496 4764 6560
rect 4828 6496 4844 6560
rect 4908 6496 4924 6560
rect 4988 6496 4996 6560
rect 4676 6495 4996 6496
rect 12140 6560 12460 6561
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 6495 12460 6496
rect 19604 6560 19924 6561
rect 19604 6496 19612 6560
rect 19676 6496 19692 6560
rect 19756 6496 19772 6560
rect 19836 6496 19852 6560
rect 19916 6496 19924 6560
rect 19604 6495 19924 6496
rect 19333 6354 19399 6357
rect 19793 6354 19859 6357
rect 19333 6352 19859 6354
rect 19333 6296 19338 6352
rect 19394 6296 19798 6352
rect 19854 6296 19859 6352
rect 19333 6294 19859 6296
rect 19333 6291 19399 6294
rect 19793 6291 19859 6294
rect 22461 6354 22527 6357
rect 23800 6354 24600 6384
rect 22461 6352 24600 6354
rect 22461 6296 22466 6352
rect 22522 6296 24600 6352
rect 22461 6294 24600 6296
rect 22461 6291 22527 6294
rect 23800 6264 24600 6294
rect 19333 6082 19399 6085
rect 23565 6082 23631 6085
rect 19333 6080 23631 6082
rect 19333 6024 19338 6080
rect 19394 6024 23570 6080
rect 23626 6024 23631 6080
rect 19333 6022 23631 6024
rect 19333 6019 19399 6022
rect 23565 6019 23631 6022
rect 8408 6016 8728 6017
rect 8408 5952 8416 6016
rect 8480 5952 8496 6016
rect 8560 5952 8576 6016
rect 8640 5952 8656 6016
rect 8720 5952 8728 6016
rect 8408 5951 8728 5952
rect 15872 6016 16192 6017
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 5951 16192 5952
rect 19425 5946 19491 5949
rect 20529 5946 20595 5949
rect 19425 5944 20595 5946
rect 19425 5888 19430 5944
rect 19486 5888 20534 5944
rect 20590 5888 20595 5944
rect 19425 5886 20595 5888
rect 19425 5883 19491 5886
rect 20529 5883 20595 5886
rect 20161 5674 20227 5677
rect 23800 5674 24600 5704
rect 20161 5672 24600 5674
rect 20161 5616 20166 5672
rect 20222 5616 24600 5672
rect 20161 5614 24600 5616
rect 20161 5611 20227 5614
rect 23800 5584 24600 5614
rect 4676 5472 4996 5473
rect 4676 5408 4684 5472
rect 4748 5408 4764 5472
rect 4828 5408 4844 5472
rect 4908 5408 4924 5472
rect 4988 5408 4996 5472
rect 4676 5407 4996 5408
rect 12140 5472 12460 5473
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 5407 12460 5408
rect 19604 5472 19924 5473
rect 19604 5408 19612 5472
rect 19676 5408 19692 5472
rect 19756 5408 19772 5472
rect 19836 5408 19852 5472
rect 19916 5408 19924 5472
rect 19604 5407 19924 5408
rect 21173 4994 21239 4997
rect 23800 4994 24600 5024
rect 21173 4992 24600 4994
rect 21173 4936 21178 4992
rect 21234 4936 24600 4992
rect 21173 4934 24600 4936
rect 21173 4931 21239 4934
rect 8408 4928 8728 4929
rect 8408 4864 8416 4928
rect 8480 4864 8496 4928
rect 8560 4864 8576 4928
rect 8640 4864 8656 4928
rect 8720 4864 8728 4928
rect 8408 4863 8728 4864
rect 15872 4928 16192 4929
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 23800 4904 24600 4934
rect 15872 4863 16192 4864
rect 4676 4384 4996 4385
rect 4676 4320 4684 4384
rect 4748 4320 4764 4384
rect 4828 4320 4844 4384
rect 4908 4320 4924 4384
rect 4988 4320 4996 4384
rect 4676 4319 4996 4320
rect 12140 4384 12460 4385
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 4319 12460 4320
rect 19604 4384 19924 4385
rect 19604 4320 19612 4384
rect 19676 4320 19692 4384
rect 19756 4320 19772 4384
rect 19836 4320 19852 4384
rect 19916 4320 19924 4384
rect 19604 4319 19924 4320
rect 20437 4314 20503 4317
rect 23800 4314 24600 4344
rect 20437 4312 24600 4314
rect 20437 4256 20442 4312
rect 20498 4256 24600 4312
rect 20437 4254 24600 4256
rect 20437 4251 20503 4254
rect 23800 4224 24600 4254
rect 8408 3840 8728 3841
rect 8408 3776 8416 3840
rect 8480 3776 8496 3840
rect 8560 3776 8576 3840
rect 8640 3776 8656 3840
rect 8720 3776 8728 3840
rect 8408 3775 8728 3776
rect 15872 3840 16192 3841
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 3775 16192 3776
rect 22553 3634 22619 3637
rect 23800 3634 24600 3664
rect 22553 3632 24600 3634
rect 22553 3576 22558 3632
rect 22614 3576 24600 3632
rect 22553 3574 24600 3576
rect 22553 3571 22619 3574
rect 23800 3544 24600 3574
rect 4676 3296 4996 3297
rect 4676 3232 4684 3296
rect 4748 3232 4764 3296
rect 4828 3232 4844 3296
rect 4908 3232 4924 3296
rect 4988 3232 4996 3296
rect 4676 3231 4996 3232
rect 12140 3296 12460 3297
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 3231 12460 3232
rect 19604 3296 19924 3297
rect 19604 3232 19612 3296
rect 19676 3232 19692 3296
rect 19756 3232 19772 3296
rect 19836 3232 19852 3296
rect 19916 3232 19924 3296
rect 19604 3231 19924 3232
rect 0 3090 800 3120
rect 1945 3090 2011 3093
rect 0 3088 2011 3090
rect 0 3032 1950 3088
rect 2006 3032 2011 3088
rect 0 3030 2011 3032
rect 0 3000 800 3030
rect 1945 3027 2011 3030
rect 23381 2954 23447 2957
rect 23800 2954 24600 2984
rect 23381 2952 24600 2954
rect 23381 2896 23386 2952
rect 23442 2896 24600 2952
rect 23381 2894 24600 2896
rect 23381 2891 23447 2894
rect 23800 2864 24600 2894
rect 8408 2752 8728 2753
rect 8408 2688 8416 2752
rect 8480 2688 8496 2752
rect 8560 2688 8576 2752
rect 8640 2688 8656 2752
rect 8720 2688 8728 2752
rect 8408 2687 8728 2688
rect 15872 2752 16192 2753
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 2687 16192 2688
rect 23565 2274 23631 2277
rect 23800 2274 24600 2304
rect 23565 2272 24600 2274
rect 23565 2216 23570 2272
rect 23626 2216 24600 2272
rect 23565 2214 24600 2216
rect 23565 2211 23631 2214
rect 4676 2208 4996 2209
rect 4676 2144 4684 2208
rect 4748 2144 4764 2208
rect 4828 2144 4844 2208
rect 4908 2144 4924 2208
rect 4988 2144 4996 2208
rect 4676 2143 4996 2144
rect 12140 2208 12460 2209
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2143 12460 2144
rect 19604 2208 19924 2209
rect 19604 2144 19612 2208
rect 19676 2144 19692 2208
rect 19756 2144 19772 2208
rect 19836 2144 19852 2208
rect 19916 2144 19924 2208
rect 23800 2184 24600 2214
rect 19604 2143 19924 2144
rect 23657 1594 23723 1597
rect 23800 1594 24600 1624
rect 23657 1592 24600 1594
rect 23657 1536 23662 1592
rect 23718 1536 24600 1592
rect 23657 1534 24600 1536
rect 23657 1531 23723 1534
rect 23800 1504 24600 1534
rect 23473 914 23539 917
rect 23800 914 24600 944
rect 23473 912 24600 914
rect 23473 856 23478 912
rect 23534 856 24600 912
rect 23473 854 24600 856
rect 23473 851 23539 854
rect 23800 824 24600 854
rect 21909 370 21975 373
rect 23800 370 24600 400
rect 21909 368 24600 370
rect 21909 312 21914 368
rect 21970 312 24600 368
rect 21909 310 24600 312
rect 21909 307 21975 310
rect 23800 280 24600 310
<< via3 >>
rect 8416 22332 8480 22336
rect 8416 22276 8420 22332
rect 8420 22276 8476 22332
rect 8476 22276 8480 22332
rect 8416 22272 8480 22276
rect 8496 22332 8560 22336
rect 8496 22276 8500 22332
rect 8500 22276 8556 22332
rect 8556 22276 8560 22332
rect 8496 22272 8560 22276
rect 8576 22332 8640 22336
rect 8576 22276 8580 22332
rect 8580 22276 8636 22332
rect 8636 22276 8640 22332
rect 8576 22272 8640 22276
rect 8656 22332 8720 22336
rect 8656 22276 8660 22332
rect 8660 22276 8716 22332
rect 8716 22276 8720 22332
rect 8656 22272 8720 22276
rect 15880 22332 15944 22336
rect 15880 22276 15884 22332
rect 15884 22276 15940 22332
rect 15940 22276 15944 22332
rect 15880 22272 15944 22276
rect 15960 22332 16024 22336
rect 15960 22276 15964 22332
rect 15964 22276 16020 22332
rect 16020 22276 16024 22332
rect 15960 22272 16024 22276
rect 16040 22332 16104 22336
rect 16040 22276 16044 22332
rect 16044 22276 16100 22332
rect 16100 22276 16104 22332
rect 16040 22272 16104 22276
rect 16120 22332 16184 22336
rect 16120 22276 16124 22332
rect 16124 22276 16180 22332
rect 16180 22276 16184 22332
rect 16120 22272 16184 22276
rect 4684 21788 4748 21792
rect 4684 21732 4688 21788
rect 4688 21732 4744 21788
rect 4744 21732 4748 21788
rect 4684 21728 4748 21732
rect 4764 21788 4828 21792
rect 4764 21732 4768 21788
rect 4768 21732 4824 21788
rect 4824 21732 4828 21788
rect 4764 21728 4828 21732
rect 4844 21788 4908 21792
rect 4844 21732 4848 21788
rect 4848 21732 4904 21788
rect 4904 21732 4908 21788
rect 4844 21728 4908 21732
rect 4924 21788 4988 21792
rect 4924 21732 4928 21788
rect 4928 21732 4984 21788
rect 4984 21732 4988 21788
rect 4924 21728 4988 21732
rect 12148 21788 12212 21792
rect 12148 21732 12152 21788
rect 12152 21732 12208 21788
rect 12208 21732 12212 21788
rect 12148 21728 12212 21732
rect 12228 21788 12292 21792
rect 12228 21732 12232 21788
rect 12232 21732 12288 21788
rect 12288 21732 12292 21788
rect 12228 21728 12292 21732
rect 12308 21788 12372 21792
rect 12308 21732 12312 21788
rect 12312 21732 12368 21788
rect 12368 21732 12372 21788
rect 12308 21728 12372 21732
rect 12388 21788 12452 21792
rect 12388 21732 12392 21788
rect 12392 21732 12448 21788
rect 12448 21732 12452 21788
rect 12388 21728 12452 21732
rect 19612 21788 19676 21792
rect 19612 21732 19616 21788
rect 19616 21732 19672 21788
rect 19672 21732 19676 21788
rect 19612 21728 19676 21732
rect 19692 21788 19756 21792
rect 19692 21732 19696 21788
rect 19696 21732 19752 21788
rect 19752 21732 19756 21788
rect 19692 21728 19756 21732
rect 19772 21788 19836 21792
rect 19772 21732 19776 21788
rect 19776 21732 19832 21788
rect 19832 21732 19836 21788
rect 19772 21728 19836 21732
rect 19852 21788 19916 21792
rect 19852 21732 19856 21788
rect 19856 21732 19912 21788
rect 19912 21732 19916 21788
rect 19852 21728 19916 21732
rect 8416 21244 8480 21248
rect 8416 21188 8420 21244
rect 8420 21188 8476 21244
rect 8476 21188 8480 21244
rect 8416 21184 8480 21188
rect 8496 21244 8560 21248
rect 8496 21188 8500 21244
rect 8500 21188 8556 21244
rect 8556 21188 8560 21244
rect 8496 21184 8560 21188
rect 8576 21244 8640 21248
rect 8576 21188 8580 21244
rect 8580 21188 8636 21244
rect 8636 21188 8640 21244
rect 8576 21184 8640 21188
rect 8656 21244 8720 21248
rect 8656 21188 8660 21244
rect 8660 21188 8716 21244
rect 8716 21188 8720 21244
rect 8656 21184 8720 21188
rect 15880 21244 15944 21248
rect 15880 21188 15884 21244
rect 15884 21188 15940 21244
rect 15940 21188 15944 21244
rect 15880 21184 15944 21188
rect 15960 21244 16024 21248
rect 15960 21188 15964 21244
rect 15964 21188 16020 21244
rect 16020 21188 16024 21244
rect 15960 21184 16024 21188
rect 16040 21244 16104 21248
rect 16040 21188 16044 21244
rect 16044 21188 16100 21244
rect 16100 21188 16104 21244
rect 16040 21184 16104 21188
rect 16120 21244 16184 21248
rect 16120 21188 16124 21244
rect 16124 21188 16180 21244
rect 16180 21188 16184 21244
rect 16120 21184 16184 21188
rect 4684 20700 4748 20704
rect 4684 20644 4688 20700
rect 4688 20644 4744 20700
rect 4744 20644 4748 20700
rect 4684 20640 4748 20644
rect 4764 20700 4828 20704
rect 4764 20644 4768 20700
rect 4768 20644 4824 20700
rect 4824 20644 4828 20700
rect 4764 20640 4828 20644
rect 4844 20700 4908 20704
rect 4844 20644 4848 20700
rect 4848 20644 4904 20700
rect 4904 20644 4908 20700
rect 4844 20640 4908 20644
rect 4924 20700 4988 20704
rect 4924 20644 4928 20700
rect 4928 20644 4984 20700
rect 4984 20644 4988 20700
rect 4924 20640 4988 20644
rect 12148 20700 12212 20704
rect 12148 20644 12152 20700
rect 12152 20644 12208 20700
rect 12208 20644 12212 20700
rect 12148 20640 12212 20644
rect 12228 20700 12292 20704
rect 12228 20644 12232 20700
rect 12232 20644 12288 20700
rect 12288 20644 12292 20700
rect 12228 20640 12292 20644
rect 12308 20700 12372 20704
rect 12308 20644 12312 20700
rect 12312 20644 12368 20700
rect 12368 20644 12372 20700
rect 12308 20640 12372 20644
rect 12388 20700 12452 20704
rect 12388 20644 12392 20700
rect 12392 20644 12448 20700
rect 12448 20644 12452 20700
rect 12388 20640 12452 20644
rect 19612 20700 19676 20704
rect 19612 20644 19616 20700
rect 19616 20644 19672 20700
rect 19672 20644 19676 20700
rect 19612 20640 19676 20644
rect 19692 20700 19756 20704
rect 19692 20644 19696 20700
rect 19696 20644 19752 20700
rect 19752 20644 19756 20700
rect 19692 20640 19756 20644
rect 19772 20700 19836 20704
rect 19772 20644 19776 20700
rect 19776 20644 19832 20700
rect 19832 20644 19836 20700
rect 19772 20640 19836 20644
rect 19852 20700 19916 20704
rect 19852 20644 19856 20700
rect 19856 20644 19912 20700
rect 19912 20644 19916 20700
rect 19852 20640 19916 20644
rect 8416 20156 8480 20160
rect 8416 20100 8420 20156
rect 8420 20100 8476 20156
rect 8476 20100 8480 20156
rect 8416 20096 8480 20100
rect 8496 20156 8560 20160
rect 8496 20100 8500 20156
rect 8500 20100 8556 20156
rect 8556 20100 8560 20156
rect 8496 20096 8560 20100
rect 8576 20156 8640 20160
rect 8576 20100 8580 20156
rect 8580 20100 8636 20156
rect 8636 20100 8640 20156
rect 8576 20096 8640 20100
rect 8656 20156 8720 20160
rect 8656 20100 8660 20156
rect 8660 20100 8716 20156
rect 8716 20100 8720 20156
rect 8656 20096 8720 20100
rect 15880 20156 15944 20160
rect 15880 20100 15884 20156
rect 15884 20100 15940 20156
rect 15940 20100 15944 20156
rect 15880 20096 15944 20100
rect 15960 20156 16024 20160
rect 15960 20100 15964 20156
rect 15964 20100 16020 20156
rect 16020 20100 16024 20156
rect 15960 20096 16024 20100
rect 16040 20156 16104 20160
rect 16040 20100 16044 20156
rect 16044 20100 16100 20156
rect 16100 20100 16104 20156
rect 16040 20096 16104 20100
rect 16120 20156 16184 20160
rect 16120 20100 16124 20156
rect 16124 20100 16180 20156
rect 16180 20100 16184 20156
rect 16120 20096 16184 20100
rect 4684 19612 4748 19616
rect 4684 19556 4688 19612
rect 4688 19556 4744 19612
rect 4744 19556 4748 19612
rect 4684 19552 4748 19556
rect 4764 19612 4828 19616
rect 4764 19556 4768 19612
rect 4768 19556 4824 19612
rect 4824 19556 4828 19612
rect 4764 19552 4828 19556
rect 4844 19612 4908 19616
rect 4844 19556 4848 19612
rect 4848 19556 4904 19612
rect 4904 19556 4908 19612
rect 4844 19552 4908 19556
rect 4924 19612 4988 19616
rect 4924 19556 4928 19612
rect 4928 19556 4984 19612
rect 4984 19556 4988 19612
rect 4924 19552 4988 19556
rect 12148 19612 12212 19616
rect 12148 19556 12152 19612
rect 12152 19556 12208 19612
rect 12208 19556 12212 19612
rect 12148 19552 12212 19556
rect 12228 19612 12292 19616
rect 12228 19556 12232 19612
rect 12232 19556 12288 19612
rect 12288 19556 12292 19612
rect 12228 19552 12292 19556
rect 12308 19612 12372 19616
rect 12308 19556 12312 19612
rect 12312 19556 12368 19612
rect 12368 19556 12372 19612
rect 12308 19552 12372 19556
rect 12388 19612 12452 19616
rect 12388 19556 12392 19612
rect 12392 19556 12448 19612
rect 12448 19556 12452 19612
rect 12388 19552 12452 19556
rect 19612 19612 19676 19616
rect 19612 19556 19616 19612
rect 19616 19556 19672 19612
rect 19672 19556 19676 19612
rect 19612 19552 19676 19556
rect 19692 19612 19756 19616
rect 19692 19556 19696 19612
rect 19696 19556 19752 19612
rect 19752 19556 19756 19612
rect 19692 19552 19756 19556
rect 19772 19612 19836 19616
rect 19772 19556 19776 19612
rect 19776 19556 19832 19612
rect 19832 19556 19836 19612
rect 19772 19552 19836 19556
rect 19852 19612 19916 19616
rect 19852 19556 19856 19612
rect 19856 19556 19912 19612
rect 19912 19556 19916 19612
rect 19852 19552 19916 19556
rect 8416 19068 8480 19072
rect 8416 19012 8420 19068
rect 8420 19012 8476 19068
rect 8476 19012 8480 19068
rect 8416 19008 8480 19012
rect 8496 19068 8560 19072
rect 8496 19012 8500 19068
rect 8500 19012 8556 19068
rect 8556 19012 8560 19068
rect 8496 19008 8560 19012
rect 8576 19068 8640 19072
rect 8576 19012 8580 19068
rect 8580 19012 8636 19068
rect 8636 19012 8640 19068
rect 8576 19008 8640 19012
rect 8656 19068 8720 19072
rect 8656 19012 8660 19068
rect 8660 19012 8716 19068
rect 8716 19012 8720 19068
rect 8656 19008 8720 19012
rect 15880 19068 15944 19072
rect 15880 19012 15884 19068
rect 15884 19012 15940 19068
rect 15940 19012 15944 19068
rect 15880 19008 15944 19012
rect 15960 19068 16024 19072
rect 15960 19012 15964 19068
rect 15964 19012 16020 19068
rect 16020 19012 16024 19068
rect 15960 19008 16024 19012
rect 16040 19068 16104 19072
rect 16040 19012 16044 19068
rect 16044 19012 16100 19068
rect 16100 19012 16104 19068
rect 16040 19008 16104 19012
rect 16120 19068 16184 19072
rect 16120 19012 16124 19068
rect 16124 19012 16180 19068
rect 16180 19012 16184 19068
rect 16120 19008 16184 19012
rect 4684 18524 4748 18528
rect 4684 18468 4688 18524
rect 4688 18468 4744 18524
rect 4744 18468 4748 18524
rect 4684 18464 4748 18468
rect 4764 18524 4828 18528
rect 4764 18468 4768 18524
rect 4768 18468 4824 18524
rect 4824 18468 4828 18524
rect 4764 18464 4828 18468
rect 4844 18524 4908 18528
rect 4844 18468 4848 18524
rect 4848 18468 4904 18524
rect 4904 18468 4908 18524
rect 4844 18464 4908 18468
rect 4924 18524 4988 18528
rect 4924 18468 4928 18524
rect 4928 18468 4984 18524
rect 4984 18468 4988 18524
rect 4924 18464 4988 18468
rect 12148 18524 12212 18528
rect 12148 18468 12152 18524
rect 12152 18468 12208 18524
rect 12208 18468 12212 18524
rect 12148 18464 12212 18468
rect 12228 18524 12292 18528
rect 12228 18468 12232 18524
rect 12232 18468 12288 18524
rect 12288 18468 12292 18524
rect 12228 18464 12292 18468
rect 12308 18524 12372 18528
rect 12308 18468 12312 18524
rect 12312 18468 12368 18524
rect 12368 18468 12372 18524
rect 12308 18464 12372 18468
rect 12388 18524 12452 18528
rect 12388 18468 12392 18524
rect 12392 18468 12448 18524
rect 12448 18468 12452 18524
rect 12388 18464 12452 18468
rect 19612 18524 19676 18528
rect 19612 18468 19616 18524
rect 19616 18468 19672 18524
rect 19672 18468 19676 18524
rect 19612 18464 19676 18468
rect 19692 18524 19756 18528
rect 19692 18468 19696 18524
rect 19696 18468 19752 18524
rect 19752 18468 19756 18524
rect 19692 18464 19756 18468
rect 19772 18524 19836 18528
rect 19772 18468 19776 18524
rect 19776 18468 19832 18524
rect 19832 18468 19836 18524
rect 19772 18464 19836 18468
rect 19852 18524 19916 18528
rect 19852 18468 19856 18524
rect 19856 18468 19912 18524
rect 19912 18468 19916 18524
rect 19852 18464 19916 18468
rect 8416 17980 8480 17984
rect 8416 17924 8420 17980
rect 8420 17924 8476 17980
rect 8476 17924 8480 17980
rect 8416 17920 8480 17924
rect 8496 17980 8560 17984
rect 8496 17924 8500 17980
rect 8500 17924 8556 17980
rect 8556 17924 8560 17980
rect 8496 17920 8560 17924
rect 8576 17980 8640 17984
rect 8576 17924 8580 17980
rect 8580 17924 8636 17980
rect 8636 17924 8640 17980
rect 8576 17920 8640 17924
rect 8656 17980 8720 17984
rect 8656 17924 8660 17980
rect 8660 17924 8716 17980
rect 8716 17924 8720 17980
rect 8656 17920 8720 17924
rect 15880 17980 15944 17984
rect 15880 17924 15884 17980
rect 15884 17924 15940 17980
rect 15940 17924 15944 17980
rect 15880 17920 15944 17924
rect 15960 17980 16024 17984
rect 15960 17924 15964 17980
rect 15964 17924 16020 17980
rect 16020 17924 16024 17980
rect 15960 17920 16024 17924
rect 16040 17980 16104 17984
rect 16040 17924 16044 17980
rect 16044 17924 16100 17980
rect 16100 17924 16104 17980
rect 16040 17920 16104 17924
rect 16120 17980 16184 17984
rect 16120 17924 16124 17980
rect 16124 17924 16180 17980
rect 16180 17924 16184 17980
rect 16120 17920 16184 17924
rect 4684 17436 4748 17440
rect 4684 17380 4688 17436
rect 4688 17380 4744 17436
rect 4744 17380 4748 17436
rect 4684 17376 4748 17380
rect 4764 17436 4828 17440
rect 4764 17380 4768 17436
rect 4768 17380 4824 17436
rect 4824 17380 4828 17436
rect 4764 17376 4828 17380
rect 4844 17436 4908 17440
rect 4844 17380 4848 17436
rect 4848 17380 4904 17436
rect 4904 17380 4908 17436
rect 4844 17376 4908 17380
rect 4924 17436 4988 17440
rect 4924 17380 4928 17436
rect 4928 17380 4984 17436
rect 4984 17380 4988 17436
rect 4924 17376 4988 17380
rect 12148 17436 12212 17440
rect 12148 17380 12152 17436
rect 12152 17380 12208 17436
rect 12208 17380 12212 17436
rect 12148 17376 12212 17380
rect 12228 17436 12292 17440
rect 12228 17380 12232 17436
rect 12232 17380 12288 17436
rect 12288 17380 12292 17436
rect 12228 17376 12292 17380
rect 12308 17436 12372 17440
rect 12308 17380 12312 17436
rect 12312 17380 12368 17436
rect 12368 17380 12372 17436
rect 12308 17376 12372 17380
rect 12388 17436 12452 17440
rect 12388 17380 12392 17436
rect 12392 17380 12448 17436
rect 12448 17380 12452 17436
rect 12388 17376 12452 17380
rect 19612 17436 19676 17440
rect 19612 17380 19616 17436
rect 19616 17380 19672 17436
rect 19672 17380 19676 17436
rect 19612 17376 19676 17380
rect 19692 17436 19756 17440
rect 19692 17380 19696 17436
rect 19696 17380 19752 17436
rect 19752 17380 19756 17436
rect 19692 17376 19756 17380
rect 19772 17436 19836 17440
rect 19772 17380 19776 17436
rect 19776 17380 19832 17436
rect 19832 17380 19836 17436
rect 19772 17376 19836 17380
rect 19852 17436 19916 17440
rect 19852 17380 19856 17436
rect 19856 17380 19912 17436
rect 19912 17380 19916 17436
rect 19852 17376 19916 17380
rect 8416 16892 8480 16896
rect 8416 16836 8420 16892
rect 8420 16836 8476 16892
rect 8476 16836 8480 16892
rect 8416 16832 8480 16836
rect 8496 16892 8560 16896
rect 8496 16836 8500 16892
rect 8500 16836 8556 16892
rect 8556 16836 8560 16892
rect 8496 16832 8560 16836
rect 8576 16892 8640 16896
rect 8576 16836 8580 16892
rect 8580 16836 8636 16892
rect 8636 16836 8640 16892
rect 8576 16832 8640 16836
rect 8656 16892 8720 16896
rect 8656 16836 8660 16892
rect 8660 16836 8716 16892
rect 8716 16836 8720 16892
rect 8656 16832 8720 16836
rect 15880 16892 15944 16896
rect 15880 16836 15884 16892
rect 15884 16836 15940 16892
rect 15940 16836 15944 16892
rect 15880 16832 15944 16836
rect 15960 16892 16024 16896
rect 15960 16836 15964 16892
rect 15964 16836 16020 16892
rect 16020 16836 16024 16892
rect 15960 16832 16024 16836
rect 16040 16892 16104 16896
rect 16040 16836 16044 16892
rect 16044 16836 16100 16892
rect 16100 16836 16104 16892
rect 16040 16832 16104 16836
rect 16120 16892 16184 16896
rect 16120 16836 16124 16892
rect 16124 16836 16180 16892
rect 16180 16836 16184 16892
rect 16120 16832 16184 16836
rect 4684 16348 4748 16352
rect 4684 16292 4688 16348
rect 4688 16292 4744 16348
rect 4744 16292 4748 16348
rect 4684 16288 4748 16292
rect 4764 16348 4828 16352
rect 4764 16292 4768 16348
rect 4768 16292 4824 16348
rect 4824 16292 4828 16348
rect 4764 16288 4828 16292
rect 4844 16348 4908 16352
rect 4844 16292 4848 16348
rect 4848 16292 4904 16348
rect 4904 16292 4908 16348
rect 4844 16288 4908 16292
rect 4924 16348 4988 16352
rect 4924 16292 4928 16348
rect 4928 16292 4984 16348
rect 4984 16292 4988 16348
rect 4924 16288 4988 16292
rect 12148 16348 12212 16352
rect 12148 16292 12152 16348
rect 12152 16292 12208 16348
rect 12208 16292 12212 16348
rect 12148 16288 12212 16292
rect 12228 16348 12292 16352
rect 12228 16292 12232 16348
rect 12232 16292 12288 16348
rect 12288 16292 12292 16348
rect 12228 16288 12292 16292
rect 12308 16348 12372 16352
rect 12308 16292 12312 16348
rect 12312 16292 12368 16348
rect 12368 16292 12372 16348
rect 12308 16288 12372 16292
rect 12388 16348 12452 16352
rect 12388 16292 12392 16348
rect 12392 16292 12448 16348
rect 12448 16292 12452 16348
rect 12388 16288 12452 16292
rect 19612 16348 19676 16352
rect 19612 16292 19616 16348
rect 19616 16292 19672 16348
rect 19672 16292 19676 16348
rect 19612 16288 19676 16292
rect 19692 16348 19756 16352
rect 19692 16292 19696 16348
rect 19696 16292 19752 16348
rect 19752 16292 19756 16348
rect 19692 16288 19756 16292
rect 19772 16348 19836 16352
rect 19772 16292 19776 16348
rect 19776 16292 19832 16348
rect 19832 16292 19836 16348
rect 19772 16288 19836 16292
rect 19852 16348 19916 16352
rect 19852 16292 19856 16348
rect 19856 16292 19912 16348
rect 19912 16292 19916 16348
rect 19852 16288 19916 16292
rect 8416 15804 8480 15808
rect 8416 15748 8420 15804
rect 8420 15748 8476 15804
rect 8476 15748 8480 15804
rect 8416 15744 8480 15748
rect 8496 15804 8560 15808
rect 8496 15748 8500 15804
rect 8500 15748 8556 15804
rect 8556 15748 8560 15804
rect 8496 15744 8560 15748
rect 8576 15804 8640 15808
rect 8576 15748 8580 15804
rect 8580 15748 8636 15804
rect 8636 15748 8640 15804
rect 8576 15744 8640 15748
rect 8656 15804 8720 15808
rect 8656 15748 8660 15804
rect 8660 15748 8716 15804
rect 8716 15748 8720 15804
rect 8656 15744 8720 15748
rect 15880 15804 15944 15808
rect 15880 15748 15884 15804
rect 15884 15748 15940 15804
rect 15940 15748 15944 15804
rect 15880 15744 15944 15748
rect 15960 15804 16024 15808
rect 15960 15748 15964 15804
rect 15964 15748 16020 15804
rect 16020 15748 16024 15804
rect 15960 15744 16024 15748
rect 16040 15804 16104 15808
rect 16040 15748 16044 15804
rect 16044 15748 16100 15804
rect 16100 15748 16104 15804
rect 16040 15744 16104 15748
rect 16120 15804 16184 15808
rect 16120 15748 16124 15804
rect 16124 15748 16180 15804
rect 16180 15748 16184 15804
rect 16120 15744 16184 15748
rect 4684 15260 4748 15264
rect 4684 15204 4688 15260
rect 4688 15204 4744 15260
rect 4744 15204 4748 15260
rect 4684 15200 4748 15204
rect 4764 15260 4828 15264
rect 4764 15204 4768 15260
rect 4768 15204 4824 15260
rect 4824 15204 4828 15260
rect 4764 15200 4828 15204
rect 4844 15260 4908 15264
rect 4844 15204 4848 15260
rect 4848 15204 4904 15260
rect 4904 15204 4908 15260
rect 4844 15200 4908 15204
rect 4924 15260 4988 15264
rect 4924 15204 4928 15260
rect 4928 15204 4984 15260
rect 4984 15204 4988 15260
rect 4924 15200 4988 15204
rect 12148 15260 12212 15264
rect 12148 15204 12152 15260
rect 12152 15204 12208 15260
rect 12208 15204 12212 15260
rect 12148 15200 12212 15204
rect 12228 15260 12292 15264
rect 12228 15204 12232 15260
rect 12232 15204 12288 15260
rect 12288 15204 12292 15260
rect 12228 15200 12292 15204
rect 12308 15260 12372 15264
rect 12308 15204 12312 15260
rect 12312 15204 12368 15260
rect 12368 15204 12372 15260
rect 12308 15200 12372 15204
rect 12388 15260 12452 15264
rect 12388 15204 12392 15260
rect 12392 15204 12448 15260
rect 12448 15204 12452 15260
rect 12388 15200 12452 15204
rect 19612 15260 19676 15264
rect 19612 15204 19616 15260
rect 19616 15204 19672 15260
rect 19672 15204 19676 15260
rect 19612 15200 19676 15204
rect 19692 15260 19756 15264
rect 19692 15204 19696 15260
rect 19696 15204 19752 15260
rect 19752 15204 19756 15260
rect 19692 15200 19756 15204
rect 19772 15260 19836 15264
rect 19772 15204 19776 15260
rect 19776 15204 19832 15260
rect 19832 15204 19836 15260
rect 19772 15200 19836 15204
rect 19852 15260 19916 15264
rect 19852 15204 19856 15260
rect 19856 15204 19912 15260
rect 19912 15204 19916 15260
rect 19852 15200 19916 15204
rect 8416 14716 8480 14720
rect 8416 14660 8420 14716
rect 8420 14660 8476 14716
rect 8476 14660 8480 14716
rect 8416 14656 8480 14660
rect 8496 14716 8560 14720
rect 8496 14660 8500 14716
rect 8500 14660 8556 14716
rect 8556 14660 8560 14716
rect 8496 14656 8560 14660
rect 8576 14716 8640 14720
rect 8576 14660 8580 14716
rect 8580 14660 8636 14716
rect 8636 14660 8640 14716
rect 8576 14656 8640 14660
rect 8656 14716 8720 14720
rect 8656 14660 8660 14716
rect 8660 14660 8716 14716
rect 8716 14660 8720 14716
rect 8656 14656 8720 14660
rect 15880 14716 15944 14720
rect 15880 14660 15884 14716
rect 15884 14660 15940 14716
rect 15940 14660 15944 14716
rect 15880 14656 15944 14660
rect 15960 14716 16024 14720
rect 15960 14660 15964 14716
rect 15964 14660 16020 14716
rect 16020 14660 16024 14716
rect 15960 14656 16024 14660
rect 16040 14716 16104 14720
rect 16040 14660 16044 14716
rect 16044 14660 16100 14716
rect 16100 14660 16104 14716
rect 16040 14656 16104 14660
rect 16120 14716 16184 14720
rect 16120 14660 16124 14716
rect 16124 14660 16180 14716
rect 16180 14660 16184 14716
rect 16120 14656 16184 14660
rect 4684 14172 4748 14176
rect 4684 14116 4688 14172
rect 4688 14116 4744 14172
rect 4744 14116 4748 14172
rect 4684 14112 4748 14116
rect 4764 14172 4828 14176
rect 4764 14116 4768 14172
rect 4768 14116 4824 14172
rect 4824 14116 4828 14172
rect 4764 14112 4828 14116
rect 4844 14172 4908 14176
rect 4844 14116 4848 14172
rect 4848 14116 4904 14172
rect 4904 14116 4908 14172
rect 4844 14112 4908 14116
rect 4924 14172 4988 14176
rect 4924 14116 4928 14172
rect 4928 14116 4984 14172
rect 4984 14116 4988 14172
rect 4924 14112 4988 14116
rect 12148 14172 12212 14176
rect 12148 14116 12152 14172
rect 12152 14116 12208 14172
rect 12208 14116 12212 14172
rect 12148 14112 12212 14116
rect 12228 14172 12292 14176
rect 12228 14116 12232 14172
rect 12232 14116 12288 14172
rect 12288 14116 12292 14172
rect 12228 14112 12292 14116
rect 12308 14172 12372 14176
rect 12308 14116 12312 14172
rect 12312 14116 12368 14172
rect 12368 14116 12372 14172
rect 12308 14112 12372 14116
rect 12388 14172 12452 14176
rect 12388 14116 12392 14172
rect 12392 14116 12448 14172
rect 12448 14116 12452 14172
rect 12388 14112 12452 14116
rect 19612 14172 19676 14176
rect 19612 14116 19616 14172
rect 19616 14116 19672 14172
rect 19672 14116 19676 14172
rect 19612 14112 19676 14116
rect 19692 14172 19756 14176
rect 19692 14116 19696 14172
rect 19696 14116 19752 14172
rect 19752 14116 19756 14172
rect 19692 14112 19756 14116
rect 19772 14172 19836 14176
rect 19772 14116 19776 14172
rect 19776 14116 19832 14172
rect 19832 14116 19836 14172
rect 19772 14112 19836 14116
rect 19852 14172 19916 14176
rect 19852 14116 19856 14172
rect 19856 14116 19912 14172
rect 19912 14116 19916 14172
rect 19852 14112 19916 14116
rect 8416 13628 8480 13632
rect 8416 13572 8420 13628
rect 8420 13572 8476 13628
rect 8476 13572 8480 13628
rect 8416 13568 8480 13572
rect 8496 13628 8560 13632
rect 8496 13572 8500 13628
rect 8500 13572 8556 13628
rect 8556 13572 8560 13628
rect 8496 13568 8560 13572
rect 8576 13628 8640 13632
rect 8576 13572 8580 13628
rect 8580 13572 8636 13628
rect 8636 13572 8640 13628
rect 8576 13568 8640 13572
rect 8656 13628 8720 13632
rect 8656 13572 8660 13628
rect 8660 13572 8716 13628
rect 8716 13572 8720 13628
rect 8656 13568 8720 13572
rect 15880 13628 15944 13632
rect 15880 13572 15884 13628
rect 15884 13572 15940 13628
rect 15940 13572 15944 13628
rect 15880 13568 15944 13572
rect 15960 13628 16024 13632
rect 15960 13572 15964 13628
rect 15964 13572 16020 13628
rect 16020 13572 16024 13628
rect 15960 13568 16024 13572
rect 16040 13628 16104 13632
rect 16040 13572 16044 13628
rect 16044 13572 16100 13628
rect 16100 13572 16104 13628
rect 16040 13568 16104 13572
rect 16120 13628 16184 13632
rect 16120 13572 16124 13628
rect 16124 13572 16180 13628
rect 16180 13572 16184 13628
rect 16120 13568 16184 13572
rect 4684 13084 4748 13088
rect 4684 13028 4688 13084
rect 4688 13028 4744 13084
rect 4744 13028 4748 13084
rect 4684 13024 4748 13028
rect 4764 13084 4828 13088
rect 4764 13028 4768 13084
rect 4768 13028 4824 13084
rect 4824 13028 4828 13084
rect 4764 13024 4828 13028
rect 4844 13084 4908 13088
rect 4844 13028 4848 13084
rect 4848 13028 4904 13084
rect 4904 13028 4908 13084
rect 4844 13024 4908 13028
rect 4924 13084 4988 13088
rect 4924 13028 4928 13084
rect 4928 13028 4984 13084
rect 4984 13028 4988 13084
rect 4924 13024 4988 13028
rect 12148 13084 12212 13088
rect 12148 13028 12152 13084
rect 12152 13028 12208 13084
rect 12208 13028 12212 13084
rect 12148 13024 12212 13028
rect 12228 13084 12292 13088
rect 12228 13028 12232 13084
rect 12232 13028 12288 13084
rect 12288 13028 12292 13084
rect 12228 13024 12292 13028
rect 12308 13084 12372 13088
rect 12308 13028 12312 13084
rect 12312 13028 12368 13084
rect 12368 13028 12372 13084
rect 12308 13024 12372 13028
rect 12388 13084 12452 13088
rect 12388 13028 12392 13084
rect 12392 13028 12448 13084
rect 12448 13028 12452 13084
rect 12388 13024 12452 13028
rect 19612 13084 19676 13088
rect 19612 13028 19616 13084
rect 19616 13028 19672 13084
rect 19672 13028 19676 13084
rect 19612 13024 19676 13028
rect 19692 13084 19756 13088
rect 19692 13028 19696 13084
rect 19696 13028 19752 13084
rect 19752 13028 19756 13084
rect 19692 13024 19756 13028
rect 19772 13084 19836 13088
rect 19772 13028 19776 13084
rect 19776 13028 19832 13084
rect 19832 13028 19836 13084
rect 19772 13024 19836 13028
rect 19852 13084 19916 13088
rect 19852 13028 19856 13084
rect 19856 13028 19912 13084
rect 19912 13028 19916 13084
rect 19852 13024 19916 13028
rect 8416 12540 8480 12544
rect 8416 12484 8420 12540
rect 8420 12484 8476 12540
rect 8476 12484 8480 12540
rect 8416 12480 8480 12484
rect 8496 12540 8560 12544
rect 8496 12484 8500 12540
rect 8500 12484 8556 12540
rect 8556 12484 8560 12540
rect 8496 12480 8560 12484
rect 8576 12540 8640 12544
rect 8576 12484 8580 12540
rect 8580 12484 8636 12540
rect 8636 12484 8640 12540
rect 8576 12480 8640 12484
rect 8656 12540 8720 12544
rect 8656 12484 8660 12540
rect 8660 12484 8716 12540
rect 8716 12484 8720 12540
rect 8656 12480 8720 12484
rect 15880 12540 15944 12544
rect 15880 12484 15884 12540
rect 15884 12484 15940 12540
rect 15940 12484 15944 12540
rect 15880 12480 15944 12484
rect 15960 12540 16024 12544
rect 15960 12484 15964 12540
rect 15964 12484 16020 12540
rect 16020 12484 16024 12540
rect 15960 12480 16024 12484
rect 16040 12540 16104 12544
rect 16040 12484 16044 12540
rect 16044 12484 16100 12540
rect 16100 12484 16104 12540
rect 16040 12480 16104 12484
rect 16120 12540 16184 12544
rect 16120 12484 16124 12540
rect 16124 12484 16180 12540
rect 16180 12484 16184 12540
rect 16120 12480 16184 12484
rect 4684 11996 4748 12000
rect 4684 11940 4688 11996
rect 4688 11940 4744 11996
rect 4744 11940 4748 11996
rect 4684 11936 4748 11940
rect 4764 11996 4828 12000
rect 4764 11940 4768 11996
rect 4768 11940 4824 11996
rect 4824 11940 4828 11996
rect 4764 11936 4828 11940
rect 4844 11996 4908 12000
rect 4844 11940 4848 11996
rect 4848 11940 4904 11996
rect 4904 11940 4908 11996
rect 4844 11936 4908 11940
rect 4924 11996 4988 12000
rect 4924 11940 4928 11996
rect 4928 11940 4984 11996
rect 4984 11940 4988 11996
rect 4924 11936 4988 11940
rect 12148 11996 12212 12000
rect 12148 11940 12152 11996
rect 12152 11940 12208 11996
rect 12208 11940 12212 11996
rect 12148 11936 12212 11940
rect 12228 11996 12292 12000
rect 12228 11940 12232 11996
rect 12232 11940 12288 11996
rect 12288 11940 12292 11996
rect 12228 11936 12292 11940
rect 12308 11996 12372 12000
rect 12308 11940 12312 11996
rect 12312 11940 12368 11996
rect 12368 11940 12372 11996
rect 12308 11936 12372 11940
rect 12388 11996 12452 12000
rect 12388 11940 12392 11996
rect 12392 11940 12448 11996
rect 12448 11940 12452 11996
rect 12388 11936 12452 11940
rect 19612 11996 19676 12000
rect 19612 11940 19616 11996
rect 19616 11940 19672 11996
rect 19672 11940 19676 11996
rect 19612 11936 19676 11940
rect 19692 11996 19756 12000
rect 19692 11940 19696 11996
rect 19696 11940 19752 11996
rect 19752 11940 19756 11996
rect 19692 11936 19756 11940
rect 19772 11996 19836 12000
rect 19772 11940 19776 11996
rect 19776 11940 19832 11996
rect 19832 11940 19836 11996
rect 19772 11936 19836 11940
rect 19852 11996 19916 12000
rect 19852 11940 19856 11996
rect 19856 11940 19912 11996
rect 19912 11940 19916 11996
rect 19852 11936 19916 11940
rect 8416 11452 8480 11456
rect 8416 11396 8420 11452
rect 8420 11396 8476 11452
rect 8476 11396 8480 11452
rect 8416 11392 8480 11396
rect 8496 11452 8560 11456
rect 8496 11396 8500 11452
rect 8500 11396 8556 11452
rect 8556 11396 8560 11452
rect 8496 11392 8560 11396
rect 8576 11452 8640 11456
rect 8576 11396 8580 11452
rect 8580 11396 8636 11452
rect 8636 11396 8640 11452
rect 8576 11392 8640 11396
rect 8656 11452 8720 11456
rect 8656 11396 8660 11452
rect 8660 11396 8716 11452
rect 8716 11396 8720 11452
rect 8656 11392 8720 11396
rect 15880 11452 15944 11456
rect 15880 11396 15884 11452
rect 15884 11396 15940 11452
rect 15940 11396 15944 11452
rect 15880 11392 15944 11396
rect 15960 11452 16024 11456
rect 15960 11396 15964 11452
rect 15964 11396 16020 11452
rect 16020 11396 16024 11452
rect 15960 11392 16024 11396
rect 16040 11452 16104 11456
rect 16040 11396 16044 11452
rect 16044 11396 16100 11452
rect 16100 11396 16104 11452
rect 16040 11392 16104 11396
rect 16120 11452 16184 11456
rect 16120 11396 16124 11452
rect 16124 11396 16180 11452
rect 16180 11396 16184 11452
rect 16120 11392 16184 11396
rect 4684 10908 4748 10912
rect 4684 10852 4688 10908
rect 4688 10852 4744 10908
rect 4744 10852 4748 10908
rect 4684 10848 4748 10852
rect 4764 10908 4828 10912
rect 4764 10852 4768 10908
rect 4768 10852 4824 10908
rect 4824 10852 4828 10908
rect 4764 10848 4828 10852
rect 4844 10908 4908 10912
rect 4844 10852 4848 10908
rect 4848 10852 4904 10908
rect 4904 10852 4908 10908
rect 4844 10848 4908 10852
rect 4924 10908 4988 10912
rect 4924 10852 4928 10908
rect 4928 10852 4984 10908
rect 4984 10852 4988 10908
rect 4924 10848 4988 10852
rect 12148 10908 12212 10912
rect 12148 10852 12152 10908
rect 12152 10852 12208 10908
rect 12208 10852 12212 10908
rect 12148 10848 12212 10852
rect 12228 10908 12292 10912
rect 12228 10852 12232 10908
rect 12232 10852 12288 10908
rect 12288 10852 12292 10908
rect 12228 10848 12292 10852
rect 12308 10908 12372 10912
rect 12308 10852 12312 10908
rect 12312 10852 12368 10908
rect 12368 10852 12372 10908
rect 12308 10848 12372 10852
rect 12388 10908 12452 10912
rect 12388 10852 12392 10908
rect 12392 10852 12448 10908
rect 12448 10852 12452 10908
rect 12388 10848 12452 10852
rect 19612 10908 19676 10912
rect 19612 10852 19616 10908
rect 19616 10852 19672 10908
rect 19672 10852 19676 10908
rect 19612 10848 19676 10852
rect 19692 10908 19756 10912
rect 19692 10852 19696 10908
rect 19696 10852 19752 10908
rect 19752 10852 19756 10908
rect 19692 10848 19756 10852
rect 19772 10908 19836 10912
rect 19772 10852 19776 10908
rect 19776 10852 19832 10908
rect 19832 10852 19836 10908
rect 19772 10848 19836 10852
rect 19852 10908 19916 10912
rect 19852 10852 19856 10908
rect 19856 10852 19912 10908
rect 19912 10852 19916 10908
rect 19852 10848 19916 10852
rect 8416 10364 8480 10368
rect 8416 10308 8420 10364
rect 8420 10308 8476 10364
rect 8476 10308 8480 10364
rect 8416 10304 8480 10308
rect 8496 10364 8560 10368
rect 8496 10308 8500 10364
rect 8500 10308 8556 10364
rect 8556 10308 8560 10364
rect 8496 10304 8560 10308
rect 8576 10364 8640 10368
rect 8576 10308 8580 10364
rect 8580 10308 8636 10364
rect 8636 10308 8640 10364
rect 8576 10304 8640 10308
rect 8656 10364 8720 10368
rect 8656 10308 8660 10364
rect 8660 10308 8716 10364
rect 8716 10308 8720 10364
rect 8656 10304 8720 10308
rect 15880 10364 15944 10368
rect 15880 10308 15884 10364
rect 15884 10308 15940 10364
rect 15940 10308 15944 10364
rect 15880 10304 15944 10308
rect 15960 10364 16024 10368
rect 15960 10308 15964 10364
rect 15964 10308 16020 10364
rect 16020 10308 16024 10364
rect 15960 10304 16024 10308
rect 16040 10364 16104 10368
rect 16040 10308 16044 10364
rect 16044 10308 16100 10364
rect 16100 10308 16104 10364
rect 16040 10304 16104 10308
rect 16120 10364 16184 10368
rect 16120 10308 16124 10364
rect 16124 10308 16180 10364
rect 16180 10308 16184 10364
rect 16120 10304 16184 10308
rect 4684 9820 4748 9824
rect 4684 9764 4688 9820
rect 4688 9764 4744 9820
rect 4744 9764 4748 9820
rect 4684 9760 4748 9764
rect 4764 9820 4828 9824
rect 4764 9764 4768 9820
rect 4768 9764 4824 9820
rect 4824 9764 4828 9820
rect 4764 9760 4828 9764
rect 4844 9820 4908 9824
rect 4844 9764 4848 9820
rect 4848 9764 4904 9820
rect 4904 9764 4908 9820
rect 4844 9760 4908 9764
rect 4924 9820 4988 9824
rect 4924 9764 4928 9820
rect 4928 9764 4984 9820
rect 4984 9764 4988 9820
rect 4924 9760 4988 9764
rect 12148 9820 12212 9824
rect 12148 9764 12152 9820
rect 12152 9764 12208 9820
rect 12208 9764 12212 9820
rect 12148 9760 12212 9764
rect 12228 9820 12292 9824
rect 12228 9764 12232 9820
rect 12232 9764 12288 9820
rect 12288 9764 12292 9820
rect 12228 9760 12292 9764
rect 12308 9820 12372 9824
rect 12308 9764 12312 9820
rect 12312 9764 12368 9820
rect 12368 9764 12372 9820
rect 12308 9760 12372 9764
rect 12388 9820 12452 9824
rect 12388 9764 12392 9820
rect 12392 9764 12448 9820
rect 12448 9764 12452 9820
rect 12388 9760 12452 9764
rect 19612 9820 19676 9824
rect 19612 9764 19616 9820
rect 19616 9764 19672 9820
rect 19672 9764 19676 9820
rect 19612 9760 19676 9764
rect 19692 9820 19756 9824
rect 19692 9764 19696 9820
rect 19696 9764 19752 9820
rect 19752 9764 19756 9820
rect 19692 9760 19756 9764
rect 19772 9820 19836 9824
rect 19772 9764 19776 9820
rect 19776 9764 19832 9820
rect 19832 9764 19836 9820
rect 19772 9760 19836 9764
rect 19852 9820 19916 9824
rect 19852 9764 19856 9820
rect 19856 9764 19912 9820
rect 19912 9764 19916 9820
rect 19852 9760 19916 9764
rect 8416 9276 8480 9280
rect 8416 9220 8420 9276
rect 8420 9220 8476 9276
rect 8476 9220 8480 9276
rect 8416 9216 8480 9220
rect 8496 9276 8560 9280
rect 8496 9220 8500 9276
rect 8500 9220 8556 9276
rect 8556 9220 8560 9276
rect 8496 9216 8560 9220
rect 8576 9276 8640 9280
rect 8576 9220 8580 9276
rect 8580 9220 8636 9276
rect 8636 9220 8640 9276
rect 8576 9216 8640 9220
rect 8656 9276 8720 9280
rect 8656 9220 8660 9276
rect 8660 9220 8716 9276
rect 8716 9220 8720 9276
rect 8656 9216 8720 9220
rect 15880 9276 15944 9280
rect 15880 9220 15884 9276
rect 15884 9220 15940 9276
rect 15940 9220 15944 9276
rect 15880 9216 15944 9220
rect 15960 9276 16024 9280
rect 15960 9220 15964 9276
rect 15964 9220 16020 9276
rect 16020 9220 16024 9276
rect 15960 9216 16024 9220
rect 16040 9276 16104 9280
rect 16040 9220 16044 9276
rect 16044 9220 16100 9276
rect 16100 9220 16104 9276
rect 16040 9216 16104 9220
rect 16120 9276 16184 9280
rect 16120 9220 16124 9276
rect 16124 9220 16180 9276
rect 16180 9220 16184 9276
rect 16120 9216 16184 9220
rect 19380 9148 19444 9212
rect 4684 8732 4748 8736
rect 4684 8676 4688 8732
rect 4688 8676 4744 8732
rect 4744 8676 4748 8732
rect 4684 8672 4748 8676
rect 4764 8732 4828 8736
rect 4764 8676 4768 8732
rect 4768 8676 4824 8732
rect 4824 8676 4828 8732
rect 4764 8672 4828 8676
rect 4844 8732 4908 8736
rect 4844 8676 4848 8732
rect 4848 8676 4904 8732
rect 4904 8676 4908 8732
rect 4844 8672 4908 8676
rect 4924 8732 4988 8736
rect 4924 8676 4928 8732
rect 4928 8676 4984 8732
rect 4984 8676 4988 8732
rect 4924 8672 4988 8676
rect 12148 8732 12212 8736
rect 12148 8676 12152 8732
rect 12152 8676 12208 8732
rect 12208 8676 12212 8732
rect 12148 8672 12212 8676
rect 12228 8732 12292 8736
rect 12228 8676 12232 8732
rect 12232 8676 12288 8732
rect 12288 8676 12292 8732
rect 12228 8672 12292 8676
rect 12308 8732 12372 8736
rect 12308 8676 12312 8732
rect 12312 8676 12368 8732
rect 12368 8676 12372 8732
rect 12308 8672 12372 8676
rect 12388 8732 12452 8736
rect 12388 8676 12392 8732
rect 12392 8676 12448 8732
rect 12448 8676 12452 8732
rect 12388 8672 12452 8676
rect 19612 8732 19676 8736
rect 19612 8676 19616 8732
rect 19616 8676 19672 8732
rect 19672 8676 19676 8732
rect 19612 8672 19676 8676
rect 19692 8732 19756 8736
rect 19692 8676 19696 8732
rect 19696 8676 19752 8732
rect 19752 8676 19756 8732
rect 19692 8672 19756 8676
rect 19772 8732 19836 8736
rect 19772 8676 19776 8732
rect 19776 8676 19832 8732
rect 19832 8676 19836 8732
rect 19772 8672 19836 8676
rect 19852 8732 19916 8736
rect 19852 8676 19856 8732
rect 19856 8676 19912 8732
rect 19912 8676 19916 8732
rect 19852 8672 19916 8676
rect 19380 8392 19444 8396
rect 19380 8336 19394 8392
rect 19394 8336 19444 8392
rect 19380 8332 19444 8336
rect 8416 8188 8480 8192
rect 8416 8132 8420 8188
rect 8420 8132 8476 8188
rect 8476 8132 8480 8188
rect 8416 8128 8480 8132
rect 8496 8188 8560 8192
rect 8496 8132 8500 8188
rect 8500 8132 8556 8188
rect 8556 8132 8560 8188
rect 8496 8128 8560 8132
rect 8576 8188 8640 8192
rect 8576 8132 8580 8188
rect 8580 8132 8636 8188
rect 8636 8132 8640 8188
rect 8576 8128 8640 8132
rect 8656 8188 8720 8192
rect 8656 8132 8660 8188
rect 8660 8132 8716 8188
rect 8716 8132 8720 8188
rect 8656 8128 8720 8132
rect 15880 8188 15944 8192
rect 15880 8132 15884 8188
rect 15884 8132 15940 8188
rect 15940 8132 15944 8188
rect 15880 8128 15944 8132
rect 15960 8188 16024 8192
rect 15960 8132 15964 8188
rect 15964 8132 16020 8188
rect 16020 8132 16024 8188
rect 15960 8128 16024 8132
rect 16040 8188 16104 8192
rect 16040 8132 16044 8188
rect 16044 8132 16100 8188
rect 16100 8132 16104 8188
rect 16040 8128 16104 8132
rect 16120 8188 16184 8192
rect 16120 8132 16124 8188
rect 16124 8132 16180 8188
rect 16180 8132 16184 8188
rect 16120 8128 16184 8132
rect 4684 7644 4748 7648
rect 4684 7588 4688 7644
rect 4688 7588 4744 7644
rect 4744 7588 4748 7644
rect 4684 7584 4748 7588
rect 4764 7644 4828 7648
rect 4764 7588 4768 7644
rect 4768 7588 4824 7644
rect 4824 7588 4828 7644
rect 4764 7584 4828 7588
rect 4844 7644 4908 7648
rect 4844 7588 4848 7644
rect 4848 7588 4904 7644
rect 4904 7588 4908 7644
rect 4844 7584 4908 7588
rect 4924 7644 4988 7648
rect 4924 7588 4928 7644
rect 4928 7588 4984 7644
rect 4984 7588 4988 7644
rect 4924 7584 4988 7588
rect 12148 7644 12212 7648
rect 12148 7588 12152 7644
rect 12152 7588 12208 7644
rect 12208 7588 12212 7644
rect 12148 7584 12212 7588
rect 12228 7644 12292 7648
rect 12228 7588 12232 7644
rect 12232 7588 12288 7644
rect 12288 7588 12292 7644
rect 12228 7584 12292 7588
rect 12308 7644 12372 7648
rect 12308 7588 12312 7644
rect 12312 7588 12368 7644
rect 12368 7588 12372 7644
rect 12308 7584 12372 7588
rect 12388 7644 12452 7648
rect 12388 7588 12392 7644
rect 12392 7588 12448 7644
rect 12448 7588 12452 7644
rect 12388 7584 12452 7588
rect 19612 7644 19676 7648
rect 19612 7588 19616 7644
rect 19616 7588 19672 7644
rect 19672 7588 19676 7644
rect 19612 7584 19676 7588
rect 19692 7644 19756 7648
rect 19692 7588 19696 7644
rect 19696 7588 19752 7644
rect 19752 7588 19756 7644
rect 19692 7584 19756 7588
rect 19772 7644 19836 7648
rect 19772 7588 19776 7644
rect 19776 7588 19832 7644
rect 19832 7588 19836 7644
rect 19772 7584 19836 7588
rect 19852 7644 19916 7648
rect 19852 7588 19856 7644
rect 19856 7588 19912 7644
rect 19912 7588 19916 7644
rect 19852 7584 19916 7588
rect 8416 7100 8480 7104
rect 8416 7044 8420 7100
rect 8420 7044 8476 7100
rect 8476 7044 8480 7100
rect 8416 7040 8480 7044
rect 8496 7100 8560 7104
rect 8496 7044 8500 7100
rect 8500 7044 8556 7100
rect 8556 7044 8560 7100
rect 8496 7040 8560 7044
rect 8576 7100 8640 7104
rect 8576 7044 8580 7100
rect 8580 7044 8636 7100
rect 8636 7044 8640 7100
rect 8576 7040 8640 7044
rect 8656 7100 8720 7104
rect 8656 7044 8660 7100
rect 8660 7044 8716 7100
rect 8716 7044 8720 7100
rect 8656 7040 8720 7044
rect 15880 7100 15944 7104
rect 15880 7044 15884 7100
rect 15884 7044 15940 7100
rect 15940 7044 15944 7100
rect 15880 7040 15944 7044
rect 15960 7100 16024 7104
rect 15960 7044 15964 7100
rect 15964 7044 16020 7100
rect 16020 7044 16024 7100
rect 15960 7040 16024 7044
rect 16040 7100 16104 7104
rect 16040 7044 16044 7100
rect 16044 7044 16100 7100
rect 16100 7044 16104 7100
rect 16040 7040 16104 7044
rect 16120 7100 16184 7104
rect 16120 7044 16124 7100
rect 16124 7044 16180 7100
rect 16180 7044 16184 7100
rect 16120 7040 16184 7044
rect 4684 6556 4748 6560
rect 4684 6500 4688 6556
rect 4688 6500 4744 6556
rect 4744 6500 4748 6556
rect 4684 6496 4748 6500
rect 4764 6556 4828 6560
rect 4764 6500 4768 6556
rect 4768 6500 4824 6556
rect 4824 6500 4828 6556
rect 4764 6496 4828 6500
rect 4844 6556 4908 6560
rect 4844 6500 4848 6556
rect 4848 6500 4904 6556
rect 4904 6500 4908 6556
rect 4844 6496 4908 6500
rect 4924 6556 4988 6560
rect 4924 6500 4928 6556
rect 4928 6500 4984 6556
rect 4984 6500 4988 6556
rect 4924 6496 4988 6500
rect 12148 6556 12212 6560
rect 12148 6500 12152 6556
rect 12152 6500 12208 6556
rect 12208 6500 12212 6556
rect 12148 6496 12212 6500
rect 12228 6556 12292 6560
rect 12228 6500 12232 6556
rect 12232 6500 12288 6556
rect 12288 6500 12292 6556
rect 12228 6496 12292 6500
rect 12308 6556 12372 6560
rect 12308 6500 12312 6556
rect 12312 6500 12368 6556
rect 12368 6500 12372 6556
rect 12308 6496 12372 6500
rect 12388 6556 12452 6560
rect 12388 6500 12392 6556
rect 12392 6500 12448 6556
rect 12448 6500 12452 6556
rect 12388 6496 12452 6500
rect 19612 6556 19676 6560
rect 19612 6500 19616 6556
rect 19616 6500 19672 6556
rect 19672 6500 19676 6556
rect 19612 6496 19676 6500
rect 19692 6556 19756 6560
rect 19692 6500 19696 6556
rect 19696 6500 19752 6556
rect 19752 6500 19756 6556
rect 19692 6496 19756 6500
rect 19772 6556 19836 6560
rect 19772 6500 19776 6556
rect 19776 6500 19832 6556
rect 19832 6500 19836 6556
rect 19772 6496 19836 6500
rect 19852 6556 19916 6560
rect 19852 6500 19856 6556
rect 19856 6500 19912 6556
rect 19912 6500 19916 6556
rect 19852 6496 19916 6500
rect 8416 6012 8480 6016
rect 8416 5956 8420 6012
rect 8420 5956 8476 6012
rect 8476 5956 8480 6012
rect 8416 5952 8480 5956
rect 8496 6012 8560 6016
rect 8496 5956 8500 6012
rect 8500 5956 8556 6012
rect 8556 5956 8560 6012
rect 8496 5952 8560 5956
rect 8576 6012 8640 6016
rect 8576 5956 8580 6012
rect 8580 5956 8636 6012
rect 8636 5956 8640 6012
rect 8576 5952 8640 5956
rect 8656 6012 8720 6016
rect 8656 5956 8660 6012
rect 8660 5956 8716 6012
rect 8716 5956 8720 6012
rect 8656 5952 8720 5956
rect 15880 6012 15944 6016
rect 15880 5956 15884 6012
rect 15884 5956 15940 6012
rect 15940 5956 15944 6012
rect 15880 5952 15944 5956
rect 15960 6012 16024 6016
rect 15960 5956 15964 6012
rect 15964 5956 16020 6012
rect 16020 5956 16024 6012
rect 15960 5952 16024 5956
rect 16040 6012 16104 6016
rect 16040 5956 16044 6012
rect 16044 5956 16100 6012
rect 16100 5956 16104 6012
rect 16040 5952 16104 5956
rect 16120 6012 16184 6016
rect 16120 5956 16124 6012
rect 16124 5956 16180 6012
rect 16180 5956 16184 6012
rect 16120 5952 16184 5956
rect 4684 5468 4748 5472
rect 4684 5412 4688 5468
rect 4688 5412 4744 5468
rect 4744 5412 4748 5468
rect 4684 5408 4748 5412
rect 4764 5468 4828 5472
rect 4764 5412 4768 5468
rect 4768 5412 4824 5468
rect 4824 5412 4828 5468
rect 4764 5408 4828 5412
rect 4844 5468 4908 5472
rect 4844 5412 4848 5468
rect 4848 5412 4904 5468
rect 4904 5412 4908 5468
rect 4844 5408 4908 5412
rect 4924 5468 4988 5472
rect 4924 5412 4928 5468
rect 4928 5412 4984 5468
rect 4984 5412 4988 5468
rect 4924 5408 4988 5412
rect 12148 5468 12212 5472
rect 12148 5412 12152 5468
rect 12152 5412 12208 5468
rect 12208 5412 12212 5468
rect 12148 5408 12212 5412
rect 12228 5468 12292 5472
rect 12228 5412 12232 5468
rect 12232 5412 12288 5468
rect 12288 5412 12292 5468
rect 12228 5408 12292 5412
rect 12308 5468 12372 5472
rect 12308 5412 12312 5468
rect 12312 5412 12368 5468
rect 12368 5412 12372 5468
rect 12308 5408 12372 5412
rect 12388 5468 12452 5472
rect 12388 5412 12392 5468
rect 12392 5412 12448 5468
rect 12448 5412 12452 5468
rect 12388 5408 12452 5412
rect 19612 5468 19676 5472
rect 19612 5412 19616 5468
rect 19616 5412 19672 5468
rect 19672 5412 19676 5468
rect 19612 5408 19676 5412
rect 19692 5468 19756 5472
rect 19692 5412 19696 5468
rect 19696 5412 19752 5468
rect 19752 5412 19756 5468
rect 19692 5408 19756 5412
rect 19772 5468 19836 5472
rect 19772 5412 19776 5468
rect 19776 5412 19832 5468
rect 19832 5412 19836 5468
rect 19772 5408 19836 5412
rect 19852 5468 19916 5472
rect 19852 5412 19856 5468
rect 19856 5412 19912 5468
rect 19912 5412 19916 5468
rect 19852 5408 19916 5412
rect 8416 4924 8480 4928
rect 8416 4868 8420 4924
rect 8420 4868 8476 4924
rect 8476 4868 8480 4924
rect 8416 4864 8480 4868
rect 8496 4924 8560 4928
rect 8496 4868 8500 4924
rect 8500 4868 8556 4924
rect 8556 4868 8560 4924
rect 8496 4864 8560 4868
rect 8576 4924 8640 4928
rect 8576 4868 8580 4924
rect 8580 4868 8636 4924
rect 8636 4868 8640 4924
rect 8576 4864 8640 4868
rect 8656 4924 8720 4928
rect 8656 4868 8660 4924
rect 8660 4868 8716 4924
rect 8716 4868 8720 4924
rect 8656 4864 8720 4868
rect 15880 4924 15944 4928
rect 15880 4868 15884 4924
rect 15884 4868 15940 4924
rect 15940 4868 15944 4924
rect 15880 4864 15944 4868
rect 15960 4924 16024 4928
rect 15960 4868 15964 4924
rect 15964 4868 16020 4924
rect 16020 4868 16024 4924
rect 15960 4864 16024 4868
rect 16040 4924 16104 4928
rect 16040 4868 16044 4924
rect 16044 4868 16100 4924
rect 16100 4868 16104 4924
rect 16040 4864 16104 4868
rect 16120 4924 16184 4928
rect 16120 4868 16124 4924
rect 16124 4868 16180 4924
rect 16180 4868 16184 4924
rect 16120 4864 16184 4868
rect 4684 4380 4748 4384
rect 4684 4324 4688 4380
rect 4688 4324 4744 4380
rect 4744 4324 4748 4380
rect 4684 4320 4748 4324
rect 4764 4380 4828 4384
rect 4764 4324 4768 4380
rect 4768 4324 4824 4380
rect 4824 4324 4828 4380
rect 4764 4320 4828 4324
rect 4844 4380 4908 4384
rect 4844 4324 4848 4380
rect 4848 4324 4904 4380
rect 4904 4324 4908 4380
rect 4844 4320 4908 4324
rect 4924 4380 4988 4384
rect 4924 4324 4928 4380
rect 4928 4324 4984 4380
rect 4984 4324 4988 4380
rect 4924 4320 4988 4324
rect 12148 4380 12212 4384
rect 12148 4324 12152 4380
rect 12152 4324 12208 4380
rect 12208 4324 12212 4380
rect 12148 4320 12212 4324
rect 12228 4380 12292 4384
rect 12228 4324 12232 4380
rect 12232 4324 12288 4380
rect 12288 4324 12292 4380
rect 12228 4320 12292 4324
rect 12308 4380 12372 4384
rect 12308 4324 12312 4380
rect 12312 4324 12368 4380
rect 12368 4324 12372 4380
rect 12308 4320 12372 4324
rect 12388 4380 12452 4384
rect 12388 4324 12392 4380
rect 12392 4324 12448 4380
rect 12448 4324 12452 4380
rect 12388 4320 12452 4324
rect 19612 4380 19676 4384
rect 19612 4324 19616 4380
rect 19616 4324 19672 4380
rect 19672 4324 19676 4380
rect 19612 4320 19676 4324
rect 19692 4380 19756 4384
rect 19692 4324 19696 4380
rect 19696 4324 19752 4380
rect 19752 4324 19756 4380
rect 19692 4320 19756 4324
rect 19772 4380 19836 4384
rect 19772 4324 19776 4380
rect 19776 4324 19832 4380
rect 19832 4324 19836 4380
rect 19772 4320 19836 4324
rect 19852 4380 19916 4384
rect 19852 4324 19856 4380
rect 19856 4324 19912 4380
rect 19912 4324 19916 4380
rect 19852 4320 19916 4324
rect 8416 3836 8480 3840
rect 8416 3780 8420 3836
rect 8420 3780 8476 3836
rect 8476 3780 8480 3836
rect 8416 3776 8480 3780
rect 8496 3836 8560 3840
rect 8496 3780 8500 3836
rect 8500 3780 8556 3836
rect 8556 3780 8560 3836
rect 8496 3776 8560 3780
rect 8576 3836 8640 3840
rect 8576 3780 8580 3836
rect 8580 3780 8636 3836
rect 8636 3780 8640 3836
rect 8576 3776 8640 3780
rect 8656 3836 8720 3840
rect 8656 3780 8660 3836
rect 8660 3780 8716 3836
rect 8716 3780 8720 3836
rect 8656 3776 8720 3780
rect 15880 3836 15944 3840
rect 15880 3780 15884 3836
rect 15884 3780 15940 3836
rect 15940 3780 15944 3836
rect 15880 3776 15944 3780
rect 15960 3836 16024 3840
rect 15960 3780 15964 3836
rect 15964 3780 16020 3836
rect 16020 3780 16024 3836
rect 15960 3776 16024 3780
rect 16040 3836 16104 3840
rect 16040 3780 16044 3836
rect 16044 3780 16100 3836
rect 16100 3780 16104 3836
rect 16040 3776 16104 3780
rect 16120 3836 16184 3840
rect 16120 3780 16124 3836
rect 16124 3780 16180 3836
rect 16180 3780 16184 3836
rect 16120 3776 16184 3780
rect 4684 3292 4748 3296
rect 4684 3236 4688 3292
rect 4688 3236 4744 3292
rect 4744 3236 4748 3292
rect 4684 3232 4748 3236
rect 4764 3292 4828 3296
rect 4764 3236 4768 3292
rect 4768 3236 4824 3292
rect 4824 3236 4828 3292
rect 4764 3232 4828 3236
rect 4844 3292 4908 3296
rect 4844 3236 4848 3292
rect 4848 3236 4904 3292
rect 4904 3236 4908 3292
rect 4844 3232 4908 3236
rect 4924 3292 4988 3296
rect 4924 3236 4928 3292
rect 4928 3236 4984 3292
rect 4984 3236 4988 3292
rect 4924 3232 4988 3236
rect 12148 3292 12212 3296
rect 12148 3236 12152 3292
rect 12152 3236 12208 3292
rect 12208 3236 12212 3292
rect 12148 3232 12212 3236
rect 12228 3292 12292 3296
rect 12228 3236 12232 3292
rect 12232 3236 12288 3292
rect 12288 3236 12292 3292
rect 12228 3232 12292 3236
rect 12308 3292 12372 3296
rect 12308 3236 12312 3292
rect 12312 3236 12368 3292
rect 12368 3236 12372 3292
rect 12308 3232 12372 3236
rect 12388 3292 12452 3296
rect 12388 3236 12392 3292
rect 12392 3236 12448 3292
rect 12448 3236 12452 3292
rect 12388 3232 12452 3236
rect 19612 3292 19676 3296
rect 19612 3236 19616 3292
rect 19616 3236 19672 3292
rect 19672 3236 19676 3292
rect 19612 3232 19676 3236
rect 19692 3292 19756 3296
rect 19692 3236 19696 3292
rect 19696 3236 19752 3292
rect 19752 3236 19756 3292
rect 19692 3232 19756 3236
rect 19772 3292 19836 3296
rect 19772 3236 19776 3292
rect 19776 3236 19832 3292
rect 19832 3236 19836 3292
rect 19772 3232 19836 3236
rect 19852 3292 19916 3296
rect 19852 3236 19856 3292
rect 19856 3236 19912 3292
rect 19912 3236 19916 3292
rect 19852 3232 19916 3236
rect 8416 2748 8480 2752
rect 8416 2692 8420 2748
rect 8420 2692 8476 2748
rect 8476 2692 8480 2748
rect 8416 2688 8480 2692
rect 8496 2748 8560 2752
rect 8496 2692 8500 2748
rect 8500 2692 8556 2748
rect 8556 2692 8560 2748
rect 8496 2688 8560 2692
rect 8576 2748 8640 2752
rect 8576 2692 8580 2748
rect 8580 2692 8636 2748
rect 8636 2692 8640 2748
rect 8576 2688 8640 2692
rect 8656 2748 8720 2752
rect 8656 2692 8660 2748
rect 8660 2692 8716 2748
rect 8716 2692 8720 2748
rect 8656 2688 8720 2692
rect 15880 2748 15944 2752
rect 15880 2692 15884 2748
rect 15884 2692 15940 2748
rect 15940 2692 15944 2748
rect 15880 2688 15944 2692
rect 15960 2748 16024 2752
rect 15960 2692 15964 2748
rect 15964 2692 16020 2748
rect 16020 2692 16024 2748
rect 15960 2688 16024 2692
rect 16040 2748 16104 2752
rect 16040 2692 16044 2748
rect 16044 2692 16100 2748
rect 16100 2692 16104 2748
rect 16040 2688 16104 2692
rect 16120 2748 16184 2752
rect 16120 2692 16124 2748
rect 16124 2692 16180 2748
rect 16180 2692 16184 2748
rect 16120 2688 16184 2692
rect 4684 2204 4748 2208
rect 4684 2148 4688 2204
rect 4688 2148 4744 2204
rect 4744 2148 4748 2204
rect 4684 2144 4748 2148
rect 4764 2204 4828 2208
rect 4764 2148 4768 2204
rect 4768 2148 4824 2204
rect 4824 2148 4828 2204
rect 4764 2144 4828 2148
rect 4844 2204 4908 2208
rect 4844 2148 4848 2204
rect 4848 2148 4904 2204
rect 4904 2148 4908 2204
rect 4844 2144 4908 2148
rect 4924 2204 4988 2208
rect 4924 2148 4928 2204
rect 4928 2148 4984 2204
rect 4984 2148 4988 2204
rect 4924 2144 4988 2148
rect 12148 2204 12212 2208
rect 12148 2148 12152 2204
rect 12152 2148 12208 2204
rect 12208 2148 12212 2204
rect 12148 2144 12212 2148
rect 12228 2204 12292 2208
rect 12228 2148 12232 2204
rect 12232 2148 12288 2204
rect 12288 2148 12292 2204
rect 12228 2144 12292 2148
rect 12308 2204 12372 2208
rect 12308 2148 12312 2204
rect 12312 2148 12368 2204
rect 12368 2148 12372 2204
rect 12308 2144 12372 2148
rect 12388 2204 12452 2208
rect 12388 2148 12392 2204
rect 12392 2148 12448 2204
rect 12448 2148 12452 2204
rect 12388 2144 12452 2148
rect 19612 2204 19676 2208
rect 19612 2148 19616 2204
rect 19616 2148 19672 2204
rect 19672 2148 19676 2204
rect 19612 2144 19676 2148
rect 19692 2204 19756 2208
rect 19692 2148 19696 2204
rect 19696 2148 19752 2204
rect 19752 2148 19756 2204
rect 19692 2144 19756 2148
rect 19772 2204 19836 2208
rect 19772 2148 19776 2204
rect 19776 2148 19832 2204
rect 19832 2148 19836 2204
rect 19772 2144 19836 2148
rect 19852 2204 19916 2208
rect 19852 2148 19856 2204
rect 19856 2148 19912 2204
rect 19912 2148 19916 2204
rect 19852 2144 19916 2148
<< metal4 >>
rect 4676 21792 4996 22352
rect 4676 21728 4684 21792
rect 4748 21728 4764 21792
rect 4828 21728 4844 21792
rect 4908 21728 4924 21792
rect 4988 21728 4996 21792
rect 4676 20704 4996 21728
rect 4676 20640 4684 20704
rect 4748 20640 4764 20704
rect 4828 20640 4844 20704
rect 4908 20640 4924 20704
rect 4988 20640 4996 20704
rect 4676 19616 4996 20640
rect 4676 19552 4684 19616
rect 4748 19552 4764 19616
rect 4828 19552 4844 19616
rect 4908 19552 4924 19616
rect 4988 19552 4996 19616
rect 4676 18528 4996 19552
rect 4676 18464 4684 18528
rect 4748 18464 4764 18528
rect 4828 18464 4844 18528
rect 4908 18464 4924 18528
rect 4988 18464 4996 18528
rect 4676 17440 4996 18464
rect 4676 17376 4684 17440
rect 4748 17376 4764 17440
rect 4828 17376 4844 17440
rect 4908 17376 4924 17440
rect 4988 17376 4996 17440
rect 4676 16352 4996 17376
rect 4676 16288 4684 16352
rect 4748 16288 4764 16352
rect 4828 16288 4844 16352
rect 4908 16288 4924 16352
rect 4988 16288 4996 16352
rect 4676 15264 4996 16288
rect 4676 15200 4684 15264
rect 4748 15200 4764 15264
rect 4828 15200 4844 15264
rect 4908 15200 4924 15264
rect 4988 15200 4996 15264
rect 4676 14176 4996 15200
rect 4676 14112 4684 14176
rect 4748 14112 4764 14176
rect 4828 14112 4844 14176
rect 4908 14112 4924 14176
rect 4988 14112 4996 14176
rect 4676 13088 4996 14112
rect 4676 13024 4684 13088
rect 4748 13024 4764 13088
rect 4828 13024 4844 13088
rect 4908 13024 4924 13088
rect 4988 13024 4996 13088
rect 4676 12000 4996 13024
rect 4676 11936 4684 12000
rect 4748 11936 4764 12000
rect 4828 11936 4844 12000
rect 4908 11936 4924 12000
rect 4988 11936 4996 12000
rect 4676 10912 4996 11936
rect 4676 10848 4684 10912
rect 4748 10848 4764 10912
rect 4828 10848 4844 10912
rect 4908 10848 4924 10912
rect 4988 10848 4996 10912
rect 4676 9824 4996 10848
rect 4676 9760 4684 9824
rect 4748 9760 4764 9824
rect 4828 9760 4844 9824
rect 4908 9760 4924 9824
rect 4988 9760 4996 9824
rect 4676 8736 4996 9760
rect 4676 8672 4684 8736
rect 4748 8672 4764 8736
rect 4828 8672 4844 8736
rect 4908 8672 4924 8736
rect 4988 8672 4996 8736
rect 4676 7648 4996 8672
rect 4676 7584 4684 7648
rect 4748 7584 4764 7648
rect 4828 7584 4844 7648
rect 4908 7584 4924 7648
rect 4988 7584 4996 7648
rect 4676 6560 4996 7584
rect 4676 6496 4684 6560
rect 4748 6496 4764 6560
rect 4828 6496 4844 6560
rect 4908 6496 4924 6560
rect 4988 6496 4996 6560
rect 4676 5472 4996 6496
rect 4676 5408 4684 5472
rect 4748 5408 4764 5472
rect 4828 5408 4844 5472
rect 4908 5408 4924 5472
rect 4988 5408 4996 5472
rect 4676 4384 4996 5408
rect 4676 4320 4684 4384
rect 4748 4320 4764 4384
rect 4828 4320 4844 4384
rect 4908 4320 4924 4384
rect 4988 4320 4996 4384
rect 4676 3296 4996 4320
rect 4676 3232 4684 3296
rect 4748 3232 4764 3296
rect 4828 3232 4844 3296
rect 4908 3232 4924 3296
rect 4988 3232 4996 3296
rect 4676 2208 4996 3232
rect 4676 2144 4684 2208
rect 4748 2144 4764 2208
rect 4828 2144 4844 2208
rect 4908 2144 4924 2208
rect 4988 2144 4996 2208
rect 4676 2128 4996 2144
rect 8408 22336 8728 22352
rect 8408 22272 8416 22336
rect 8480 22272 8496 22336
rect 8560 22272 8576 22336
rect 8640 22272 8656 22336
rect 8720 22272 8728 22336
rect 8408 21248 8728 22272
rect 8408 21184 8416 21248
rect 8480 21184 8496 21248
rect 8560 21184 8576 21248
rect 8640 21184 8656 21248
rect 8720 21184 8728 21248
rect 8408 20160 8728 21184
rect 8408 20096 8416 20160
rect 8480 20096 8496 20160
rect 8560 20096 8576 20160
rect 8640 20096 8656 20160
rect 8720 20096 8728 20160
rect 8408 19072 8728 20096
rect 8408 19008 8416 19072
rect 8480 19008 8496 19072
rect 8560 19008 8576 19072
rect 8640 19008 8656 19072
rect 8720 19008 8728 19072
rect 8408 17984 8728 19008
rect 8408 17920 8416 17984
rect 8480 17920 8496 17984
rect 8560 17920 8576 17984
rect 8640 17920 8656 17984
rect 8720 17920 8728 17984
rect 8408 16896 8728 17920
rect 8408 16832 8416 16896
rect 8480 16832 8496 16896
rect 8560 16832 8576 16896
rect 8640 16832 8656 16896
rect 8720 16832 8728 16896
rect 8408 15808 8728 16832
rect 8408 15744 8416 15808
rect 8480 15744 8496 15808
rect 8560 15744 8576 15808
rect 8640 15744 8656 15808
rect 8720 15744 8728 15808
rect 8408 14720 8728 15744
rect 8408 14656 8416 14720
rect 8480 14656 8496 14720
rect 8560 14656 8576 14720
rect 8640 14656 8656 14720
rect 8720 14656 8728 14720
rect 8408 13632 8728 14656
rect 8408 13568 8416 13632
rect 8480 13568 8496 13632
rect 8560 13568 8576 13632
rect 8640 13568 8656 13632
rect 8720 13568 8728 13632
rect 8408 12544 8728 13568
rect 8408 12480 8416 12544
rect 8480 12480 8496 12544
rect 8560 12480 8576 12544
rect 8640 12480 8656 12544
rect 8720 12480 8728 12544
rect 8408 11456 8728 12480
rect 8408 11392 8416 11456
rect 8480 11392 8496 11456
rect 8560 11392 8576 11456
rect 8640 11392 8656 11456
rect 8720 11392 8728 11456
rect 8408 10368 8728 11392
rect 8408 10304 8416 10368
rect 8480 10304 8496 10368
rect 8560 10304 8576 10368
rect 8640 10304 8656 10368
rect 8720 10304 8728 10368
rect 8408 9280 8728 10304
rect 8408 9216 8416 9280
rect 8480 9216 8496 9280
rect 8560 9216 8576 9280
rect 8640 9216 8656 9280
rect 8720 9216 8728 9280
rect 8408 8192 8728 9216
rect 8408 8128 8416 8192
rect 8480 8128 8496 8192
rect 8560 8128 8576 8192
rect 8640 8128 8656 8192
rect 8720 8128 8728 8192
rect 8408 7104 8728 8128
rect 8408 7040 8416 7104
rect 8480 7040 8496 7104
rect 8560 7040 8576 7104
rect 8640 7040 8656 7104
rect 8720 7040 8728 7104
rect 8408 6016 8728 7040
rect 8408 5952 8416 6016
rect 8480 5952 8496 6016
rect 8560 5952 8576 6016
rect 8640 5952 8656 6016
rect 8720 5952 8728 6016
rect 8408 4928 8728 5952
rect 8408 4864 8416 4928
rect 8480 4864 8496 4928
rect 8560 4864 8576 4928
rect 8640 4864 8656 4928
rect 8720 4864 8728 4928
rect 8408 3840 8728 4864
rect 8408 3776 8416 3840
rect 8480 3776 8496 3840
rect 8560 3776 8576 3840
rect 8640 3776 8656 3840
rect 8720 3776 8728 3840
rect 8408 2752 8728 3776
rect 8408 2688 8416 2752
rect 8480 2688 8496 2752
rect 8560 2688 8576 2752
rect 8640 2688 8656 2752
rect 8720 2688 8728 2752
rect 8408 2128 8728 2688
rect 12140 21792 12460 22352
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 20704 12460 21728
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 19616 12460 20640
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 18528 12460 19552
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 17440 12460 18464
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 16352 12460 17376
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 15264 12460 16288
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 14176 12460 15200
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 13088 12460 14112
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 12000 12460 13024
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 10912 12460 11936
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 9824 12460 10848
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 8736 12460 9760
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 7648 12460 8672
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 6560 12460 7584
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 5472 12460 6496
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 4384 12460 5408
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 3296 12460 4320
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 2208 12460 3232
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2128 12460 2144
rect 15872 22336 16192 22352
rect 15872 22272 15880 22336
rect 15944 22272 15960 22336
rect 16024 22272 16040 22336
rect 16104 22272 16120 22336
rect 16184 22272 16192 22336
rect 15872 21248 16192 22272
rect 15872 21184 15880 21248
rect 15944 21184 15960 21248
rect 16024 21184 16040 21248
rect 16104 21184 16120 21248
rect 16184 21184 16192 21248
rect 15872 20160 16192 21184
rect 15872 20096 15880 20160
rect 15944 20096 15960 20160
rect 16024 20096 16040 20160
rect 16104 20096 16120 20160
rect 16184 20096 16192 20160
rect 15872 19072 16192 20096
rect 15872 19008 15880 19072
rect 15944 19008 15960 19072
rect 16024 19008 16040 19072
rect 16104 19008 16120 19072
rect 16184 19008 16192 19072
rect 15872 17984 16192 19008
rect 15872 17920 15880 17984
rect 15944 17920 15960 17984
rect 16024 17920 16040 17984
rect 16104 17920 16120 17984
rect 16184 17920 16192 17984
rect 15872 16896 16192 17920
rect 15872 16832 15880 16896
rect 15944 16832 15960 16896
rect 16024 16832 16040 16896
rect 16104 16832 16120 16896
rect 16184 16832 16192 16896
rect 15872 15808 16192 16832
rect 15872 15744 15880 15808
rect 15944 15744 15960 15808
rect 16024 15744 16040 15808
rect 16104 15744 16120 15808
rect 16184 15744 16192 15808
rect 15872 14720 16192 15744
rect 15872 14656 15880 14720
rect 15944 14656 15960 14720
rect 16024 14656 16040 14720
rect 16104 14656 16120 14720
rect 16184 14656 16192 14720
rect 15872 13632 16192 14656
rect 15872 13568 15880 13632
rect 15944 13568 15960 13632
rect 16024 13568 16040 13632
rect 16104 13568 16120 13632
rect 16184 13568 16192 13632
rect 15872 12544 16192 13568
rect 15872 12480 15880 12544
rect 15944 12480 15960 12544
rect 16024 12480 16040 12544
rect 16104 12480 16120 12544
rect 16184 12480 16192 12544
rect 15872 11456 16192 12480
rect 15872 11392 15880 11456
rect 15944 11392 15960 11456
rect 16024 11392 16040 11456
rect 16104 11392 16120 11456
rect 16184 11392 16192 11456
rect 15872 10368 16192 11392
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 9280 16192 10304
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 8192 16192 9216
rect 19604 21792 19924 22352
rect 19604 21728 19612 21792
rect 19676 21728 19692 21792
rect 19756 21728 19772 21792
rect 19836 21728 19852 21792
rect 19916 21728 19924 21792
rect 19604 20704 19924 21728
rect 19604 20640 19612 20704
rect 19676 20640 19692 20704
rect 19756 20640 19772 20704
rect 19836 20640 19852 20704
rect 19916 20640 19924 20704
rect 19604 19616 19924 20640
rect 19604 19552 19612 19616
rect 19676 19552 19692 19616
rect 19756 19552 19772 19616
rect 19836 19552 19852 19616
rect 19916 19552 19924 19616
rect 19604 18528 19924 19552
rect 19604 18464 19612 18528
rect 19676 18464 19692 18528
rect 19756 18464 19772 18528
rect 19836 18464 19852 18528
rect 19916 18464 19924 18528
rect 19604 17440 19924 18464
rect 19604 17376 19612 17440
rect 19676 17376 19692 17440
rect 19756 17376 19772 17440
rect 19836 17376 19852 17440
rect 19916 17376 19924 17440
rect 19604 16352 19924 17376
rect 19604 16288 19612 16352
rect 19676 16288 19692 16352
rect 19756 16288 19772 16352
rect 19836 16288 19852 16352
rect 19916 16288 19924 16352
rect 19604 15264 19924 16288
rect 19604 15200 19612 15264
rect 19676 15200 19692 15264
rect 19756 15200 19772 15264
rect 19836 15200 19852 15264
rect 19916 15200 19924 15264
rect 19604 14176 19924 15200
rect 19604 14112 19612 14176
rect 19676 14112 19692 14176
rect 19756 14112 19772 14176
rect 19836 14112 19852 14176
rect 19916 14112 19924 14176
rect 19604 13088 19924 14112
rect 19604 13024 19612 13088
rect 19676 13024 19692 13088
rect 19756 13024 19772 13088
rect 19836 13024 19852 13088
rect 19916 13024 19924 13088
rect 19604 12000 19924 13024
rect 19604 11936 19612 12000
rect 19676 11936 19692 12000
rect 19756 11936 19772 12000
rect 19836 11936 19852 12000
rect 19916 11936 19924 12000
rect 19604 10912 19924 11936
rect 19604 10848 19612 10912
rect 19676 10848 19692 10912
rect 19756 10848 19772 10912
rect 19836 10848 19852 10912
rect 19916 10848 19924 10912
rect 19604 9824 19924 10848
rect 19604 9760 19612 9824
rect 19676 9760 19692 9824
rect 19756 9760 19772 9824
rect 19836 9760 19852 9824
rect 19916 9760 19924 9824
rect 19379 9212 19445 9213
rect 19379 9148 19380 9212
rect 19444 9148 19445 9212
rect 19379 9147 19445 9148
rect 19382 8397 19442 9147
rect 19604 8736 19924 9760
rect 19604 8672 19612 8736
rect 19676 8672 19692 8736
rect 19756 8672 19772 8736
rect 19836 8672 19852 8736
rect 19916 8672 19924 8736
rect 19379 8396 19445 8397
rect 19379 8332 19380 8396
rect 19444 8332 19445 8396
rect 19379 8331 19445 8332
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 15872 7104 16192 8128
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 6016 16192 7040
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 4928 16192 5952
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 15872 3840 16192 4864
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 2752 16192 3776
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 2128 16192 2688
rect 19604 7648 19924 8672
rect 19604 7584 19612 7648
rect 19676 7584 19692 7648
rect 19756 7584 19772 7648
rect 19836 7584 19852 7648
rect 19916 7584 19924 7648
rect 19604 6560 19924 7584
rect 19604 6496 19612 6560
rect 19676 6496 19692 6560
rect 19756 6496 19772 6560
rect 19836 6496 19852 6560
rect 19916 6496 19924 6560
rect 19604 5472 19924 6496
rect 19604 5408 19612 5472
rect 19676 5408 19692 5472
rect 19756 5408 19772 5472
rect 19836 5408 19852 5472
rect 19916 5408 19924 5472
rect 19604 4384 19924 5408
rect 19604 4320 19612 4384
rect 19676 4320 19692 4384
rect 19756 4320 19772 4384
rect 19836 4320 19852 4384
rect 19916 4320 19924 4384
rect 19604 3296 19924 4320
rect 19604 3232 19612 3296
rect 19676 3232 19692 3296
rect 19756 3232 19772 3296
rect 19836 3232 19852 3296
rect 19916 3232 19924 3296
rect 19604 2208 19924 3232
rect 19604 2144 19612 2208
rect 19676 2144 19692 2208
rect 19756 2144 19772 2208
rect 19836 2144 19852 2208
rect 19916 2144 19924 2208
rect 19604 2128 19924 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1608910539
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_21 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3036 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_33
timestamp 1608910539
transform 1 0 4140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_45 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _64_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_55
timestamp 1608910539
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608910539
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608910539
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608910539
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608910539
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 16468 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1608910539
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608910539
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1608910539
transform 1 0 19228 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_207
timestamp 1608910539
transform 1 0 20148 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1608910539
transform 1 0 19780 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 20792 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 19320 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 20240 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_239
timestamp 1608910539
transform 1 0 23092 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 23460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 23460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608910539
transform 1 0 22632 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 22264 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608910539
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1608910539
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 16468 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 17940 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1608910539
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 20240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 19412 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 23460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 22356 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608910539
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608910539
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608910539
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_159
timestamp 1608910539
transform 1 0 15732 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 16284 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608910539
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 18216 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_3_218
timestamp 1608910539
transform 1 0 21160 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 19688 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_237
timestamp 1608910539
transform 1 0 22908 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1608910539
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 21436 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608910539
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_126
timestamp 1608910539
transform 1 0 12696 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_114
timestamp 1608910539
transform 1 0 11592 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1608910539
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_138
timestamp 1608910539
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16376 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17848 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608910539
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 19504 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608910539
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 21344 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 23000 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 23460 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 21528 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608910539
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608910539
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1608910539
transform 1 0 10856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_98
timestamp 1608910539
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 10948 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1608910539
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_145
timestamp 1608910539
transform 1 0 14444 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_139
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1608910539
transform 1 0 15548 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15916 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1608910539
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 18860 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_211
timestamp 1608910539
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 20700 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A
timestamp 1608910539
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 21528 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_82
timestamp 1608910539
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_74
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1608910539
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1608910539
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 8924 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 9936 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1608910539
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1608910539
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 12696 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 12880 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 11408 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 14168 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 14352 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_163
timestamp 1608910539
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17112 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15640 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16376 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_6_191
timestamp 1608910539
transform 1 0 18676 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18676 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18952 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 18308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19504 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 20976 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 23460 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 23460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 21712 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 22724 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 21804 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1608910539
transform 1 0 22172 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608910539
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608910539
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 13984 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16744 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_191
timestamp 1608910539
transform 1 0 18676 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18952 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608910539
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1608910539
transform 1 0 23092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 23460 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 21896 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 22724 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608910539
transform 1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_86
timestamp 1608910539
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 9292 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1608910539
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 11592 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1608910539
transform 1 0 13616 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 13708 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14168 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15364 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_200
timestamp 1608910539
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 20424 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_239
timestamp 1608910539
transform 1 0 23092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 23460 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 21896 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 22724 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608910539
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608910539
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608910539
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_86
timestamp 1608910539
transform 1 0 9016 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_68
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_FTB00_A
timestamp 1608910539
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  Test_en_FTB00
timestamp 1608910539
transform 1 0 7728 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 11132 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_118
timestamp 1608910539
transform 1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12236 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1608910539
transform 1 0 13892 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 13984 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1608910539
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 16008 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608910539
transform 1 0 15640 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608910539
transform 1 0 17940 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 18492 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1608910539
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 21160 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608910539
transform 1 0 20424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 23460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01
timestamp 1608910539
transform 1 0 22632 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1608910539
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1608910539
transform 1 0 1748 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608910539
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608910539
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1608910539
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1608910539
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13892 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 14720 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17112 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608910539
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1608910539
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18492 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 19964 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 1608910539
transform 1 0 23092 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 23460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 22724 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 21896 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608910539
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608910539
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_109
timestamp 1608910539
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11776 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 11408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13248 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 16744 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17020 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18492 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1608910539
transform 1 0 21068 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19964 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_239
timestamp 1608910539
transform 1 0 23092 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 23460 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 21620 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608910539
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608910539
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608910539
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608910539
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_68
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_86
timestamp 1608910539
transform 1 0 9016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608910539
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1608910539
transform 1 0 9936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1608910539
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_119
timestamp 1608910539
transform 1 0 12052 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_111
timestamp 1608910539
transform 1 0 11316 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_112
timestamp 1608910539
transform 1 0 11408 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 12328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 12880 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1608910539
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14168 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_170
timestamp 1608910539
transform 1 0 16744 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1608910539
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17112 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 17480 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608910539
transform 1 0 17204 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1608910539
transform 1 0 20332 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_199
timestamp 1608910539
transform 1 0 19412 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19504 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 19780 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608910539
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1608910539
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_E_FTB01_A
timestamp 1608910539
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 23460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 22356 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 21252 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 22264 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_17
timestamp 1608910539
transform 1 0 2668 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_5
timestamp 1608910539
transform 1 0 1564 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_41
timestamp 1608910539
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_29
timestamp 1608910539
transform 1 0 3772 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1608910539
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_83
timestamp 1608910539
transform 1 0 8740 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1608910539
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 7268 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 10764 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 9292 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608910539
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 12696 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14996 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 16468 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1608910539
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_198
timestamp 1608910539
transform 1 0 19320 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 19412 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_15_239
timestamp 1608910539
transform 1 0 23092 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 21344 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608910539
transform 1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_19
timestamp 1608910539
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1608910539
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 6808 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 8280 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 9844 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_124
timestamp 1608910539
transform 1 0 12512 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1608910539
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 12880 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14352 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_171
timestamp 1608910539
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17112 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15364 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18768 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1608910539
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608910539
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 23460 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 21712 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1608910539
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1608910539
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_38
timestamp 1608910539
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3128 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1608910539
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_50
timestamp 1608910539
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 6992 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1608910539
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 10396 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608910539
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1608910539
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 12880 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1608910539
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16468 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_176
timestamp 1608910539
transform 1 0 17296 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_204
timestamp 1608910539
transform 1 0 19872 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 20148 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 19504 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 22080 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1608910539
transform 1 0 22908 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1608910539
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608910539
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_26
timestamp 1608910539
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8464 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_96
timestamp 1608910539
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 10120 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11592 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 13432 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.clb_clk
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16376 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15548 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1608910539
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19044 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 18216 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_204
timestamp 1608910539
transform 1 0 19872 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19964 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 21160 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_234
timestamp 1608910539
transform 1 0 22632 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 23460 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1608910539
transform 1 0 4876 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1608910539
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4048 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 4968 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_55
timestamp 1608910539
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6992 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1608910539
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 7268 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_102
timestamp 1608910539
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1608910539
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 10856 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 10580 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1608910539
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 12972 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 13156 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1608910539
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14444 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 16744 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 16100 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 15272 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 18216 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_202
timestamp 1608910539
transform 1 0 19688 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1608910539
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19964 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 20516 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1608910539
transform 1 0 23092 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 23460 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 22356 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1608910539
transform 1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 1472 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 2944 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_42
timestamp 1608910539
transform 1 0 4968 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 4600 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3772 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5060 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5888 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1608910539
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7360 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1608910539
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.clb_clk
timestamp 1608910539
transform 1 0 13800 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 15640 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 17112 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608910539
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 19964 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 19504 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_21_238
timestamp 1608910539
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 23460 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 21896 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1608910539
transform 1 0 22724 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 1748 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1608910539
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_23
timestamp 1608910539
transform 1 0 3220 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_59
timestamp 1608910539
transform 1 0 6532 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 5704 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1608910539
transform 1 0 8740 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 8832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11316 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 12788 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 13340 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1608910539
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 16284 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 18124 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18400 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 17756 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1608910539
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 20332 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 20148 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 19872 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_239
timestamp 1608910539
transform 1 0 23092 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 23460 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 21620 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1608910539
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 2024 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 4968 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 3496 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 8832 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10120 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9292 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_130
timestamp 1608910539
transform 1 0 13064 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1608910539
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.clb_clk
timestamp 1608910539
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13156 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 11776 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1608910539
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 16468 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_190
timestamp 1608910539
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1608910539
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 17664 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 18676 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 17296 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1608910539
transform 1 0 20976 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 20148 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1608910539
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 21344 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 22816 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 1564 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3036 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608910539
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1608910539
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 5520 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 7084 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7544 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1608910539
transform 1 0 9016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10764 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 12236 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608910539
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1608910539
transform 1 0 16744 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1608910539
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 17296 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 18952 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608910539
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 23460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 21344 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 22816 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1608910539
transform 1 0 1932 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 2024 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 3496 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 4324 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5520 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8280 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 9108 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 9476 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1608910539
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13892 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1608910539
transform 1 0 14720 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17112 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 15180 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 21160 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 20332 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 19504 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 23460 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 22816 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1608910539
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 1840 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 1656 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1608910539
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4508 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 3312 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4784 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4784 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 3128 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1608910539
transform 1 0 6808 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6900 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 6256 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8188 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8372 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 7636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10672 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9844 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9752 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608910539
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_125
timestamp 1608910539
transform 1 0 12604 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_110
timestamp 1608910539
transform 1 0 11224 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1608910539
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1608910539
transform 1 0 13892 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1608910539
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1608910539
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1608910539
transform 1 0 13984 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13524 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1608910539
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1608910539
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_174
timestamp 1608910539
transform 1 0 17112 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp 1608910539
transform 1 0 15548 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15640 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1608910539
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 17388 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 17664 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1608910539
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 21160 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 20516 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 19964 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 19504 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1608910539
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 23460 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 23460 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 21528 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 22356 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 21528 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 2116 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608910539
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4784 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_56
timestamp 1608910539
transform 1 0 6256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6992 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8464 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1608910539
transform 1 0 11684 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1608910539
transform 1 0 11316 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12604 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1608910539
transform 1 0 14076 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1608910539
transform 1 0 16744 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17112 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 17940 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1608910539
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 21068 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 19412 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 23460 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 21528 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_39
timestamp 1608910539
transform 1 0 4692 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 3220 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4784 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1608910539
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 8832 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1608910539
transform 1 0 8556 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1608910539
transform 1 0 8280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608910539
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1608910539
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11592 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1608910539
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1608910539
transform 1 0 14904 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13248 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1608910539
transform 1 0 16376 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1608910539
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 18584 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 20056 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1608910539
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 21344 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 22816 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 1656 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4416 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 3128 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1608910539
transform 1 0 6440 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 6072 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5244 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 7360 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1608910539
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 13064 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1608910539
transform 1 0 11592 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_150
timestamp 1608910539
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_167
timestamp 1608910539
transform 1 0 16468 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1608910539
transform 1 0 16100 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 16560 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_30_192
timestamp 1608910539
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 18952 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608910539
transform 1 0 18492 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 22356 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1608910539
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 1840 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 2208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 2576 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_34
timestamp 1608910539
transform 1 0 4232 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4508 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3404 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5336 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 6164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1608910539
transform 1 0 7636 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10028 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1608910539
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_116
timestamp 1608910539
transform 1 0 11776 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1608910539
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1608910539
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp 1608910539
transform 1 0 13892 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1608910539
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16468 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1608910539
transform 1 0 18216 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 21160 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 19688 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1608910539
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 23460 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 22632 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 1564 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3036 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608910539
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4876 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6716 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5704 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1608910539
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 8188 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_32_121
timestamp 1608910539
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_113
timestamp 1608910539
transform 1 0 11500 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1608910539
transform 1 0 12512 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1608910539
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14168 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1608910539
transform 1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_195
timestamp 1608910539
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17572 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608910539
transform 1 0 17296 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_215
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1608910539
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 20976 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1608910539
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1608910539
transform 1 0 21804 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 23460 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 21896 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 22632 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 22264 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1608910539
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1608910539
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 1932 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 1564 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 3036 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608910539
transform 1 0 1564 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1608910539
transform 1 0 5060 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1608910539
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1608910539
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 4048 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 3864 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608910539
transform 1 0 4692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608910539
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1608910539
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1608910539
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7084 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6164 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 5520 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 1608910539
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7636 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1608910539
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 11132 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9292 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1608910539
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_114
timestamp 1608910539
transform 1 0 11592 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1608910539
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1608910539
transform 1 0 13156 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1608910539
transform 1 0 11684 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1608910539
transform 1 0 12420 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_147
timestamp 1608910539
transform 1 0 14628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1608910539
transform 1 0 14260 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1608910539
transform 1 0 14352 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1608910539
transform 1 0 14720 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1608910539
transform 1 0 13892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1608910539
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16744 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1608910539
transform 1 0 15824 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1608910539
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1608910539
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18216 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1608910539
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1608910539
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_209
timestamp 1608910539
transform 1 0 20332 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1608910539
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 19504 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_33_221
timestamp 1608910539
transform 1 0 21436 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_227
timestamp 1608910539
transform 1 0 21988 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_227
timestamp 1608910539
transform 1 0 21988 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1608910539
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1608910539
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 22264 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 22264 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_238
timestamp 1608910539
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 23000 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 22632 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1608910539
transform -1 0 23460 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1608910539
transform 1 0 1748 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1608910539
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1608910539
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 2576 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608910539
transform 1 0 2208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608910539
transform 1 0 1840 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_36
timestamp 1608910539
transform 1 0 4416 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4508 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608910539
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1608910539
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 6992 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 6348 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608910539
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1608910539
transform 1 0 8648 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1608910539
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7544 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9016 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1608910539
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10488 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1608910539
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1608910539
transform 1 0 12420 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1608910539
transform 1 0 11960 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1608910539
transform 1 0 13892 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_168
timestamp 1608910539
transform 1 0 16560 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 16192 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1608910539
transform 1 0 15364 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1608910539
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1608910539
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  clk_0_FTB00
timestamp 1608910539
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 17480 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608910539
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_213
timestamp 1608910539
transform 1 0 20700 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_201
timestamp 1608910539
transform 1 0 19596 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1608910539
transform 1 0 21804 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1608910539
transform 1 0 22080 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1608910539
transform -1 0 23460 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 22632 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 22264 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_18
timestamp 1608910539
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_14
timestamp 1608910539
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_11
timestamp 1608910539
transform 1 0 2116 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1608910539
transform 1 0 1380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1608910539
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1608910539
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1608910539
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_43
timestamp 1608910539
transform 1 0 5060 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_38
timestamp 1608910539
transform 1 0 4600 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1608910539
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1608910539
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1608910539
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1608910539
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1608910539
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608910539
transform 1 0 4692 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_65
timestamp 1608910539
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1608910539
transform 1 0 6716 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 6900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1608910539
transform 1 0 6808 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5888 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 5152 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 5520 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_78
timestamp 1608910539
transform 1 0 8280 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 8096 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_36_106
timestamp 1608910539
transform 1 0 10856 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_90
timestamp 1608910539
transform 1 0 9384 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1608910539
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9752 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1608910539
transform 1 0 10580 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_125
timestamp 1608910539
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1608910539
transform 1 0 11960 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1608910539
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1608910539
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1608910539
transform 1 0 12880 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1608910539
transform 1 0 13708 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1608910539
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1608910539
transform 1 0 13984 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_36_174
timestamp 1608910539
transform 1 0 17112 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_166
timestamp 1608910539
transform 1 0 16376 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1608910539
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1608910539
transform 1 0 15180 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1608910539
transform 1 0 15364 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1608910539
transform 1 0 15824 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1608910539
transform 1 0 15456 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_189
timestamp 1608910539
transform 1 0 18492 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1608910539
transform 1 0 18308 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1608910539
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 17388 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_36_218
timestamp 1608910539
transform 1 0 21160 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1608910539
transform 1 0 20700 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1608910539
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1608910539
transform 1 0 21068 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_238
timestamp 1608910539
transform 1 0 23000 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_230
timestamp 1608910539
transform 1 0 22264 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1608910539
transform -1 0 23460 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal2 s 17038 23800 17094 24600 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 17682 23800 17738 24600 6 SC_OUT_TOP
port 2 nsew signal tristate
rlabel metal3 s 23800 6808 24600 6928 6 Test_en_E_in
port 3 nsew signal input
rlabel metal3 s 23800 6264 24600 6384 6 Test_en_E_out
port 4 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 Test_en_W_in
port 5 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 Test_en_W_out
port 6 nsew signal tristate
rlabel metal2 s 2042 0 2098 800 6 bottom_width_0_height_0__pin_50_
port 7 nsew signal tristate
rlabel metal2 s 6090 0 6146 800 6 bottom_width_0_height_0__pin_51_
port 8 nsew signal tristate
rlabel metal3 s 0 9120 800 9240 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 23800 5584 24600 5704 6 ccff_tail
port 10 nsew signal tristate
rlabel metal2 s 18326 23800 18382 24600 6 clk_0_N_in
port 11 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 clk_0_S_in
port 12 nsew signal input
rlabel metal3 s 23800 8168 24600 8288 6 prog_clk_0_E_out
port 13 nsew signal tristate
rlabel metal3 s 23800 7488 24600 7608 6 prog_clk_0_N_in
port 14 nsew signal input
rlabel metal2 s 18970 23800 19026 24600 6 prog_clk_0_N_out
port 15 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 prog_clk_0_S_in
port 16 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 prog_clk_0_S_out
port 17 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 prog_clk_0_W_out
port 18 nsew signal tristate
rlabel metal3 s 23800 8848 24600 8968 6 right_width_0_height_0__pin_16_
port 19 nsew signal input
rlabel metal3 s 23800 9528 24600 9648 6 right_width_0_height_0__pin_17_
port 20 nsew signal input
rlabel metal3 s 23800 10208 24600 10328 6 right_width_0_height_0__pin_18_
port 21 nsew signal input
rlabel metal3 s 23800 10888 24600 11008 6 right_width_0_height_0__pin_19_
port 22 nsew signal input
rlabel metal3 s 23800 11568 24600 11688 6 right_width_0_height_0__pin_20_
port 23 nsew signal input
rlabel metal3 s 23800 12248 24600 12368 6 right_width_0_height_0__pin_21_
port 24 nsew signal input
rlabel metal3 s 23800 12792 24600 12912 6 right_width_0_height_0__pin_22_
port 25 nsew signal input
rlabel metal3 s 23800 13472 24600 13592 6 right_width_0_height_0__pin_23_
port 26 nsew signal input
rlabel metal3 s 23800 14152 24600 14272 6 right_width_0_height_0__pin_24_
port 27 nsew signal input
rlabel metal3 s 23800 14832 24600 14952 6 right_width_0_height_0__pin_25_
port 28 nsew signal input
rlabel metal3 s 23800 15512 24600 15632 6 right_width_0_height_0__pin_26_
port 29 nsew signal input
rlabel metal3 s 23800 16192 24600 16312 6 right_width_0_height_0__pin_27_
port 30 nsew signal input
rlabel metal3 s 23800 16872 24600 16992 6 right_width_0_height_0__pin_28_
port 31 nsew signal input
rlabel metal3 s 23800 17552 24600 17672 6 right_width_0_height_0__pin_29_
port 32 nsew signal input
rlabel metal3 s 23800 18232 24600 18352 6 right_width_0_height_0__pin_30_
port 33 nsew signal input
rlabel metal3 s 23800 18776 24600 18896 6 right_width_0_height_0__pin_31_
port 34 nsew signal input
rlabel metal3 s 23800 280 24600 400 6 right_width_0_height_0__pin_42_lower
port 35 nsew signal tristate
rlabel metal3 s 23800 19456 24600 19576 6 right_width_0_height_0__pin_42_upper
port 36 nsew signal tristate
rlabel metal3 s 23800 824 24600 944 6 right_width_0_height_0__pin_43_lower
port 37 nsew signal tristate
rlabel metal3 s 23800 20136 24600 20256 6 right_width_0_height_0__pin_43_upper
port 38 nsew signal tristate
rlabel metal3 s 23800 1504 24600 1624 6 right_width_0_height_0__pin_44_lower
port 39 nsew signal tristate
rlabel metal3 s 23800 20816 24600 20936 6 right_width_0_height_0__pin_44_upper
port 40 nsew signal tristate
rlabel metal3 s 23800 2184 24600 2304 6 right_width_0_height_0__pin_45_lower
port 41 nsew signal tristate
rlabel metal3 s 23800 21496 24600 21616 6 right_width_0_height_0__pin_45_upper
port 42 nsew signal tristate
rlabel metal3 s 23800 2864 24600 2984 6 right_width_0_height_0__pin_46_lower
port 43 nsew signal tristate
rlabel metal3 s 23800 22176 24600 22296 6 right_width_0_height_0__pin_46_upper
port 44 nsew signal tristate
rlabel metal3 s 23800 3544 24600 3664 6 right_width_0_height_0__pin_47_lower
port 45 nsew signal tristate
rlabel metal3 s 23800 22856 24600 22976 6 right_width_0_height_0__pin_47_upper
port 46 nsew signal tristate
rlabel metal3 s 23800 4224 24600 4344 6 right_width_0_height_0__pin_48_lower
port 47 nsew signal tristate
rlabel metal3 s 23800 23536 24600 23656 6 right_width_0_height_0__pin_48_upper
port 48 nsew signal tristate
rlabel metal3 s 23800 4904 24600 5024 6 right_width_0_height_0__pin_49_lower
port 49 nsew signal tristate
rlabel metal3 s 23800 24216 24600 24336 6 right_width_0_height_0__pin_49_upper
port 50 nsew signal tristate
rlabel metal2 s 5446 23800 5502 24600 6 top_width_0_height_0__pin_0_
port 51 nsew signal input
rlabel metal2 s 11886 23800 11942 24600 6 top_width_0_height_0__pin_10_
port 52 nsew signal input
rlabel metal2 s 12530 23800 12586 24600 6 top_width_0_height_0__pin_11_
port 53 nsew signal input
rlabel metal2 s 13174 23800 13230 24600 6 top_width_0_height_0__pin_12_
port 54 nsew signal input
rlabel metal2 s 13818 23800 13874 24600 6 top_width_0_height_0__pin_13_
port 55 nsew signal input
rlabel metal2 s 14462 23800 14518 24600 6 top_width_0_height_0__pin_14_
port 56 nsew signal input
rlabel metal2 s 15106 23800 15162 24600 6 top_width_0_height_0__pin_15_
port 57 nsew signal input
rlabel metal2 s 6090 23800 6146 24600 6 top_width_0_height_0__pin_1_
port 58 nsew signal input
rlabel metal2 s 6734 23800 6790 24600 6 top_width_0_height_0__pin_2_
port 59 nsew signal input
rlabel metal2 s 15750 23800 15806 24600 6 top_width_0_height_0__pin_32_
port 60 nsew signal input
rlabel metal2 s 16394 23800 16450 24600 6 top_width_0_height_0__pin_33_
port 61 nsew signal input
rlabel metal2 s 19614 23800 19670 24600 6 top_width_0_height_0__pin_34_lower
port 62 nsew signal tristate
rlabel metal2 s 294 23800 350 24600 6 top_width_0_height_0__pin_34_upper
port 63 nsew signal tristate
rlabel metal2 s 20258 23800 20314 24600 6 top_width_0_height_0__pin_35_lower
port 64 nsew signal tristate
rlabel metal2 s 938 23800 994 24600 6 top_width_0_height_0__pin_35_upper
port 65 nsew signal tristate
rlabel metal2 s 20902 23800 20958 24600 6 top_width_0_height_0__pin_36_lower
port 66 nsew signal tristate
rlabel metal2 s 1582 23800 1638 24600 6 top_width_0_height_0__pin_36_upper
port 67 nsew signal tristate
rlabel metal2 s 21546 23800 21602 24600 6 top_width_0_height_0__pin_37_lower
port 68 nsew signal tristate
rlabel metal2 s 2226 23800 2282 24600 6 top_width_0_height_0__pin_37_upper
port 69 nsew signal tristate
rlabel metal2 s 22190 23800 22246 24600 6 top_width_0_height_0__pin_38_lower
port 70 nsew signal tristate
rlabel metal2 s 2870 23800 2926 24600 6 top_width_0_height_0__pin_38_upper
port 71 nsew signal tristate
rlabel metal2 s 22834 23800 22890 24600 6 top_width_0_height_0__pin_39_lower
port 72 nsew signal tristate
rlabel metal2 s 3514 23800 3570 24600 6 top_width_0_height_0__pin_39_upper
port 73 nsew signal tristate
rlabel metal2 s 7378 23800 7434 24600 6 top_width_0_height_0__pin_3_
port 74 nsew signal input
rlabel metal2 s 23478 23800 23534 24600 6 top_width_0_height_0__pin_40_lower
port 75 nsew signal tristate
rlabel metal2 s 4158 23800 4214 24600 6 top_width_0_height_0__pin_40_upper
port 76 nsew signal tristate
rlabel metal2 s 24122 23800 24178 24600 6 top_width_0_height_0__pin_41_lower
port 77 nsew signal tristate
rlabel metal2 s 4802 23800 4858 24600 6 top_width_0_height_0__pin_41_upper
port 78 nsew signal tristate
rlabel metal2 s 8022 23800 8078 24600 6 top_width_0_height_0__pin_4_
port 79 nsew signal input
rlabel metal2 s 8666 23800 8722 24600 6 top_width_0_height_0__pin_5_
port 80 nsew signal input
rlabel metal2 s 9310 23800 9366 24600 6 top_width_0_height_0__pin_6_
port 81 nsew signal input
rlabel metal2 s 9954 23800 10010 24600 6 top_width_0_height_0__pin_7_
port 82 nsew signal input
rlabel metal2 s 10598 23800 10654 24600 6 top_width_0_height_0__pin_8_
port 83 nsew signal input
rlabel metal2 s 11242 23800 11298 24600 6 top_width_0_height_0__pin_9_
port 84 nsew signal input
rlabel metal4 s 19604 2128 19924 22352 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 12140 2128 12460 22352 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 4676 2128 4996 22352 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 15872 2128 16192 22352 6 VGND
port 88 nsew ground bidirectional
rlabel metal4 s 8408 2128 8728 22352 6 VGND
port 89 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24600 24600
<< end >>
