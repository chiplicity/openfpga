magic
tech sky130A
magscale 1 2
timestamp 1605121657
<< viali >>
rect 23029 25169 23063 25203
rect 24777 25169 24811 25203
rect 22845 25033 22879 25067
rect 24593 25033 24627 25067
rect 11437 24829 11471 24863
rect 11989 24489 12023 24523
rect 23489 24489 23523 24523
rect 11897 24421 11931 24455
rect 22569 24421 22603 24455
rect 23121 24421 23155 24455
rect 23673 24421 23707 24455
rect 24961 24421 24995 24455
rect 25513 24421 25547 24455
rect 23949 24353 23983 24387
rect 11253 24285 11287 24319
rect 11437 24285 11471 24319
rect 11805 24285 11839 24319
rect 16497 24285 16531 24319
rect 17417 24285 17451 24319
rect 22753 24285 22787 24319
rect 24409 24285 24443 24319
rect 24777 24285 24811 24319
rect 25145 24285 25179 24319
rect 21557 24081 21591 24115
rect 23949 24013 23983 24047
rect 14177 23945 14211 23979
rect 16681 23945 16715 23979
rect 19257 23945 19291 23979
rect 21373 23945 21407 23979
rect 21925 23945 21959 23979
rect 22477 23945 22511 23979
rect 23029 23945 23063 23979
rect 23673 23945 23707 23979
rect 24961 23945 24995 23979
rect 13921 23877 13955 23911
rect 16773 23877 16807 23911
rect 16865 23877 16899 23911
rect 19349 23877 19383 23911
rect 19533 23877 19567 23911
rect 16221 23809 16255 23843
rect 20913 23809 20947 23843
rect 22661 23809 22695 23843
rect 25145 23809 25179 23843
rect 11437 23741 11471 23775
rect 13737 23741 13771 23775
rect 15301 23741 15335 23775
rect 16313 23741 16347 23775
rect 18337 23741 18371 23775
rect 18705 23741 18739 23775
rect 18889 23741 18923 23775
rect 20545 23741 20579 23775
rect 24409 23741 24443 23775
rect 13185 23537 13219 23571
rect 13461 23537 13495 23571
rect 16221 23537 16255 23571
rect 18153 23537 18187 23571
rect 18429 23537 18463 23571
rect 19993 23537 20027 23571
rect 20913 23537 20947 23571
rect 23673 23537 23707 23571
rect 24961 23537 24995 23571
rect 22109 23469 22143 23503
rect 14105 23401 14139 23435
rect 14289 23401 14323 23435
rect 21373 23401 21407 23435
rect 21465 23401 21499 23435
rect 23121 23401 23155 23435
rect 24409 23401 24443 23435
rect 11345 23333 11379 23367
rect 11437 23333 11471 23367
rect 16405 23333 16439 23367
rect 18613 23333 18647 23367
rect 20269 23333 20303 23367
rect 22937 23333 22971 23367
rect 24133 23333 24167 23367
rect 10977 23265 11011 23299
rect 11682 23265 11716 23299
rect 14749 23265 14783 23299
rect 15945 23265 15979 23299
rect 16672 23265 16706 23299
rect 18858 23265 18892 23299
rect 22385 23265 22419 23299
rect 23029 23265 23063 23299
rect 12817 23197 12851 23231
rect 13645 23197 13679 23231
rect 14013 23197 14047 23231
rect 15301 23197 15335 23231
rect 17785 23197 17819 23231
rect 20729 23197 20763 23231
rect 21281 23197 21315 23231
rect 22569 23197 22603 23231
rect 9781 22993 9815 23027
rect 11253 22993 11287 23027
rect 15301 22993 15335 23027
rect 16773 22993 16807 23027
rect 19441 22993 19475 23027
rect 24133 22993 24167 23027
rect 25421 22993 25455 23027
rect 14188 22925 14222 22959
rect 15669 22925 15703 22959
rect 16865 22925 16899 22959
rect 19717 22925 19751 22959
rect 20913 22925 20947 22959
rect 24041 22925 24075 22959
rect 11161 22857 11195 22891
rect 12449 22857 12483 22891
rect 18317 22857 18351 22891
rect 21353 22857 21387 22891
rect 25237 22857 25271 22891
rect 11437 22789 11471 22823
rect 12725 22789 12759 22823
rect 13921 22789 13955 22823
rect 17049 22789 17083 22823
rect 18061 22789 18095 22823
rect 21097 22789 21131 22823
rect 24225 22789 24259 22823
rect 10793 22721 10827 22755
rect 16405 22721 16439 22755
rect 13737 22653 13771 22687
rect 16037 22653 16071 22687
rect 20545 22653 20579 22687
rect 22477 22653 22511 22687
rect 22845 22653 22879 22687
rect 23673 22653 23707 22687
rect 10885 22449 10919 22483
rect 12725 22449 12759 22483
rect 13001 22449 13035 22483
rect 14289 22449 14323 22483
rect 17325 22449 17359 22483
rect 17601 22449 17635 22483
rect 18153 22449 18187 22483
rect 18429 22449 18463 22483
rect 20361 22449 20395 22483
rect 22017 22449 22051 22483
rect 22477 22449 22511 22483
rect 23949 22449 23983 22483
rect 24593 22449 24627 22483
rect 11253 22313 11287 22347
rect 11345 22313 11379 22347
rect 14013 22313 14047 22347
rect 15853 22313 15887 22347
rect 15945 22313 15979 22347
rect 19533 22313 19567 22347
rect 21465 22313 21499 22347
rect 22569 22313 22603 22347
rect 11612 22245 11646 22279
rect 16201 22245 16235 22279
rect 24777 22245 24811 22279
rect 25329 22245 25363 22279
rect 10517 22177 10551 22211
rect 20729 22177 20763 22211
rect 21373 22177 21407 22211
rect 22836 22177 22870 22211
rect 20913 22109 20947 22143
rect 21281 22109 21315 22143
rect 24225 22109 24259 22143
rect 24961 22109 24995 22143
rect 25697 22109 25731 22143
rect 11437 21905 11471 21939
rect 14657 21905 14691 21939
rect 17233 21905 17267 21939
rect 22569 21905 22603 21939
rect 20514 21837 20548 21871
rect 23949 21837 23983 21871
rect 10885 21769 10919 21803
rect 14749 21769 14783 21803
rect 16589 21769 16623 21803
rect 18061 21769 18095 21803
rect 18337 21769 18371 21803
rect 24593 21769 24627 21803
rect 14841 21701 14875 21735
rect 16681 21701 16715 21735
rect 16865 21701 16899 21735
rect 20269 21701 20303 21735
rect 14289 21633 14323 21667
rect 16221 21633 16255 21667
rect 18797 21633 18831 21667
rect 11805 21565 11839 21599
rect 15761 21565 15795 21599
rect 16129 21565 16163 21599
rect 21649 21565 21683 21599
rect 23121 21565 23155 21599
rect 24777 21565 24811 21599
rect 11529 21361 11563 21395
rect 14381 21361 14415 21395
rect 14749 21361 14783 21395
rect 15577 21361 15611 21395
rect 16037 21361 16071 21395
rect 19993 21361 20027 21395
rect 22937 21361 22971 21395
rect 24593 21361 24627 21395
rect 15117 21293 15151 21327
rect 22293 21293 22327 21327
rect 12173 21225 12207 21259
rect 12357 21225 12391 21259
rect 16589 21225 16623 21259
rect 18705 21225 18739 21259
rect 21465 21225 21499 21259
rect 21925 21225 21959 21259
rect 23397 21225 23431 21259
rect 24041 21225 24075 21259
rect 13277 21157 13311 21191
rect 21373 21157 21407 21191
rect 22753 21157 22787 21191
rect 23857 21157 23891 21191
rect 25145 21157 25179 21191
rect 25697 21157 25731 21191
rect 13553 21089 13587 21123
rect 16497 21089 16531 21123
rect 18521 21089 18555 21123
rect 20729 21089 20763 21123
rect 21281 21089 21315 21123
rect 11713 21021 11747 21055
rect 12081 21021 12115 21055
rect 13093 21021 13127 21055
rect 15853 21021 15887 21055
rect 16405 21021 16439 21055
rect 17049 21021 17083 21055
rect 17601 21021 17635 21055
rect 18061 21021 18095 21055
rect 18153 21021 18187 21055
rect 18613 21021 18647 21055
rect 19165 21021 19199 21055
rect 20269 21021 20303 21055
rect 20913 21021 20947 21055
rect 23673 21021 23707 21055
rect 25329 21021 25363 21055
rect 14289 20817 14323 20851
rect 14657 20817 14691 20851
rect 17049 20817 17083 20851
rect 18061 20817 18095 20851
rect 12694 20749 12728 20783
rect 18429 20749 18463 20783
rect 20444 20749 20478 20783
rect 15925 20681 15959 20715
rect 23857 20681 23891 20715
rect 25145 20681 25179 20715
rect 12449 20613 12483 20647
rect 15669 20613 15703 20647
rect 18521 20613 18555 20647
rect 18705 20613 18739 20647
rect 20177 20613 20211 20647
rect 24133 20613 24167 20647
rect 25421 20613 25455 20647
rect 11805 20477 11839 20511
rect 13829 20477 13863 20511
rect 15393 20477 15427 20511
rect 21557 20477 21591 20511
rect 22845 20477 22879 20511
rect 12541 20273 12575 20307
rect 14749 20273 14783 20307
rect 16681 20273 16715 20307
rect 17969 20273 18003 20307
rect 19441 20273 19475 20307
rect 20545 20273 20579 20307
rect 24409 20273 24443 20307
rect 25145 20273 25179 20307
rect 25513 20273 25547 20307
rect 19809 20205 19843 20239
rect 24133 20205 24167 20239
rect 17233 20137 17267 20171
rect 20913 20137 20947 20171
rect 10425 20069 10459 20103
rect 10517 20069 10551 20103
rect 12173 20069 12207 20103
rect 12725 20069 12759 20103
rect 12992 20069 13026 20103
rect 15301 20069 15335 20103
rect 15557 20069 15591 20103
rect 18061 20069 18095 20103
rect 18328 20069 18362 20103
rect 22109 20069 22143 20103
rect 22753 20069 22787 20103
rect 23009 20069 23043 20103
rect 24961 20069 24995 20103
rect 10784 20001 10818 20035
rect 20177 20001 20211 20035
rect 11897 19933 11931 19967
rect 14105 19933 14139 19967
rect 15025 19933 15059 19967
rect 17509 19933 17543 19967
rect 22661 19933 22695 19967
rect 24869 19933 24903 19967
rect 10609 19729 10643 19763
rect 12081 19729 12115 19763
rect 13001 19729 13035 19763
rect 13277 19729 13311 19763
rect 15301 19729 15335 19763
rect 18337 19729 18371 19763
rect 22017 19729 22051 19763
rect 24133 19729 24167 19763
rect 25421 19729 25455 19763
rect 13737 19661 13771 19695
rect 14166 19661 14200 19695
rect 13921 19593 13955 19627
rect 15761 19593 15795 19627
rect 18705 19593 18739 19627
rect 18981 19593 19015 19627
rect 22385 19593 22419 19627
rect 24041 19593 24075 19627
rect 25237 19593 25271 19627
rect 12449 19525 12483 19559
rect 16129 19525 16163 19559
rect 22477 19525 22511 19559
rect 22569 19525 22603 19559
rect 24225 19525 24259 19559
rect 21005 19389 21039 19423
rect 21833 19389 21867 19423
rect 23673 19389 23707 19423
rect 14749 19185 14783 19219
rect 18705 19185 18739 19219
rect 24409 19185 24443 19219
rect 24777 19185 24811 19219
rect 25881 19185 25915 19219
rect 20913 19117 20947 19151
rect 22109 19117 22143 19151
rect 24133 19117 24167 19151
rect 12541 19049 12575 19083
rect 12725 19049 12759 19083
rect 14197 19049 14231 19083
rect 15853 19049 15887 19083
rect 21465 19049 21499 19083
rect 22753 19049 22787 19083
rect 11989 18981 12023 19015
rect 12449 18981 12483 19015
rect 15117 18981 15151 19015
rect 15669 18981 15703 19015
rect 18245 18981 18279 19015
rect 24961 18981 24995 19015
rect 25513 18981 25547 19015
rect 13461 18913 13495 18947
rect 14105 18913 14139 18947
rect 21373 18913 21407 18947
rect 22998 18913 23032 18947
rect 12081 18845 12115 18879
rect 13645 18845 13679 18879
rect 14013 18845 14047 18879
rect 15301 18845 15335 18879
rect 15761 18845 15795 18879
rect 20729 18845 20763 18879
rect 21281 18845 21315 18879
rect 22569 18845 22603 18879
rect 25145 18845 25179 18879
rect 12173 18641 12207 18675
rect 13737 18641 13771 18675
rect 14105 18641 14139 18675
rect 15393 18641 15427 18675
rect 15761 18641 15795 18675
rect 20269 18641 20303 18675
rect 22753 18641 22787 18675
rect 23029 18641 23063 18675
rect 25329 18641 25363 18675
rect 16773 18573 16807 18607
rect 23949 18573 23983 18607
rect 18317 18505 18351 18539
rect 21640 18505 21674 18539
rect 24041 18505 24075 18539
rect 16865 18437 16899 18471
rect 17049 18437 17083 18471
rect 18061 18437 18095 18471
rect 20361 18437 20395 18471
rect 21373 18437 21407 18471
rect 24317 18437 24351 18471
rect 16129 18301 16163 18335
rect 16405 18301 16439 18335
rect 19441 18301 19475 18335
rect 21005 18301 21039 18335
rect 15393 18097 15427 18131
rect 16865 18097 16899 18131
rect 17233 18097 17267 18131
rect 17601 18097 17635 18131
rect 22293 18097 22327 18131
rect 22569 18097 22603 18131
rect 24593 18097 24627 18131
rect 25329 18097 25363 18131
rect 15117 17961 15151 17995
rect 15945 17961 15979 17995
rect 16405 17893 16439 17927
rect 18429 17893 18463 17927
rect 20913 17893 20947 17927
rect 21169 17893 21203 17927
rect 23857 17893 23891 17927
rect 25145 17893 25179 17927
rect 25697 17893 25731 17927
rect 15761 17825 15795 17859
rect 18674 17825 18708 17859
rect 20085 17825 20119 17859
rect 24133 17825 24167 17859
rect 14749 17757 14783 17791
rect 15853 17757 15887 17791
rect 17969 17757 18003 17791
rect 18245 17757 18279 17791
rect 19809 17757 19843 17791
rect 20729 17757 20763 17791
rect 23673 17757 23707 17791
rect 14565 17553 14599 17587
rect 17141 17553 17175 17587
rect 18521 17553 18555 17587
rect 21005 17553 21039 17587
rect 21833 17553 21867 17587
rect 22293 17553 22327 17587
rect 24777 17553 24811 17587
rect 16006 17485 16040 17519
rect 21373 17485 21407 17519
rect 14657 17417 14691 17451
rect 15761 17417 15795 17451
rect 18429 17417 18463 17451
rect 19625 17417 19659 17451
rect 19892 17417 19926 17451
rect 22201 17417 22235 17451
rect 24593 17417 24627 17451
rect 14749 17349 14783 17383
rect 18613 17349 18647 17383
rect 19441 17349 19475 17383
rect 22385 17349 22419 17383
rect 14197 17213 14231 17247
rect 15393 17213 15427 17247
rect 18061 17213 18095 17247
rect 19073 17213 19107 17247
rect 15025 17009 15059 17043
rect 16681 17009 16715 17043
rect 17509 17009 17543 17043
rect 19625 17009 19659 17043
rect 21373 17009 21407 17043
rect 25053 17009 25087 17043
rect 25421 17009 25455 17043
rect 18061 16941 18095 16975
rect 23305 16941 23339 16975
rect 15301 16873 15335 16907
rect 18429 16873 18463 16907
rect 19165 16873 19199 16907
rect 22477 16873 22511 16907
rect 14197 16805 14231 16839
rect 15557 16805 15591 16839
rect 17601 16805 17635 16839
rect 18981 16805 19015 16839
rect 23949 16805 23983 16839
rect 24225 16805 24259 16839
rect 25237 16805 25271 16839
rect 25789 16805 25823 16839
rect 13921 16737 13955 16771
rect 19993 16737 20027 16771
rect 21833 16737 21867 16771
rect 22293 16737 22327 16771
rect 24685 16737 24719 16771
rect 14657 16669 14691 16703
rect 18613 16669 18647 16703
rect 19073 16669 19107 16703
rect 21925 16669 21959 16703
rect 22385 16669 22419 16703
rect 22937 16669 22971 16703
rect 15669 16465 15703 16499
rect 16313 16465 16347 16499
rect 18337 16465 18371 16499
rect 18705 16465 18739 16499
rect 19165 16465 19199 16499
rect 20729 16465 20763 16499
rect 25421 16465 25455 16499
rect 14556 16397 14590 16431
rect 16957 16397 16991 16431
rect 21189 16397 21223 16431
rect 21925 16397 21959 16431
rect 15945 16329 15979 16363
rect 19073 16329 19107 16363
rect 21097 16329 21131 16363
rect 22569 16329 22603 16363
rect 23949 16329 23983 16363
rect 24225 16329 24259 16363
rect 25237 16329 25271 16363
rect 14289 16261 14323 16295
rect 16497 16261 16531 16295
rect 19257 16261 19291 16295
rect 21281 16261 21315 16295
rect 22293 16261 22327 16295
rect 14013 15921 14047 15955
rect 15301 15921 15335 15955
rect 16405 15921 16439 15955
rect 19993 15921 20027 15955
rect 21189 15921 21223 15955
rect 23949 15921 23983 15955
rect 24777 15921 24811 15955
rect 25513 15921 25547 15955
rect 16865 15853 16899 15887
rect 15761 15785 15795 15819
rect 15853 15785 15887 15819
rect 17417 15785 17451 15819
rect 18521 15785 18555 15819
rect 19165 15785 19199 15819
rect 22017 15785 22051 15819
rect 17233 15717 17267 15751
rect 17325 15717 17359 15751
rect 22201 15717 22235 15751
rect 22457 15717 22491 15751
rect 24593 15717 24627 15751
rect 25145 15717 25179 15751
rect 16773 15649 16807 15683
rect 18153 15649 18187 15683
rect 19073 15649 19107 15683
rect 20729 15649 20763 15683
rect 14289 15581 14323 15615
rect 14749 15581 14783 15615
rect 15117 15581 15151 15615
rect 15669 15581 15703 15615
rect 18613 15581 18647 15615
rect 18981 15581 19015 15615
rect 19625 15581 19659 15615
rect 21557 15581 21591 15615
rect 23581 15581 23615 15615
rect 15025 15377 15059 15411
rect 15393 15377 15427 15411
rect 16405 15377 16439 15411
rect 18429 15377 18463 15411
rect 18797 15377 18831 15411
rect 20361 15377 20395 15411
rect 22569 15377 22603 15411
rect 22845 15377 22879 15411
rect 24133 15377 24167 15411
rect 25421 15377 25455 15411
rect 19248 15309 19282 15343
rect 13912 15241 13946 15275
rect 16313 15241 16347 15275
rect 21189 15241 21223 15275
rect 21456 15241 21490 15275
rect 24041 15241 24075 15275
rect 25237 15241 25271 15275
rect 13645 15173 13679 15207
rect 16497 15173 16531 15207
rect 18981 15173 19015 15207
rect 24225 15173 24259 15207
rect 15853 15105 15887 15139
rect 16957 15105 16991 15139
rect 15945 15037 15979 15071
rect 23673 15037 23707 15071
rect 14013 14833 14047 14867
rect 15117 14833 15151 14867
rect 15485 14833 15519 14867
rect 16037 14833 16071 14867
rect 18889 14833 18923 14867
rect 19901 14833 19935 14867
rect 21373 14833 21407 14867
rect 21741 14833 21775 14867
rect 23765 14833 23799 14867
rect 24869 14833 24903 14867
rect 25513 14833 25547 14867
rect 25881 14833 25915 14867
rect 16497 14765 16531 14799
rect 22477 14765 22511 14799
rect 16681 14697 16715 14731
rect 19349 14697 19383 14731
rect 19533 14697 19567 14731
rect 20269 14697 20303 14731
rect 20729 14697 20763 14731
rect 23029 14697 23063 14731
rect 24317 14697 24351 14731
rect 15301 14629 15335 14663
rect 22845 14629 22879 14663
rect 24041 14629 24075 14663
rect 25329 14629 25363 14663
rect 16926 14561 16960 14595
rect 18705 14561 18739 14595
rect 13645 14493 13679 14527
rect 18061 14493 18095 14527
rect 18429 14493 18463 14527
rect 19257 14493 19291 14527
rect 20913 14493 20947 14527
rect 22385 14493 22419 14527
rect 22937 14493 22971 14527
rect 25145 14493 25179 14527
rect 13645 14289 13679 14323
rect 16957 14289 16991 14323
rect 19717 14289 19751 14323
rect 22569 14289 22603 14323
rect 22937 14289 22971 14323
rect 23489 14289 23523 14323
rect 24593 14289 24627 14323
rect 25329 14289 25363 14323
rect 21097 14221 21131 14255
rect 24133 14221 24167 14255
rect 13461 14153 13495 14187
rect 15577 14153 15611 14187
rect 15844 14153 15878 14187
rect 18604 14153 18638 14187
rect 20821 14153 20855 14187
rect 23857 14153 23891 14187
rect 25145 14153 25179 14187
rect 18337 14085 18371 14119
rect 15393 13949 15427 13983
rect 13461 13745 13495 13779
rect 16037 13745 16071 13779
rect 16405 13745 16439 13779
rect 16865 13745 16899 13779
rect 17693 13745 17727 13779
rect 18521 13745 18555 13779
rect 19533 13745 19567 13779
rect 20269 13745 20303 13779
rect 23857 13745 23891 13779
rect 24777 13745 24811 13779
rect 25605 13745 25639 13779
rect 17969 13677 18003 13711
rect 19993 13677 20027 13711
rect 20913 13677 20947 13711
rect 13001 13609 13035 13643
rect 15485 13609 15519 13643
rect 18981 13609 19015 13643
rect 19165 13609 19199 13643
rect 21465 13609 21499 13643
rect 25237 13609 25271 13643
rect 12725 13541 12759 13575
rect 15117 13541 15151 13575
rect 15301 13541 15335 13575
rect 16681 13541 16715 13575
rect 17233 13541 17267 13575
rect 18337 13541 18371 13575
rect 21373 13541 21407 13575
rect 21925 13541 21959 13575
rect 24593 13541 24627 13575
rect 18889 13473 18923 13507
rect 20729 13473 20763 13507
rect 21281 13473 21315 13507
rect 12633 13405 12667 13439
rect 18797 13201 18831 13235
rect 21833 13201 21867 13235
rect 24777 13201 24811 13235
rect 16957 13133 16991 13167
rect 16681 13065 16715 13099
rect 19625 13065 19659 13099
rect 19892 13065 19926 13099
rect 24593 13065 24627 13099
rect 12725 12997 12759 13031
rect 18245 12997 18279 13031
rect 13277 12861 13311 12895
rect 15393 12861 15427 12895
rect 21005 12861 21039 12895
rect 21373 12861 21407 12895
rect 13001 12657 13035 12691
rect 13185 12657 13219 12691
rect 15301 12657 15335 12691
rect 18061 12657 18095 12691
rect 19625 12657 19659 12691
rect 20637 12657 20671 12691
rect 22293 12657 22327 12691
rect 24225 12657 24259 12691
rect 25053 12657 25087 12691
rect 16773 12589 16807 12623
rect 18153 12589 18187 12623
rect 13737 12521 13771 12555
rect 15853 12521 15887 12555
rect 17325 12521 17359 12555
rect 18613 12521 18647 12555
rect 18705 12521 18739 12555
rect 20913 12521 20947 12555
rect 24685 12521 24719 12555
rect 13553 12453 13587 12487
rect 18521 12453 18555 12487
rect 19993 12453 20027 12487
rect 24041 12453 24075 12487
rect 12725 12385 12759 12419
rect 13645 12385 13679 12419
rect 15117 12385 15151 12419
rect 15669 12385 15703 12419
rect 21180 12385 21214 12419
rect 14749 12317 14783 12351
rect 15761 12317 15795 12351
rect 17693 12317 17727 12351
rect 16589 12113 16623 12147
rect 19533 12113 19567 12147
rect 20821 12113 20855 12147
rect 24777 12113 24811 12147
rect 13268 12045 13302 12079
rect 13001 11977 13035 12011
rect 15209 11977 15243 12011
rect 15465 11977 15499 12011
rect 18409 11977 18443 12011
rect 21189 11977 21223 12011
rect 21281 11977 21315 12011
rect 24593 11977 24627 12011
rect 18153 11909 18187 11943
rect 21373 11909 21407 11943
rect 14381 11773 14415 11807
rect 13921 11569 13955 11603
rect 14197 11569 14231 11603
rect 15025 11569 15059 11603
rect 15945 11569 15979 11603
rect 16589 11569 16623 11603
rect 18337 11569 18371 11603
rect 18889 11569 18923 11603
rect 20729 11569 20763 11603
rect 21465 11569 21499 11603
rect 24685 11569 24719 11603
rect 12541 11433 12575 11467
rect 15393 11433 15427 11467
rect 16681 11433 16715 11467
rect 19441 11433 19475 11467
rect 10333 11365 10367 11399
rect 11989 11365 12023 11399
rect 12357 11365 12391 11399
rect 16937 11365 16971 11399
rect 19349 11365 19383 11399
rect 21189 11365 21223 11399
rect 10149 11297 10183 11331
rect 10578 11297 10612 11331
rect 12808 11297 12842 11331
rect 11713 11229 11747 11263
rect 18061 11229 18095 11263
rect 18797 11229 18831 11263
rect 19257 11229 19291 11263
rect 10333 11025 10367 11059
rect 13093 11025 13127 11059
rect 15577 11025 15611 11059
rect 16773 11025 16807 11059
rect 18337 11025 18371 11059
rect 19349 11025 19383 11059
rect 24777 11025 24811 11059
rect 16037 10957 16071 10991
rect 18981 10957 19015 10991
rect 13461 10889 13495 10923
rect 15945 10889 15979 10923
rect 24593 10889 24627 10923
rect 13553 10821 13587 10855
rect 13737 10821 13771 10855
rect 16129 10821 16163 10855
rect 12725 10753 12759 10787
rect 13829 10481 13863 10515
rect 16037 10481 16071 10515
rect 16313 10481 16347 10515
rect 24501 10481 24535 10515
rect 13553 10413 13587 10447
rect 24777 10413 24811 10447
rect 24593 10277 24627 10311
rect 13185 10141 13219 10175
rect 15669 10141 15703 10175
rect 25237 10141 25271 10175
rect 24777 9937 24811 9971
rect 24593 9801 24627 9835
rect 24777 9325 24811 9359
rect 25237 9325 25271 9359
rect 24593 9189 24627 9223
rect 24501 9053 24535 9087
rect 24777 8849 24811 8883
rect 24593 8713 24627 8747
rect 24685 8305 24719 8339
rect 24593 7625 24627 7659
rect 24777 7489 24811 7523
rect 17785 7217 17819 7251
rect 24685 7217 24719 7251
rect 18245 7081 18279 7115
rect 17601 7013 17635 7047
rect 16405 6129 16439 6163
rect 16221 5925 16255 5959
rect 16865 5857 16899 5891
rect 15485 5041 15519 5075
rect 15301 4837 15335 4871
rect 15945 4769 15979 4803
rect 24593 3749 24627 3783
rect 24777 3613 24811 3647
rect 25237 3613 25271 3647
<< metal1 >>
rect 290 27132 296 27184
rect 348 27172 354 27184
rect 474 27172 480 27184
rect 348 27144 480 27172
rect 348 27132 354 27144
rect 474 27132 480 27144
rect 532 27132 538 27184
rect 1104 25314 26864 25336
rect 1104 25262 10315 25314
rect 10367 25262 10379 25314
rect 10431 25262 10443 25314
rect 10495 25262 10507 25314
rect 10559 25262 19648 25314
rect 19700 25262 19712 25314
rect 19764 25262 19776 25314
rect 19828 25262 19840 25314
rect 19892 25262 26864 25314
rect 1104 25240 26864 25262
rect 23017 25203 23075 25209
rect 23017 25169 23029 25203
rect 23063 25200 23075 25203
rect 23566 25200 23572 25212
rect 23063 25172 23572 25200
rect 23063 25169 23075 25172
rect 23017 25163 23075 25169
rect 23566 25160 23572 25172
rect 23624 25160 23630 25212
rect 24762 25200 24768 25212
rect 24723 25172 24768 25200
rect 24762 25160 24768 25172
rect 24820 25160 24826 25212
rect 22830 25064 22836 25076
rect 22791 25036 22836 25064
rect 22830 25024 22836 25036
rect 22888 25024 22894 25076
rect 24581 25067 24639 25073
rect 24581 25033 24593 25067
rect 24627 25064 24639 25067
rect 24627 25036 24808 25064
rect 24627 25033 24639 25036
rect 24581 25027 24639 25033
rect 24780 25008 24808 25036
rect 24762 24956 24768 25008
rect 24820 24956 24826 25008
rect 11422 24860 11428 24872
rect 11383 24832 11428 24860
rect 11422 24820 11428 24832
rect 11480 24820 11486 24872
rect 1104 24770 26864 24792
rect 1104 24718 5648 24770
rect 5700 24718 5712 24770
rect 5764 24718 5776 24770
rect 5828 24718 5840 24770
rect 5892 24718 14982 24770
rect 15034 24718 15046 24770
rect 15098 24718 15110 24770
rect 15162 24718 15174 24770
rect 15226 24718 24315 24770
rect 24367 24718 24379 24770
rect 24431 24718 24443 24770
rect 24495 24718 24507 24770
rect 24559 24718 26864 24770
rect 1104 24696 26864 24718
rect 22830 24548 22836 24600
rect 22888 24588 22894 24600
rect 22888 24560 23428 24588
rect 22888 24548 22894 24560
rect 11238 24480 11244 24532
rect 11296 24520 11302 24532
rect 11977 24523 12035 24529
rect 11977 24520 11989 24523
rect 11296 24492 11989 24520
rect 11296 24480 11302 24492
rect 11977 24489 11989 24492
rect 12023 24489 12035 24523
rect 11977 24483 12035 24489
rect 15286 24480 15292 24532
rect 15344 24520 15350 24532
rect 16206 24520 16212 24532
rect 15344 24492 16212 24520
rect 15344 24480 15350 24492
rect 16206 24480 16212 24492
rect 16264 24480 16270 24532
rect 18690 24480 18696 24532
rect 18748 24520 18754 24532
rect 19150 24520 19156 24532
rect 18748 24492 19156 24520
rect 18748 24480 18754 24492
rect 19150 24480 19156 24492
rect 19208 24480 19214 24532
rect 21358 24480 21364 24532
rect 21416 24520 21422 24532
rect 22002 24520 22008 24532
rect 21416 24492 22008 24520
rect 21416 24480 21422 24492
rect 22002 24480 22008 24492
rect 22060 24480 22066 24532
rect 23400 24520 23428 24560
rect 23477 24523 23535 24529
rect 23477 24520 23489 24523
rect 23400 24492 23489 24520
rect 23477 24489 23489 24492
rect 23523 24489 23535 24523
rect 23477 24483 23535 24489
rect 23750 24480 23756 24532
rect 23808 24520 23814 24532
rect 24670 24520 24676 24532
rect 23808 24492 24676 24520
rect 23808 24480 23814 24492
rect 24670 24480 24676 24492
rect 24728 24480 24734 24532
rect 11054 24412 11060 24464
rect 11112 24452 11118 24464
rect 11422 24452 11428 24464
rect 11112 24424 11428 24452
rect 11112 24412 11118 24424
rect 11422 24412 11428 24424
rect 11480 24452 11486 24464
rect 11885 24455 11943 24461
rect 11885 24452 11897 24455
rect 11480 24424 11897 24452
rect 11480 24412 11486 24424
rect 11885 24421 11897 24424
rect 11931 24421 11943 24455
rect 11885 24415 11943 24421
rect 20714 24412 20720 24464
rect 20772 24452 20778 24464
rect 21634 24452 21640 24464
rect 20772 24424 21640 24452
rect 20772 24412 20778 24424
rect 21634 24412 21640 24424
rect 21692 24412 21698 24464
rect 22554 24452 22560 24464
rect 22515 24424 22560 24452
rect 22554 24412 22560 24424
rect 22612 24452 22618 24464
rect 23109 24455 23167 24461
rect 23109 24452 23121 24455
rect 22612 24424 23121 24452
rect 22612 24412 22618 24424
rect 23109 24421 23121 24424
rect 23155 24421 23167 24455
rect 23109 24415 23167 24421
rect 23661 24455 23719 24461
rect 23661 24421 23673 24455
rect 23707 24452 23719 24455
rect 23842 24452 23848 24464
rect 23707 24424 23848 24452
rect 23707 24421 23719 24424
rect 23661 24415 23719 24421
rect 23842 24412 23848 24424
rect 23900 24412 23906 24464
rect 24210 24412 24216 24464
rect 24268 24452 24274 24464
rect 24949 24455 25007 24461
rect 24949 24452 24961 24455
rect 24268 24424 24961 24452
rect 24268 24412 24274 24424
rect 24949 24421 24961 24424
rect 24995 24452 25007 24455
rect 25501 24455 25559 24461
rect 25501 24452 25513 24455
rect 24995 24424 25513 24452
rect 24995 24421 25007 24424
rect 24949 24415 25007 24421
rect 25501 24421 25513 24424
rect 25547 24421 25559 24455
rect 25501 24415 25559 24421
rect 12342 24384 12348 24396
rect 11440 24356 12348 24384
rect 11238 24316 11244 24328
rect 11199 24288 11244 24316
rect 11238 24276 11244 24288
rect 11296 24276 11302 24328
rect 11440 24325 11468 24356
rect 12342 24344 12348 24356
rect 12400 24344 12406 24396
rect 23937 24387 23995 24393
rect 23937 24353 23949 24387
rect 23983 24384 23995 24387
rect 24670 24384 24676 24396
rect 23983 24356 24676 24384
rect 23983 24353 23995 24356
rect 23937 24347 23995 24353
rect 24670 24344 24676 24356
rect 24728 24344 24734 24396
rect 11425 24319 11483 24325
rect 11425 24285 11437 24319
rect 11471 24285 11483 24319
rect 11790 24316 11796 24328
rect 11751 24288 11796 24316
rect 11425 24279 11483 24285
rect 11790 24276 11796 24288
rect 11848 24276 11854 24328
rect 16485 24319 16543 24325
rect 16485 24285 16497 24319
rect 16531 24316 16543 24319
rect 16850 24316 16856 24328
rect 16531 24288 16856 24316
rect 16531 24285 16543 24288
rect 16485 24279 16543 24285
rect 16850 24276 16856 24288
rect 16908 24276 16914 24328
rect 17402 24316 17408 24328
rect 17363 24288 17408 24316
rect 17402 24276 17408 24288
rect 17460 24276 17466 24328
rect 22741 24319 22799 24325
rect 22741 24285 22753 24319
rect 22787 24316 22799 24319
rect 23382 24316 23388 24328
rect 22787 24288 23388 24316
rect 22787 24285 22799 24288
rect 22741 24279 22799 24285
rect 23382 24276 23388 24288
rect 23440 24276 23446 24328
rect 23842 24276 23848 24328
rect 23900 24316 23906 24328
rect 24397 24319 24455 24325
rect 24397 24316 24409 24319
rect 23900 24288 24409 24316
rect 23900 24276 23906 24288
rect 24397 24285 24409 24288
rect 24443 24285 24455 24319
rect 24762 24316 24768 24328
rect 24723 24288 24768 24316
rect 24397 24279 24455 24285
rect 24762 24276 24768 24288
rect 24820 24276 24826 24328
rect 25130 24316 25136 24328
rect 25091 24288 25136 24316
rect 25130 24276 25136 24288
rect 25188 24276 25194 24328
rect 1104 24226 26864 24248
rect 1104 24174 10315 24226
rect 10367 24174 10379 24226
rect 10431 24174 10443 24226
rect 10495 24174 10507 24226
rect 10559 24174 19648 24226
rect 19700 24174 19712 24226
rect 19764 24174 19776 24226
rect 19828 24174 19840 24226
rect 19892 24174 26864 24226
rect 1104 24152 26864 24174
rect 21545 24115 21603 24121
rect 21545 24081 21557 24115
rect 21591 24112 21603 24115
rect 22738 24112 22744 24124
rect 21591 24084 22744 24112
rect 21591 24081 21603 24084
rect 21545 24075 21603 24081
rect 22738 24072 22744 24084
rect 22796 24072 22802 24124
rect 23937 24047 23995 24053
rect 23937 24013 23949 24047
rect 23983 24044 23995 24047
rect 24210 24044 24216 24056
rect 23983 24016 24216 24044
rect 23983 24013 23995 24016
rect 23937 24007 23995 24013
rect 24210 24004 24216 24016
rect 24268 24004 24274 24056
rect 13170 23936 13176 23988
rect 13228 23976 13234 23988
rect 14165 23979 14223 23985
rect 14165 23976 14177 23979
rect 13228 23948 14177 23976
rect 13228 23936 13234 23948
rect 14165 23945 14177 23948
rect 14211 23976 14223 23979
rect 15102 23976 15108 23988
rect 14211 23948 15108 23976
rect 14211 23945 14223 23948
rect 14165 23939 14223 23945
rect 15102 23936 15108 23948
rect 15160 23936 15166 23988
rect 15470 23936 15476 23988
rect 15528 23976 15534 23988
rect 15930 23976 15936 23988
rect 15528 23948 15936 23976
rect 15528 23936 15534 23948
rect 15930 23936 15936 23948
rect 15988 23936 15994 23988
rect 16669 23979 16727 23985
rect 16669 23945 16681 23979
rect 16715 23976 16727 23979
rect 18138 23976 18144 23988
rect 16715 23948 18144 23976
rect 16715 23945 16727 23948
rect 16669 23939 16727 23945
rect 18138 23936 18144 23948
rect 18196 23936 18202 23988
rect 19242 23976 19248 23988
rect 19203 23948 19248 23976
rect 19242 23936 19248 23948
rect 19300 23936 19306 23988
rect 21082 23936 21088 23988
rect 21140 23976 21146 23988
rect 21361 23979 21419 23985
rect 21361 23976 21373 23979
rect 21140 23948 21373 23976
rect 21140 23936 21146 23948
rect 21361 23945 21373 23948
rect 21407 23976 21419 23979
rect 21913 23979 21971 23985
rect 21913 23976 21925 23979
rect 21407 23948 21925 23976
rect 21407 23945 21419 23948
rect 21361 23939 21419 23945
rect 21913 23945 21925 23948
rect 21959 23945 21971 23979
rect 21913 23939 21971 23945
rect 22278 23936 22284 23988
rect 22336 23976 22342 23988
rect 22465 23979 22523 23985
rect 22465 23976 22477 23979
rect 22336 23948 22477 23976
rect 22336 23936 22342 23948
rect 22465 23945 22477 23948
rect 22511 23976 22523 23979
rect 23017 23979 23075 23985
rect 23017 23976 23029 23979
rect 22511 23948 23029 23976
rect 22511 23945 22523 23948
rect 22465 23939 22523 23945
rect 23017 23945 23029 23948
rect 23063 23945 23075 23979
rect 23658 23976 23664 23988
rect 23619 23948 23664 23976
rect 23017 23939 23075 23945
rect 23658 23936 23664 23948
rect 23716 23936 23722 23988
rect 24670 23936 24676 23988
rect 24728 23976 24734 23988
rect 24949 23979 25007 23985
rect 24949 23976 24961 23979
rect 24728 23948 24961 23976
rect 24728 23936 24734 23948
rect 24949 23945 24961 23948
rect 24995 23945 25007 23979
rect 24949 23939 25007 23945
rect 13814 23868 13820 23920
rect 13872 23908 13878 23920
rect 13909 23911 13967 23917
rect 13909 23908 13921 23911
rect 13872 23880 13921 23908
rect 13872 23868 13878 23880
rect 13909 23877 13921 23880
rect 13955 23877 13967 23911
rect 13909 23871 13967 23877
rect 16114 23868 16120 23920
rect 16172 23908 16178 23920
rect 16761 23911 16819 23917
rect 16761 23908 16773 23911
rect 16172 23880 16773 23908
rect 16172 23868 16178 23880
rect 16761 23877 16773 23880
rect 16807 23877 16819 23911
rect 16761 23871 16819 23877
rect 16850 23868 16856 23920
rect 16908 23908 16914 23920
rect 16908 23880 16953 23908
rect 16908 23868 16914 23880
rect 18414 23868 18420 23920
rect 18472 23908 18478 23920
rect 19337 23911 19395 23917
rect 19337 23908 19349 23911
rect 18472 23880 19349 23908
rect 18472 23868 18478 23880
rect 19337 23877 19349 23880
rect 19383 23877 19395 23911
rect 19337 23871 19395 23877
rect 19521 23911 19579 23917
rect 19521 23877 19533 23911
rect 19567 23877 19579 23911
rect 19521 23871 19579 23877
rect 16209 23843 16267 23849
rect 16209 23809 16221 23843
rect 16255 23840 16267 23843
rect 16868 23840 16896 23868
rect 19426 23840 19432 23852
rect 16255 23812 16896 23840
rect 18340 23812 19432 23840
rect 16255 23809 16267 23812
rect 16209 23803 16267 23809
rect 18340 23784 18368 23812
rect 19426 23800 19432 23812
rect 19484 23840 19490 23852
rect 19536 23840 19564 23871
rect 19484 23812 19564 23840
rect 19484 23800 19490 23812
rect 19978 23800 19984 23852
rect 20036 23840 20042 23852
rect 20901 23843 20959 23849
rect 20901 23840 20913 23843
rect 20036 23812 20913 23840
rect 20036 23800 20042 23812
rect 20901 23809 20913 23812
rect 20947 23840 20959 23843
rect 21450 23840 21456 23852
rect 20947 23812 21456 23840
rect 20947 23809 20959 23812
rect 20901 23803 20959 23809
rect 21450 23800 21456 23812
rect 21508 23800 21514 23852
rect 22649 23843 22707 23849
rect 22649 23809 22661 23843
rect 22695 23840 22707 23843
rect 23290 23840 23296 23852
rect 22695 23812 23296 23840
rect 22695 23809 22707 23812
rect 22649 23803 22707 23809
rect 23290 23800 23296 23812
rect 23348 23800 23354 23852
rect 25130 23840 25136 23852
rect 25091 23812 25136 23840
rect 25130 23800 25136 23812
rect 25188 23800 25194 23852
rect 25222 23800 25228 23852
rect 25280 23840 25286 23852
rect 26142 23840 26148 23852
rect 25280 23812 26148 23840
rect 25280 23800 25286 23812
rect 26142 23800 26148 23812
rect 26200 23800 26206 23852
rect 11054 23732 11060 23784
rect 11112 23772 11118 23784
rect 11425 23775 11483 23781
rect 11425 23772 11437 23775
rect 11112 23744 11437 23772
rect 11112 23732 11118 23744
rect 11425 23741 11437 23744
rect 11471 23772 11483 23775
rect 11790 23772 11796 23784
rect 11471 23744 11796 23772
rect 11471 23741 11483 23744
rect 11425 23735 11483 23741
rect 11790 23732 11796 23744
rect 11848 23732 11854 23784
rect 13725 23775 13783 23781
rect 13725 23741 13737 23775
rect 13771 23772 13783 23775
rect 14274 23772 14280 23784
rect 13771 23744 14280 23772
rect 13771 23741 13783 23744
rect 13725 23735 13783 23741
rect 14274 23732 14280 23744
rect 14332 23772 14338 23784
rect 15289 23775 15347 23781
rect 15289 23772 15301 23775
rect 14332 23744 15301 23772
rect 14332 23732 14338 23744
rect 15289 23741 15301 23744
rect 15335 23741 15347 23775
rect 16298 23772 16304 23784
rect 16259 23744 16304 23772
rect 15289 23735 15347 23741
rect 16298 23732 16304 23744
rect 16356 23732 16362 23784
rect 18322 23772 18328 23784
rect 18283 23744 18328 23772
rect 18322 23732 18328 23744
rect 18380 23732 18386 23784
rect 18690 23772 18696 23784
rect 18651 23744 18696 23772
rect 18690 23732 18696 23744
rect 18748 23732 18754 23784
rect 18877 23775 18935 23781
rect 18877 23741 18889 23775
rect 18923 23772 18935 23775
rect 20530 23772 20536 23784
rect 18923 23744 20536 23772
rect 18923 23741 18935 23744
rect 18877 23735 18935 23741
rect 20530 23732 20536 23744
rect 20588 23732 20594 23784
rect 24210 23732 24216 23784
rect 24268 23772 24274 23784
rect 24397 23775 24455 23781
rect 24397 23772 24409 23775
rect 24268 23744 24409 23772
rect 24268 23732 24274 23744
rect 24397 23741 24409 23744
rect 24443 23741 24455 23775
rect 24397 23735 24455 23741
rect 1104 23682 26864 23704
rect 1104 23630 5648 23682
rect 5700 23630 5712 23682
rect 5764 23630 5776 23682
rect 5828 23630 5840 23682
rect 5892 23630 14982 23682
rect 15034 23630 15046 23682
rect 15098 23630 15110 23682
rect 15162 23630 15174 23682
rect 15226 23630 24315 23682
rect 24367 23630 24379 23682
rect 24431 23630 24443 23682
rect 24495 23630 24507 23682
rect 24559 23630 26864 23682
rect 1104 23608 26864 23630
rect 13170 23568 13176 23580
rect 13131 23540 13176 23568
rect 13170 23528 13176 23540
rect 13228 23528 13234 23580
rect 13446 23568 13452 23580
rect 13407 23540 13452 23568
rect 13446 23528 13452 23540
rect 13504 23568 13510 23580
rect 13504 23540 14136 23568
rect 13504 23528 13510 23540
rect 14108 23441 14136 23540
rect 16114 23528 16120 23580
rect 16172 23568 16178 23580
rect 16209 23571 16267 23577
rect 16209 23568 16221 23571
rect 16172 23540 16221 23568
rect 16172 23528 16178 23540
rect 16209 23537 16221 23540
rect 16255 23537 16267 23571
rect 18138 23568 18144 23580
rect 18099 23540 18144 23568
rect 16209 23531 16267 23537
rect 18138 23528 18144 23540
rect 18196 23528 18202 23580
rect 18414 23568 18420 23580
rect 18375 23540 18420 23568
rect 18414 23528 18420 23540
rect 18472 23528 18478 23580
rect 19978 23568 19984 23580
rect 19939 23540 19984 23568
rect 19978 23528 19984 23540
rect 20036 23528 20042 23580
rect 20901 23571 20959 23577
rect 20901 23537 20913 23571
rect 20947 23568 20959 23571
rect 23658 23568 23664 23580
rect 20947 23540 23664 23568
rect 20947 23537 20959 23540
rect 20901 23531 20959 23537
rect 23658 23528 23664 23540
rect 23716 23528 23722 23580
rect 24670 23528 24676 23580
rect 24728 23568 24734 23580
rect 24949 23571 25007 23577
rect 24949 23568 24961 23571
rect 24728 23540 24961 23568
rect 24728 23528 24734 23540
rect 24949 23537 24961 23540
rect 24995 23537 25007 23571
rect 24949 23531 25007 23537
rect 22094 23460 22100 23512
rect 22152 23500 22158 23512
rect 22152 23472 22197 23500
rect 22152 23460 22158 23472
rect 14093 23435 14151 23441
rect 14093 23401 14105 23435
rect 14139 23401 14151 23435
rect 14274 23432 14280 23444
rect 14235 23404 14280 23432
rect 14093 23395 14151 23401
rect 14274 23392 14280 23404
rect 14332 23392 14338 23444
rect 20530 23392 20536 23444
rect 20588 23432 20594 23444
rect 21361 23435 21419 23441
rect 21361 23432 21373 23435
rect 20588 23404 21373 23432
rect 20588 23392 20594 23404
rect 21361 23401 21373 23404
rect 21407 23401 21419 23435
rect 21361 23395 21419 23401
rect 21450 23392 21456 23444
rect 21508 23432 21514 23444
rect 21508 23404 21553 23432
rect 21508 23392 21514 23404
rect 11330 23364 11336 23376
rect 11243 23336 11336 23364
rect 11330 23324 11336 23336
rect 11388 23364 11394 23376
rect 11425 23367 11483 23373
rect 11425 23364 11437 23367
rect 11388 23336 11437 23364
rect 11388 23324 11394 23336
rect 11425 23333 11437 23336
rect 11471 23364 11483 23367
rect 11471 23336 12388 23364
rect 11471 23333 11483 23336
rect 11425 23327 11483 23333
rect 10965 23299 11023 23305
rect 10965 23265 10977 23299
rect 11011 23296 11023 23299
rect 11670 23299 11728 23305
rect 11670 23296 11682 23299
rect 11011 23268 11682 23296
rect 11011 23265 11023 23268
rect 10965 23259 11023 23265
rect 11670 23265 11682 23268
rect 11716 23296 11728 23299
rect 12158 23296 12164 23308
rect 11716 23268 12164 23296
rect 11716 23265 11728 23268
rect 11670 23259 11728 23265
rect 12158 23256 12164 23268
rect 12216 23256 12222 23308
rect 12360 23296 12388 23336
rect 13814 23324 13820 23376
rect 13872 23324 13878 23376
rect 16393 23367 16451 23373
rect 16393 23364 16405 23367
rect 15948 23336 16405 23364
rect 13832 23296 13860 23324
rect 15948 23308 15976 23336
rect 16393 23333 16405 23336
rect 16439 23364 16451 23367
rect 18138 23364 18144 23376
rect 16439 23336 18144 23364
rect 16439 23333 16451 23336
rect 16393 23327 16451 23333
rect 18138 23324 18144 23336
rect 18196 23364 18202 23376
rect 18601 23367 18659 23373
rect 18601 23364 18613 23367
rect 18196 23336 18613 23364
rect 18196 23324 18202 23336
rect 18601 23333 18613 23336
rect 18647 23364 18659 23367
rect 18690 23364 18696 23376
rect 18647 23336 18696 23364
rect 18647 23333 18659 23336
rect 18601 23327 18659 23333
rect 18690 23324 18696 23336
rect 18748 23324 18754 23376
rect 19426 23324 19432 23376
rect 19484 23364 19490 23376
rect 20257 23367 20315 23373
rect 20257 23364 20269 23367
rect 19484 23336 20269 23364
rect 19484 23324 19490 23336
rect 20257 23333 20269 23336
rect 20303 23333 20315 23367
rect 22112 23364 22140 23460
rect 22830 23392 22836 23444
rect 22888 23432 22894 23444
rect 23109 23435 23167 23441
rect 23109 23432 23121 23435
rect 22888 23404 23121 23432
rect 22888 23392 22894 23404
rect 23109 23401 23121 23404
rect 23155 23401 23167 23435
rect 23109 23395 23167 23401
rect 24397 23435 24455 23441
rect 24397 23401 24409 23435
rect 24443 23432 24455 23435
rect 24762 23432 24768 23444
rect 24443 23404 24768 23432
rect 24443 23401 24455 23404
rect 24397 23395 24455 23401
rect 24762 23392 24768 23404
rect 24820 23392 24826 23444
rect 22925 23367 22983 23373
rect 22925 23364 22937 23367
rect 22112 23336 22937 23364
rect 20257 23327 20315 23333
rect 22925 23333 22937 23336
rect 22971 23333 22983 23367
rect 22925 23327 22983 23333
rect 23658 23324 23664 23376
rect 23716 23364 23722 23376
rect 24121 23367 24179 23373
rect 24121 23364 24133 23367
rect 23716 23336 24133 23364
rect 23716 23324 23722 23336
rect 24121 23333 24133 23336
rect 24167 23364 24179 23367
rect 24210 23364 24216 23376
rect 24167 23336 24216 23364
rect 24167 23333 24179 23336
rect 24121 23327 24179 23333
rect 24210 23324 24216 23336
rect 24268 23324 24274 23376
rect 14737 23299 14795 23305
rect 14737 23296 14749 23299
rect 12360 23268 14749 23296
rect 14737 23265 14749 23268
rect 14783 23296 14795 23299
rect 15930 23296 15936 23308
rect 14783 23268 15936 23296
rect 14783 23265 14795 23268
rect 14737 23259 14795 23265
rect 15930 23256 15936 23268
rect 15988 23256 15994 23308
rect 16660 23299 16718 23305
rect 16660 23265 16672 23299
rect 16706 23296 16718 23299
rect 16850 23296 16856 23308
rect 16706 23268 16856 23296
rect 16706 23265 16718 23268
rect 16660 23259 16718 23265
rect 16850 23256 16856 23268
rect 16908 23296 16914 23308
rect 17310 23296 17316 23308
rect 16908 23268 17316 23296
rect 16908 23256 16914 23268
rect 17310 23256 17316 23268
rect 17368 23256 17374 23308
rect 18322 23256 18328 23308
rect 18380 23296 18386 23308
rect 18846 23299 18904 23305
rect 18846 23296 18858 23299
rect 18380 23268 18858 23296
rect 18380 23256 18386 23268
rect 18846 23265 18858 23268
rect 18892 23265 18904 23299
rect 18846 23259 18904 23265
rect 19334 23256 19340 23308
rect 19392 23296 19398 23308
rect 20530 23296 20536 23308
rect 19392 23268 20536 23296
rect 19392 23256 19398 23268
rect 20530 23256 20536 23268
rect 20588 23256 20594 23308
rect 22370 23296 22376 23308
rect 22331 23268 22376 23296
rect 22370 23256 22376 23268
rect 22428 23296 22434 23308
rect 23017 23299 23075 23305
rect 23017 23296 23029 23299
rect 22428 23268 23029 23296
rect 22428 23256 22434 23268
rect 23017 23265 23029 23268
rect 23063 23265 23075 23299
rect 23017 23259 23075 23265
rect 12250 23188 12256 23240
rect 12308 23228 12314 23240
rect 12805 23231 12863 23237
rect 12805 23228 12817 23231
rect 12308 23200 12817 23228
rect 12308 23188 12314 23200
rect 12805 23197 12817 23200
rect 12851 23197 12863 23231
rect 12805 23191 12863 23197
rect 13633 23231 13691 23237
rect 13633 23197 13645 23231
rect 13679 23228 13691 23231
rect 13814 23228 13820 23240
rect 13679 23200 13820 23228
rect 13679 23197 13691 23200
rect 13633 23191 13691 23197
rect 13814 23188 13820 23200
rect 13872 23188 13878 23240
rect 13998 23228 14004 23240
rect 13959 23200 14004 23228
rect 13998 23188 14004 23200
rect 14056 23188 14062 23240
rect 15286 23228 15292 23240
rect 15247 23200 15292 23228
rect 15286 23188 15292 23200
rect 15344 23188 15350 23240
rect 17218 23188 17224 23240
rect 17276 23228 17282 23240
rect 17773 23231 17831 23237
rect 17773 23228 17785 23231
rect 17276 23200 17785 23228
rect 17276 23188 17282 23200
rect 17773 23197 17785 23200
rect 17819 23197 17831 23231
rect 20714 23228 20720 23240
rect 20675 23200 20720 23228
rect 17773 23191 17831 23197
rect 20714 23188 20720 23200
rect 20772 23228 20778 23240
rect 21269 23231 21327 23237
rect 21269 23228 21281 23231
rect 20772 23200 21281 23228
rect 20772 23188 20778 23200
rect 21269 23197 21281 23200
rect 21315 23197 21327 23231
rect 21269 23191 21327 23197
rect 22557 23231 22615 23237
rect 22557 23197 22569 23231
rect 22603 23228 22615 23231
rect 23566 23228 23572 23240
rect 22603 23200 23572 23228
rect 22603 23197 22615 23200
rect 22557 23191 22615 23197
rect 23566 23188 23572 23200
rect 23624 23188 23630 23240
rect 1104 23138 26864 23160
rect 1104 23086 10315 23138
rect 10367 23086 10379 23138
rect 10431 23086 10443 23138
rect 10495 23086 10507 23138
rect 10559 23086 19648 23138
rect 19700 23086 19712 23138
rect 19764 23086 19776 23138
rect 19828 23086 19840 23138
rect 19892 23086 26864 23138
rect 1104 23064 26864 23086
rect 9769 23027 9827 23033
rect 9769 22993 9781 23027
rect 9815 23024 9827 23027
rect 10962 23024 10968 23036
rect 9815 22996 10968 23024
rect 9815 22993 9827 22996
rect 9769 22987 9827 22993
rect 10962 22984 10968 22996
rect 11020 22984 11026 23036
rect 11054 22984 11060 23036
rect 11112 23024 11118 23036
rect 11241 23027 11299 23033
rect 11241 23024 11253 23027
rect 11112 22996 11253 23024
rect 11112 22984 11118 22996
rect 11241 22993 11253 22996
rect 11287 23024 11299 23027
rect 11882 23024 11888 23036
rect 11287 22996 11888 23024
rect 11287 22993 11299 22996
rect 11241 22987 11299 22993
rect 11882 22984 11888 22996
rect 11940 22984 11946 23036
rect 15194 22984 15200 23036
rect 15252 23024 15258 23036
rect 15289 23027 15347 23033
rect 15289 23024 15301 23027
rect 15252 22996 15301 23024
rect 15252 22984 15258 22996
rect 15289 22993 15301 22996
rect 15335 22993 15347 23027
rect 15289 22987 15347 22993
rect 16761 23027 16819 23033
rect 16761 22993 16773 23027
rect 16807 23024 16819 23027
rect 17402 23024 17408 23036
rect 16807 22996 17408 23024
rect 16807 22993 16819 22996
rect 16761 22987 16819 22993
rect 17402 22984 17408 22996
rect 17460 22984 17466 23036
rect 19426 23024 19432 23036
rect 19387 22996 19432 23024
rect 19426 22984 19432 22996
rect 19484 22984 19490 23036
rect 23566 22984 23572 23036
rect 23624 23024 23630 23036
rect 24118 23024 24124 23036
rect 23624 22996 24124 23024
rect 23624 22984 23630 22996
rect 24118 22984 24124 22996
rect 24176 22984 24182 23036
rect 25406 23024 25412 23036
rect 25367 22996 25412 23024
rect 25406 22984 25412 22996
rect 25464 22984 25470 23036
rect 14176 22959 14234 22965
rect 14176 22925 14188 22959
rect 14222 22956 14234 22959
rect 14274 22956 14280 22968
rect 14222 22928 14280 22956
rect 14222 22925 14234 22928
rect 14176 22919 14234 22925
rect 14274 22916 14280 22928
rect 14332 22916 14338 22968
rect 15657 22959 15715 22965
rect 15657 22925 15669 22959
rect 15703 22956 15715 22959
rect 16298 22956 16304 22968
rect 15703 22928 16304 22956
rect 15703 22925 15715 22928
rect 15657 22919 15715 22925
rect 16298 22916 16304 22928
rect 16356 22956 16362 22968
rect 16853 22959 16911 22965
rect 16853 22956 16865 22959
rect 16356 22928 16865 22956
rect 16356 22916 16362 22928
rect 16853 22925 16865 22928
rect 16899 22925 16911 22959
rect 16853 22919 16911 22925
rect 19334 22916 19340 22968
rect 19392 22956 19398 22968
rect 19705 22959 19763 22965
rect 19705 22956 19717 22959
rect 19392 22928 19717 22956
rect 19392 22916 19398 22928
rect 19705 22925 19717 22928
rect 19751 22956 19763 22959
rect 20901 22959 20959 22965
rect 20901 22956 20913 22959
rect 19751 22928 20913 22956
rect 19751 22925 19763 22928
rect 19705 22919 19763 22925
rect 20901 22925 20913 22928
rect 20947 22956 20959 22959
rect 21174 22956 21180 22968
rect 20947 22928 21180 22956
rect 20947 22925 20959 22928
rect 20901 22919 20959 22925
rect 21174 22916 21180 22928
rect 21232 22916 21238 22968
rect 24029 22959 24087 22965
rect 24029 22925 24041 22959
rect 24075 22956 24087 22959
rect 24210 22956 24216 22968
rect 24075 22928 24216 22956
rect 24075 22925 24087 22928
rect 24029 22919 24087 22925
rect 24210 22916 24216 22928
rect 24268 22916 24274 22968
rect 11146 22888 11152 22900
rect 11107 22860 11152 22888
rect 11146 22848 11152 22860
rect 11204 22848 11210 22900
rect 12434 22848 12440 22900
rect 12492 22888 12498 22900
rect 12986 22888 12992 22900
rect 12492 22860 12992 22888
rect 12492 22848 12498 22860
rect 12986 22848 12992 22860
rect 13044 22848 13050 22900
rect 18322 22897 18328 22900
rect 18305 22891 18328 22897
rect 18305 22888 18317 22891
rect 17236 22860 18317 22888
rect 17236 22832 17264 22860
rect 18305 22857 18317 22860
rect 18380 22888 18386 22900
rect 18380 22860 18453 22888
rect 18305 22851 18328 22857
rect 18322 22848 18328 22851
rect 18380 22848 18386 22860
rect 20346 22848 20352 22900
rect 20404 22888 20410 22900
rect 21358 22897 21364 22900
rect 21341 22891 21364 22897
rect 21341 22888 21353 22891
rect 20404 22860 21353 22888
rect 20404 22848 20410 22860
rect 21341 22857 21353 22860
rect 21416 22888 21422 22900
rect 25225 22891 25283 22897
rect 21416 22860 21489 22888
rect 21341 22851 21364 22857
rect 21358 22848 21364 22851
rect 21416 22848 21422 22860
rect 25225 22857 25237 22891
rect 25271 22888 25283 22891
rect 25682 22888 25688 22900
rect 25271 22860 25688 22888
rect 25271 22857 25283 22860
rect 25225 22851 25283 22857
rect 25682 22848 25688 22860
rect 25740 22848 25746 22900
rect 11425 22823 11483 22829
rect 11425 22789 11437 22823
rect 11471 22820 11483 22823
rect 11606 22820 11612 22832
rect 11471 22792 11612 22820
rect 11471 22789 11483 22792
rect 11425 22783 11483 22789
rect 11606 22780 11612 22792
rect 11664 22820 11670 22832
rect 12250 22820 12256 22832
rect 11664 22792 12256 22820
rect 11664 22780 11670 22792
rect 12250 22780 12256 22792
rect 12308 22780 12314 22832
rect 12713 22823 12771 22829
rect 12713 22789 12725 22823
rect 12759 22820 12771 22823
rect 13722 22820 13728 22832
rect 12759 22792 13728 22820
rect 12759 22789 12771 22792
rect 12713 22783 12771 22789
rect 13722 22780 13728 22792
rect 13780 22780 13786 22832
rect 13909 22823 13967 22829
rect 13909 22789 13921 22823
rect 13955 22789 13967 22823
rect 13909 22783 13967 22789
rect 17037 22823 17095 22829
rect 17037 22789 17049 22823
rect 17083 22820 17095 22823
rect 17218 22820 17224 22832
rect 17083 22792 17224 22820
rect 17083 22789 17095 22792
rect 17037 22783 17095 22789
rect 10781 22755 10839 22761
rect 10781 22721 10793 22755
rect 10827 22752 10839 22755
rect 10870 22752 10876 22764
rect 10827 22724 10876 22752
rect 10827 22721 10839 22724
rect 10781 22715 10839 22721
rect 10870 22712 10876 22724
rect 10928 22712 10934 22764
rect 13722 22684 13728 22696
rect 13683 22656 13728 22684
rect 13722 22644 13728 22656
rect 13780 22644 13786 22696
rect 13924 22684 13952 22783
rect 17218 22780 17224 22792
rect 17276 22780 17282 22832
rect 18046 22820 18052 22832
rect 18007 22792 18052 22820
rect 18046 22780 18052 22792
rect 18104 22780 18110 22832
rect 20990 22780 20996 22832
rect 21048 22820 21054 22832
rect 21085 22823 21143 22829
rect 21085 22820 21097 22823
rect 21048 22792 21097 22820
rect 21048 22780 21054 22792
rect 21085 22789 21097 22792
rect 21131 22789 21143 22823
rect 21085 22783 21143 22789
rect 23934 22780 23940 22832
rect 23992 22820 23998 22832
rect 24213 22823 24271 22829
rect 24213 22820 24225 22823
rect 23992 22792 24225 22820
rect 23992 22780 23998 22792
rect 24213 22789 24225 22792
rect 24259 22789 24271 22823
rect 24213 22783 24271 22789
rect 16390 22752 16396 22764
rect 16351 22724 16396 22752
rect 16390 22712 16396 22724
rect 16448 22712 16454 22764
rect 14090 22684 14096 22696
rect 13924 22656 14096 22684
rect 14090 22644 14096 22656
rect 14148 22644 14154 22696
rect 16022 22684 16028 22696
rect 15983 22656 16028 22684
rect 16022 22644 16028 22656
rect 16080 22644 16086 22696
rect 20438 22644 20444 22696
rect 20496 22684 20502 22696
rect 20533 22687 20591 22693
rect 20533 22684 20545 22687
rect 20496 22656 20545 22684
rect 20496 22644 20502 22656
rect 20533 22653 20545 22656
rect 20579 22653 20591 22687
rect 22462 22684 22468 22696
rect 22423 22656 22468 22684
rect 20533 22647 20591 22653
rect 22462 22644 22468 22656
rect 22520 22644 22526 22696
rect 22830 22684 22836 22696
rect 22791 22656 22836 22684
rect 22830 22644 22836 22656
rect 22888 22644 22894 22696
rect 23661 22687 23719 22693
rect 23661 22653 23673 22687
rect 23707 22684 23719 22687
rect 24854 22684 24860 22696
rect 23707 22656 24860 22684
rect 23707 22653 23719 22656
rect 23661 22647 23719 22653
rect 24854 22644 24860 22656
rect 24912 22644 24918 22696
rect 1104 22594 26864 22616
rect 1104 22542 5648 22594
rect 5700 22542 5712 22594
rect 5764 22542 5776 22594
rect 5828 22542 5840 22594
rect 5892 22542 14982 22594
rect 15034 22542 15046 22594
rect 15098 22542 15110 22594
rect 15162 22542 15174 22594
rect 15226 22542 24315 22594
rect 24367 22542 24379 22594
rect 24431 22542 24443 22594
rect 24495 22542 24507 22594
rect 24559 22542 26864 22594
rect 1104 22520 26864 22542
rect 10873 22483 10931 22489
rect 10873 22449 10885 22483
rect 10919 22480 10931 22483
rect 11054 22480 11060 22492
rect 10919 22452 11060 22480
rect 10919 22449 10931 22452
rect 10873 22443 10931 22449
rect 11054 22440 11060 22452
rect 11112 22440 11118 22492
rect 12710 22480 12716 22492
rect 12671 22452 12716 22480
rect 12710 22440 12716 22452
rect 12768 22440 12774 22492
rect 12986 22480 12992 22492
rect 12947 22452 12992 22480
rect 12986 22440 12992 22452
rect 13044 22440 13050 22492
rect 14274 22480 14280 22492
rect 14235 22452 14280 22480
rect 14274 22440 14280 22452
rect 14332 22440 14338 22492
rect 17310 22480 17316 22492
rect 17271 22452 17316 22480
rect 17310 22440 17316 22452
rect 17368 22440 17374 22492
rect 17402 22440 17408 22492
rect 17460 22480 17466 22492
rect 17589 22483 17647 22489
rect 17589 22480 17601 22483
rect 17460 22452 17601 22480
rect 17460 22440 17466 22452
rect 17589 22449 17601 22452
rect 17635 22449 17647 22483
rect 18138 22480 18144 22492
rect 18099 22452 18144 22480
rect 17589 22443 17647 22449
rect 18138 22440 18144 22452
rect 18196 22440 18202 22492
rect 18322 22440 18328 22492
rect 18380 22480 18386 22492
rect 18417 22483 18475 22489
rect 18417 22480 18429 22483
rect 18380 22452 18429 22480
rect 18380 22440 18386 22452
rect 18417 22449 18429 22452
rect 18463 22449 18475 22483
rect 20346 22480 20352 22492
rect 20307 22452 20352 22480
rect 18417 22443 18475 22449
rect 20346 22440 20352 22452
rect 20404 22440 20410 22492
rect 20990 22440 20996 22492
rect 21048 22480 21054 22492
rect 22005 22483 22063 22489
rect 22005 22480 22017 22483
rect 21048 22452 22017 22480
rect 21048 22440 21054 22452
rect 22005 22449 22017 22452
rect 22051 22480 22063 22483
rect 22465 22483 22523 22489
rect 22465 22480 22477 22483
rect 22051 22452 22477 22480
rect 22051 22449 22063 22452
rect 22005 22443 22063 22449
rect 22465 22449 22477 22452
rect 22511 22480 22523 22483
rect 23198 22480 23204 22492
rect 22511 22452 23204 22480
rect 22511 22449 22523 22452
rect 22465 22443 22523 22449
rect 11241 22347 11299 22353
rect 11241 22313 11253 22347
rect 11287 22344 11299 22347
rect 11330 22344 11336 22356
rect 11287 22316 11336 22344
rect 11287 22313 11299 22316
rect 11241 22307 11299 22313
rect 11330 22304 11336 22316
rect 11388 22304 11394 22356
rect 14001 22347 14059 22353
rect 14001 22313 14013 22347
rect 14047 22344 14059 22347
rect 14090 22344 14096 22356
rect 14047 22316 14096 22344
rect 14047 22313 14059 22316
rect 14001 22307 14059 22313
rect 14090 22304 14096 22316
rect 14148 22344 14154 22356
rect 15378 22344 15384 22356
rect 14148 22316 15384 22344
rect 14148 22304 14154 22316
rect 15378 22304 15384 22316
rect 15436 22344 15442 22356
rect 15841 22347 15899 22353
rect 15841 22344 15853 22347
rect 15436 22316 15853 22344
rect 15436 22304 15442 22316
rect 15841 22313 15853 22316
rect 15887 22344 15899 22347
rect 15930 22344 15936 22356
rect 15887 22316 15936 22344
rect 15887 22313 15899 22316
rect 15841 22307 15899 22313
rect 15930 22304 15936 22316
rect 15988 22304 15994 22356
rect 19521 22347 19579 22353
rect 19521 22313 19533 22347
rect 19567 22344 19579 22347
rect 20622 22344 20628 22356
rect 19567 22316 20628 22344
rect 19567 22313 19579 22316
rect 19521 22307 19579 22313
rect 20622 22304 20628 22316
rect 20680 22304 20686 22356
rect 21453 22347 21511 22353
rect 21453 22313 21465 22347
rect 21499 22344 21511 22347
rect 22462 22344 22468 22356
rect 21499 22316 22468 22344
rect 21499 22313 21511 22316
rect 21453 22307 21511 22313
rect 11146 22236 11152 22288
rect 11204 22236 11210 22288
rect 11606 22285 11612 22288
rect 11600 22276 11612 22285
rect 11567 22248 11612 22276
rect 11600 22239 11612 22248
rect 11606 22236 11612 22239
rect 11664 22236 11670 22288
rect 16022 22236 16028 22288
rect 16080 22276 16086 22288
rect 16189 22279 16247 22285
rect 16189 22276 16201 22279
rect 16080 22248 16201 22276
rect 16080 22236 16086 22248
rect 16189 22245 16201 22248
rect 16235 22276 16247 22279
rect 16482 22276 16488 22288
rect 16235 22248 16488 22276
rect 16235 22245 16247 22248
rect 16189 22239 16247 22245
rect 16482 22236 16488 22248
rect 16540 22236 16546 22288
rect 20438 22236 20444 22288
rect 20496 22276 20502 22288
rect 21468 22276 21496 22307
rect 22462 22304 22468 22316
rect 22520 22304 22526 22356
rect 22572 22353 22600 22452
rect 23198 22440 23204 22452
rect 23256 22440 23262 22492
rect 23934 22480 23940 22492
rect 23895 22452 23940 22480
rect 23934 22440 23940 22452
rect 23992 22440 23998 22492
rect 24118 22440 24124 22492
rect 24176 22480 24182 22492
rect 24581 22483 24639 22489
rect 24581 22480 24593 22483
rect 24176 22452 24593 22480
rect 24176 22440 24182 22452
rect 24581 22449 24593 22452
rect 24627 22449 24639 22483
rect 24581 22443 24639 22449
rect 22557 22347 22615 22353
rect 22557 22313 22569 22347
rect 22603 22313 22615 22347
rect 22557 22307 22615 22313
rect 24762 22276 24768 22288
rect 20496 22248 21496 22276
rect 24723 22248 24768 22276
rect 20496 22236 20502 22248
rect 24762 22236 24768 22248
rect 24820 22276 24826 22288
rect 25317 22279 25375 22285
rect 25317 22276 25329 22279
rect 24820 22248 25329 22276
rect 24820 22236 24826 22248
rect 25317 22245 25329 22248
rect 25363 22245 25375 22279
rect 25317 22239 25375 22245
rect 10505 22211 10563 22217
rect 10505 22177 10517 22211
rect 10551 22208 10563 22211
rect 11164 22208 11192 22236
rect 11790 22208 11796 22220
rect 10551 22180 11796 22208
rect 10551 22177 10563 22180
rect 10505 22171 10563 22177
rect 11790 22168 11796 22180
rect 11848 22168 11854 22220
rect 15562 22168 15568 22220
rect 15620 22208 15626 22220
rect 16040 22208 16068 22236
rect 20714 22208 20720 22220
rect 15620 22180 16068 22208
rect 20675 22180 20720 22208
rect 15620 22168 15626 22180
rect 20714 22168 20720 22180
rect 20772 22208 20778 22220
rect 22830 22217 22836 22220
rect 21361 22211 21419 22217
rect 21361 22208 21373 22211
rect 20772 22180 21373 22208
rect 20772 22168 20778 22180
rect 21361 22177 21373 22180
rect 21407 22177 21419 22211
rect 22824 22208 22836 22217
rect 22743 22180 22836 22208
rect 21361 22171 21419 22177
rect 22824 22171 22836 22180
rect 22888 22208 22894 22220
rect 23382 22208 23388 22220
rect 22888 22180 23388 22208
rect 22830 22168 22836 22171
rect 22888 22168 22894 22180
rect 23382 22168 23388 22180
rect 23440 22168 23446 22220
rect 20898 22140 20904 22152
rect 20859 22112 20904 22140
rect 20898 22100 20904 22112
rect 20956 22100 20962 22152
rect 21174 22100 21180 22152
rect 21232 22140 21238 22152
rect 21269 22143 21327 22149
rect 21269 22140 21281 22143
rect 21232 22112 21281 22140
rect 21232 22100 21238 22112
rect 21269 22109 21281 22112
rect 21315 22140 21327 22143
rect 21726 22140 21732 22152
rect 21315 22112 21732 22140
rect 21315 22109 21327 22112
rect 21269 22103 21327 22109
rect 21726 22100 21732 22112
rect 21784 22100 21790 22152
rect 24210 22140 24216 22152
rect 24171 22112 24216 22140
rect 24210 22100 24216 22112
rect 24268 22100 24274 22152
rect 24946 22140 24952 22152
rect 24907 22112 24952 22140
rect 24946 22100 24952 22112
rect 25004 22100 25010 22152
rect 25682 22140 25688 22152
rect 25643 22112 25688 22140
rect 25682 22100 25688 22112
rect 25740 22100 25746 22152
rect 1104 22050 26864 22072
rect 1104 21998 10315 22050
rect 10367 21998 10379 22050
rect 10431 21998 10443 22050
rect 10495 21998 10507 22050
rect 10559 21998 19648 22050
rect 19700 21998 19712 22050
rect 19764 21998 19776 22050
rect 19828 21998 19840 22050
rect 19892 21998 26864 22050
rect 1104 21976 26864 21998
rect 11425 21939 11483 21945
rect 11425 21905 11437 21939
rect 11471 21936 11483 21939
rect 11606 21936 11612 21948
rect 11471 21908 11612 21936
rect 11471 21905 11483 21908
rect 11425 21899 11483 21905
rect 474 21828 480 21880
rect 532 21828 538 21880
rect 492 21744 520 21828
rect 10873 21803 10931 21809
rect 10873 21769 10885 21803
rect 10919 21800 10931 21803
rect 11440 21800 11468 21899
rect 11606 21896 11612 21908
rect 11664 21896 11670 21948
rect 14366 21896 14372 21948
rect 14424 21936 14430 21948
rect 14645 21939 14703 21945
rect 14645 21936 14657 21939
rect 14424 21908 14657 21936
rect 14424 21896 14430 21908
rect 14645 21905 14657 21908
rect 14691 21936 14703 21939
rect 15102 21936 15108 21948
rect 14691 21908 15108 21936
rect 14691 21905 14703 21908
rect 14645 21899 14703 21905
rect 15102 21896 15108 21908
rect 15160 21896 15166 21948
rect 17218 21936 17224 21948
rect 17179 21908 17224 21936
rect 17218 21896 17224 21908
rect 17276 21896 17282 21948
rect 22557 21939 22615 21945
rect 22557 21905 22569 21939
rect 22603 21936 22615 21939
rect 24210 21936 24216 21948
rect 22603 21908 24216 21936
rect 22603 21905 22615 21908
rect 22557 21899 22615 21905
rect 24210 21896 24216 21908
rect 24268 21896 24274 21948
rect 19978 21828 19984 21880
rect 20036 21868 20042 21880
rect 20438 21868 20444 21880
rect 20036 21840 20444 21868
rect 20036 21828 20042 21840
rect 20438 21828 20444 21840
rect 20496 21877 20502 21880
rect 20496 21871 20560 21877
rect 20496 21837 20514 21871
rect 20548 21837 20560 21871
rect 23934 21868 23940 21880
rect 23895 21840 23940 21868
rect 20496 21831 20560 21837
rect 20496 21828 20502 21831
rect 23934 21828 23940 21840
rect 23992 21828 23998 21880
rect 10919 21772 11468 21800
rect 10919 21769 10931 21772
rect 10873 21763 10931 21769
rect 13814 21760 13820 21812
rect 13872 21800 13878 21812
rect 14737 21803 14795 21809
rect 14737 21800 14749 21803
rect 13872 21772 14749 21800
rect 13872 21760 13878 21772
rect 14737 21769 14749 21772
rect 14783 21769 14795 21803
rect 14737 21763 14795 21769
rect 16577 21803 16635 21809
rect 16577 21769 16589 21803
rect 16623 21800 16635 21803
rect 17034 21800 17040 21812
rect 16623 21772 17040 21800
rect 16623 21769 16635 21772
rect 16577 21763 16635 21769
rect 17034 21760 17040 21772
rect 17092 21760 17098 21812
rect 18049 21803 18107 21809
rect 18049 21769 18061 21803
rect 18095 21769 18107 21803
rect 18322 21800 18328 21812
rect 18283 21772 18328 21800
rect 18049 21763 18107 21769
rect 474 21692 480 21744
rect 532 21692 538 21744
rect 14826 21692 14832 21744
rect 14884 21732 14890 21744
rect 14884 21704 14929 21732
rect 14884 21692 14890 21704
rect 16022 21692 16028 21744
rect 16080 21732 16086 21744
rect 16669 21735 16727 21741
rect 16669 21732 16681 21735
rect 16080 21704 16681 21732
rect 16080 21692 16086 21704
rect 16669 21701 16681 21704
rect 16715 21701 16727 21735
rect 16850 21732 16856 21744
rect 16811 21704 16856 21732
rect 16669 21695 16727 21701
rect 16850 21692 16856 21704
rect 16908 21692 16914 21744
rect 14274 21664 14280 21676
rect 14235 21636 14280 21664
rect 14274 21624 14280 21636
rect 14332 21624 14338 21676
rect 16209 21667 16267 21673
rect 16209 21633 16221 21667
rect 16255 21664 16267 21667
rect 18064 21664 18092 21763
rect 18322 21760 18328 21772
rect 18380 21760 18386 21812
rect 24118 21760 24124 21812
rect 24176 21800 24182 21812
rect 24581 21803 24639 21809
rect 24581 21800 24593 21803
rect 24176 21772 24593 21800
rect 24176 21760 24182 21772
rect 24581 21769 24593 21772
rect 24627 21769 24639 21803
rect 24581 21763 24639 21769
rect 20162 21692 20168 21744
rect 20220 21732 20226 21744
rect 20257 21735 20315 21741
rect 20257 21732 20269 21735
rect 20220 21704 20269 21732
rect 20220 21692 20226 21704
rect 20257 21701 20269 21704
rect 20303 21701 20315 21735
rect 20257 21695 20315 21701
rect 18785 21667 18843 21673
rect 18785 21664 18797 21667
rect 16255 21636 18797 21664
rect 16255 21633 16267 21636
rect 16209 21627 16267 21633
rect 18785 21633 18797 21636
rect 18831 21633 18843 21667
rect 18785 21627 18843 21633
rect 11793 21599 11851 21605
rect 11793 21565 11805 21599
rect 11839 21596 11851 21599
rect 12618 21596 12624 21608
rect 11839 21568 12624 21596
rect 11839 21565 11851 21568
rect 11793 21559 11851 21565
rect 12618 21556 12624 21568
rect 12676 21556 12682 21608
rect 15746 21596 15752 21608
rect 15707 21568 15752 21596
rect 15746 21556 15752 21568
rect 15804 21556 15810 21608
rect 16117 21599 16175 21605
rect 16117 21565 16129 21599
rect 16163 21596 16175 21599
rect 16390 21596 16396 21608
rect 16163 21568 16396 21596
rect 16163 21565 16175 21568
rect 16117 21559 16175 21565
rect 16390 21556 16396 21568
rect 16448 21556 16454 21608
rect 16482 21556 16488 21608
rect 16540 21596 16546 21608
rect 16850 21596 16856 21608
rect 16540 21568 16856 21596
rect 16540 21556 16546 21568
rect 16850 21556 16856 21568
rect 16908 21556 16914 21608
rect 21542 21556 21548 21608
rect 21600 21596 21606 21608
rect 21637 21599 21695 21605
rect 21637 21596 21649 21599
rect 21600 21568 21649 21596
rect 21600 21556 21606 21568
rect 21637 21565 21649 21568
rect 21683 21565 21695 21599
rect 21637 21559 21695 21565
rect 23109 21599 23167 21605
rect 23109 21565 23121 21599
rect 23155 21596 23167 21599
rect 23382 21596 23388 21608
rect 23155 21568 23388 21596
rect 23155 21565 23167 21568
rect 23109 21559 23167 21565
rect 23382 21556 23388 21568
rect 23440 21556 23446 21608
rect 24762 21596 24768 21608
rect 24723 21568 24768 21596
rect 24762 21556 24768 21568
rect 24820 21556 24826 21608
rect 1104 21506 26864 21528
rect 1104 21454 5648 21506
rect 5700 21454 5712 21506
rect 5764 21454 5776 21506
rect 5828 21454 5840 21506
rect 5892 21454 14982 21506
rect 15034 21454 15046 21506
rect 15098 21454 15110 21506
rect 15162 21454 15174 21506
rect 15226 21454 24315 21506
rect 24367 21454 24379 21506
rect 24431 21454 24443 21506
rect 24495 21454 24507 21506
rect 24559 21454 26864 21506
rect 1104 21432 26864 21454
rect 11514 21392 11520 21404
rect 11475 21364 11520 21392
rect 11514 21352 11520 21364
rect 11572 21392 11578 21404
rect 14366 21392 14372 21404
rect 11572 21364 12204 21392
rect 14327 21364 14372 21392
rect 11572 21352 11578 21364
rect 12176 21265 12204 21364
rect 14366 21352 14372 21364
rect 14424 21352 14430 21404
rect 14737 21395 14795 21401
rect 14737 21361 14749 21395
rect 14783 21392 14795 21395
rect 14826 21392 14832 21404
rect 14783 21364 14832 21392
rect 14783 21361 14795 21364
rect 14737 21355 14795 21361
rect 14826 21352 14832 21364
rect 14884 21352 14890 21404
rect 15562 21392 15568 21404
rect 15523 21364 15568 21392
rect 15562 21352 15568 21364
rect 15620 21352 15626 21404
rect 16022 21392 16028 21404
rect 15983 21364 16028 21392
rect 16022 21352 16028 21364
rect 16080 21352 16086 21404
rect 19978 21392 19984 21404
rect 19939 21364 19984 21392
rect 19978 21352 19984 21364
rect 20036 21352 20042 21404
rect 22922 21392 22928 21404
rect 22883 21364 22928 21392
rect 22922 21352 22928 21364
rect 22980 21352 22986 21404
rect 24118 21352 24124 21404
rect 24176 21392 24182 21404
rect 24581 21395 24639 21401
rect 24581 21392 24593 21395
rect 24176 21364 24593 21392
rect 24176 21352 24182 21364
rect 24581 21361 24593 21364
rect 24627 21361 24639 21395
rect 24581 21355 24639 21361
rect 15105 21327 15163 21333
rect 15105 21293 15117 21327
rect 15151 21324 15163 21327
rect 16040 21324 16068 21352
rect 22281 21327 22339 21333
rect 22281 21324 22293 21327
rect 15151 21296 16068 21324
rect 22020 21296 22293 21324
rect 15151 21293 15163 21296
rect 15105 21287 15163 21293
rect 12161 21259 12219 21265
rect 12161 21225 12173 21259
rect 12207 21225 12219 21259
rect 12161 21219 12219 21225
rect 12345 21259 12403 21265
rect 12345 21225 12357 21259
rect 12391 21256 12403 21259
rect 12618 21256 12624 21268
rect 12391 21228 12624 21256
rect 12391 21225 12403 21228
rect 12345 21219 12403 21225
rect 12618 21216 12624 21228
rect 12676 21216 12682 21268
rect 16482 21216 16488 21268
rect 16540 21256 16546 21268
rect 16577 21259 16635 21265
rect 16577 21256 16589 21259
rect 16540 21228 16589 21256
rect 16540 21216 16546 21228
rect 16577 21225 16589 21228
rect 16623 21225 16635 21259
rect 16577 21219 16635 21225
rect 17586 21216 17592 21268
rect 17644 21256 17650 21268
rect 18693 21259 18751 21265
rect 18693 21256 18705 21259
rect 17644 21228 18705 21256
rect 17644 21216 17650 21228
rect 18693 21225 18705 21228
rect 18739 21256 18751 21259
rect 19242 21256 19248 21268
rect 18739 21228 19248 21256
rect 18739 21225 18751 21228
rect 18693 21219 18751 21225
rect 19242 21216 19248 21228
rect 19300 21216 19306 21268
rect 20530 21216 20536 21268
rect 20588 21256 20594 21268
rect 21453 21259 21511 21265
rect 21453 21256 21465 21259
rect 20588 21228 21465 21256
rect 20588 21216 20594 21228
rect 21453 21225 21465 21228
rect 21499 21256 21511 21259
rect 21542 21256 21548 21268
rect 21499 21228 21548 21256
rect 21499 21225 21511 21228
rect 21453 21219 21511 21225
rect 21542 21216 21548 21228
rect 21600 21256 21606 21268
rect 21913 21259 21971 21265
rect 21913 21256 21925 21259
rect 21600 21228 21925 21256
rect 21600 21216 21606 21228
rect 21913 21225 21925 21228
rect 21959 21225 21971 21259
rect 21913 21219 21971 21225
rect 13265 21191 13323 21197
rect 13265 21188 13277 21191
rect 13096 21160 13277 21188
rect 11698 21052 11704 21064
rect 11659 21024 11704 21052
rect 11698 21012 11704 21024
rect 11756 21012 11762 21064
rect 11790 21012 11796 21064
rect 11848 21052 11854 21064
rect 12069 21055 12127 21061
rect 12069 21052 12081 21055
rect 11848 21024 12081 21052
rect 11848 21012 11854 21024
rect 12069 21021 12081 21024
rect 12115 21021 12127 21055
rect 12069 21015 12127 21021
rect 12434 21012 12440 21064
rect 12492 21052 12498 21064
rect 13096 21061 13124 21160
rect 13265 21157 13277 21160
rect 13311 21157 13323 21191
rect 13265 21151 13323 21157
rect 20898 21148 20904 21200
rect 20956 21188 20962 21200
rect 21361 21191 21419 21197
rect 21361 21188 21373 21191
rect 20956 21160 21373 21188
rect 20956 21148 20962 21160
rect 21361 21157 21373 21160
rect 21407 21188 21419 21191
rect 22020 21188 22048 21296
rect 22281 21293 22293 21296
rect 22327 21293 22339 21327
rect 22281 21287 22339 21293
rect 23385 21259 23443 21265
rect 23385 21256 23397 21259
rect 22756 21228 23397 21256
rect 22756 21197 22784 21228
rect 23385 21225 23397 21228
rect 23431 21256 23443 21259
rect 24029 21259 24087 21265
rect 24029 21256 24041 21259
rect 23431 21228 24041 21256
rect 23431 21225 23443 21228
rect 23385 21219 23443 21225
rect 24029 21225 24041 21228
rect 24075 21225 24087 21259
rect 24029 21219 24087 21225
rect 21407 21160 22048 21188
rect 22741 21191 22799 21197
rect 21407 21157 21419 21160
rect 21361 21151 21419 21157
rect 22741 21157 22753 21191
rect 22787 21157 22799 21191
rect 23845 21191 23903 21197
rect 23845 21188 23857 21191
rect 22741 21151 22799 21157
rect 23676 21160 23857 21188
rect 13538 21120 13544 21132
rect 13499 21092 13544 21120
rect 13538 21080 13544 21092
rect 13596 21080 13602 21132
rect 16485 21123 16543 21129
rect 16485 21120 16497 21123
rect 15856 21092 16497 21120
rect 15856 21064 15884 21092
rect 16485 21089 16497 21092
rect 16531 21089 16543 21123
rect 18509 21123 18567 21129
rect 18509 21120 18521 21123
rect 16485 21083 16543 21089
rect 18064 21092 18521 21120
rect 18064 21064 18092 21092
rect 18509 21089 18521 21092
rect 18555 21089 18567 21123
rect 18509 21083 18567 21089
rect 20717 21123 20775 21129
rect 20717 21089 20729 21123
rect 20763 21120 20775 21123
rect 20990 21120 20996 21132
rect 20763 21092 20996 21120
rect 20763 21089 20775 21092
rect 20717 21083 20775 21089
rect 20990 21080 20996 21092
rect 21048 21120 21054 21132
rect 21269 21123 21327 21129
rect 21269 21120 21281 21123
rect 21048 21092 21281 21120
rect 21048 21080 21054 21092
rect 21269 21089 21281 21092
rect 21315 21089 21327 21123
rect 21269 21083 21327 21089
rect 23676 21064 23704 21160
rect 23845 21157 23857 21160
rect 23891 21157 23903 21191
rect 25130 21188 25136 21200
rect 25091 21160 25136 21188
rect 23845 21151 23903 21157
rect 25130 21148 25136 21160
rect 25188 21188 25194 21200
rect 25685 21191 25743 21197
rect 25685 21188 25697 21191
rect 25188 21160 25697 21188
rect 25188 21148 25194 21160
rect 25685 21157 25697 21160
rect 25731 21157 25743 21191
rect 25685 21151 25743 21157
rect 26234 21080 26240 21132
rect 26292 21120 26298 21132
rect 27522 21120 27528 21132
rect 26292 21092 27528 21120
rect 26292 21080 26298 21092
rect 27522 21080 27528 21092
rect 27580 21080 27586 21132
rect 13081 21055 13139 21061
rect 13081 21052 13093 21055
rect 12492 21024 13093 21052
rect 12492 21012 12498 21024
rect 13081 21021 13093 21024
rect 13127 21021 13139 21055
rect 15838 21052 15844 21064
rect 15799 21024 15844 21052
rect 13081 21015 13139 21021
rect 15838 21012 15844 21024
rect 15896 21012 15902 21064
rect 16390 21052 16396 21064
rect 16351 21024 16396 21052
rect 16390 21012 16396 21024
rect 16448 21012 16454 21064
rect 17034 21052 17040 21064
rect 16995 21024 17040 21052
rect 17034 21012 17040 21024
rect 17092 21012 17098 21064
rect 17586 21052 17592 21064
rect 17547 21024 17592 21052
rect 17586 21012 17592 21024
rect 17644 21012 17650 21064
rect 18046 21052 18052 21064
rect 18007 21024 18052 21052
rect 18046 21012 18052 21024
rect 18104 21012 18110 21064
rect 18138 21012 18144 21064
rect 18196 21052 18202 21064
rect 18196 21024 18241 21052
rect 18196 21012 18202 21024
rect 18598 21012 18604 21064
rect 18656 21052 18662 21064
rect 19153 21055 19211 21061
rect 19153 21052 19165 21055
rect 18656 21024 19165 21052
rect 18656 21012 18662 21024
rect 19153 21021 19165 21024
rect 19199 21021 19211 21055
rect 19153 21015 19211 21021
rect 20162 21012 20168 21064
rect 20220 21052 20226 21064
rect 20257 21055 20315 21061
rect 20257 21052 20269 21055
rect 20220 21024 20269 21052
rect 20220 21012 20226 21024
rect 20257 21021 20269 21024
rect 20303 21021 20315 21055
rect 20898 21052 20904 21064
rect 20859 21024 20904 21052
rect 20257 21015 20315 21021
rect 20898 21012 20904 21024
rect 20956 21012 20962 21064
rect 23658 21052 23664 21064
rect 23619 21024 23664 21052
rect 23658 21012 23664 21024
rect 23716 21012 23722 21064
rect 25314 21052 25320 21064
rect 25275 21024 25320 21052
rect 25314 21012 25320 21024
rect 25372 21012 25378 21064
rect 1104 20962 26864 20984
rect 1104 20910 10315 20962
rect 10367 20910 10379 20962
rect 10431 20910 10443 20962
rect 10495 20910 10507 20962
rect 10559 20910 19648 20962
rect 19700 20910 19712 20962
rect 19764 20910 19776 20962
rect 19828 20910 19840 20962
rect 19892 20910 26864 20962
rect 1104 20888 26864 20910
rect 13814 20808 13820 20860
rect 13872 20848 13878 20860
rect 14277 20851 14335 20857
rect 14277 20848 14289 20851
rect 13872 20820 14289 20848
rect 13872 20808 13878 20820
rect 14277 20817 14289 20820
rect 14323 20817 14335 20851
rect 14642 20848 14648 20860
rect 14603 20820 14648 20848
rect 14277 20811 14335 20817
rect 14642 20808 14648 20820
rect 14700 20808 14706 20860
rect 16850 20808 16856 20860
rect 16908 20848 16914 20860
rect 17037 20851 17095 20857
rect 17037 20848 17049 20851
rect 16908 20820 17049 20848
rect 16908 20808 16914 20820
rect 17037 20817 17049 20820
rect 17083 20817 17095 20851
rect 17037 20811 17095 20817
rect 18049 20851 18107 20857
rect 18049 20817 18061 20851
rect 18095 20848 18107 20851
rect 18598 20848 18604 20860
rect 18095 20820 18604 20848
rect 18095 20817 18107 20820
rect 18049 20811 18107 20817
rect 18598 20808 18604 20820
rect 18656 20808 18662 20860
rect 22186 20808 22192 20860
rect 22244 20848 22250 20860
rect 24670 20848 24676 20860
rect 22244 20820 24676 20848
rect 22244 20808 22250 20820
rect 24670 20808 24676 20820
rect 24728 20808 24734 20860
rect 12618 20740 12624 20792
rect 12676 20789 12682 20792
rect 12676 20783 12740 20789
rect 12676 20749 12694 20783
rect 12728 20749 12740 20783
rect 18414 20780 18420 20792
rect 18375 20752 18420 20780
rect 12676 20743 12740 20749
rect 12676 20740 12682 20743
rect 18414 20740 18420 20752
rect 18472 20740 18478 20792
rect 20432 20783 20490 20789
rect 20432 20749 20444 20783
rect 20478 20780 20490 20783
rect 20530 20780 20536 20792
rect 20478 20752 20536 20780
rect 20478 20749 20490 20752
rect 20432 20743 20490 20749
rect 20530 20740 20536 20752
rect 20588 20740 20594 20792
rect 24854 20740 24860 20792
rect 24912 20740 24918 20792
rect 15286 20672 15292 20724
rect 15344 20712 15350 20724
rect 15746 20712 15752 20724
rect 15344 20684 15752 20712
rect 15344 20672 15350 20684
rect 15746 20672 15752 20684
rect 15804 20712 15810 20724
rect 15913 20715 15971 20721
rect 15913 20712 15925 20715
rect 15804 20684 15925 20712
rect 15804 20672 15810 20684
rect 15913 20681 15925 20684
rect 15959 20712 15971 20715
rect 16482 20712 16488 20724
rect 15959 20684 16488 20712
rect 15959 20681 15971 20684
rect 15913 20675 15971 20681
rect 16482 20672 16488 20684
rect 16540 20672 16546 20724
rect 23842 20712 23848 20724
rect 23803 20684 23848 20712
rect 23842 20672 23848 20684
rect 23900 20672 23906 20724
rect 24872 20712 24900 20740
rect 25133 20715 25191 20721
rect 25133 20712 25145 20715
rect 24872 20684 25145 20712
rect 25133 20681 25145 20684
rect 25179 20712 25191 20715
rect 25314 20712 25320 20724
rect 25179 20684 25320 20712
rect 25179 20681 25191 20684
rect 25133 20675 25191 20681
rect 25314 20672 25320 20684
rect 25372 20672 25378 20724
rect 12434 20604 12440 20656
rect 12492 20644 12498 20656
rect 12492 20616 12537 20644
rect 12492 20604 12498 20616
rect 15378 20604 15384 20656
rect 15436 20644 15442 20656
rect 15654 20644 15660 20656
rect 15436 20616 15660 20644
rect 15436 20604 15442 20616
rect 15654 20604 15660 20616
rect 15712 20604 15718 20656
rect 17954 20604 17960 20656
rect 18012 20644 18018 20656
rect 18509 20647 18567 20653
rect 18509 20644 18521 20647
rect 18012 20616 18521 20644
rect 18012 20604 18018 20616
rect 18509 20613 18521 20616
rect 18555 20613 18567 20647
rect 18509 20607 18567 20613
rect 18693 20647 18751 20653
rect 18693 20613 18705 20647
rect 18739 20644 18751 20647
rect 19058 20644 19064 20656
rect 18739 20616 19064 20644
rect 18739 20613 18751 20616
rect 18693 20607 18751 20613
rect 19058 20604 19064 20616
rect 19116 20604 19122 20656
rect 20162 20644 20168 20656
rect 20123 20616 20168 20644
rect 20162 20604 20168 20616
rect 20220 20604 20226 20656
rect 24121 20647 24179 20653
rect 24121 20613 24133 20647
rect 24167 20644 24179 20647
rect 24854 20644 24860 20656
rect 24167 20616 24860 20644
rect 24167 20613 24179 20616
rect 24121 20607 24179 20613
rect 24854 20604 24860 20616
rect 24912 20604 24918 20656
rect 25409 20647 25467 20653
rect 25409 20613 25421 20647
rect 25455 20644 25467 20647
rect 25498 20644 25504 20656
rect 25455 20616 25504 20644
rect 25455 20613 25467 20616
rect 25409 20607 25467 20613
rect 25498 20604 25504 20616
rect 25556 20604 25562 20656
rect 11790 20508 11796 20520
rect 11751 20480 11796 20508
rect 11790 20468 11796 20480
rect 11848 20468 11854 20520
rect 13814 20508 13820 20520
rect 13775 20480 13820 20508
rect 13814 20468 13820 20480
rect 13872 20468 13878 20520
rect 15378 20508 15384 20520
rect 15339 20480 15384 20508
rect 15378 20468 15384 20480
rect 15436 20468 15442 20520
rect 20806 20468 20812 20520
rect 20864 20508 20870 20520
rect 21545 20511 21603 20517
rect 21545 20508 21557 20511
rect 20864 20480 21557 20508
rect 20864 20468 20870 20480
rect 21545 20477 21557 20480
rect 21591 20477 21603 20511
rect 22830 20508 22836 20520
rect 22791 20480 22836 20508
rect 21545 20471 21603 20477
rect 22830 20468 22836 20480
rect 22888 20468 22894 20520
rect 1104 20418 26864 20440
rect 1104 20366 5648 20418
rect 5700 20366 5712 20418
rect 5764 20366 5776 20418
rect 5828 20366 5840 20418
rect 5892 20366 14982 20418
rect 15034 20366 15046 20418
rect 15098 20366 15110 20418
rect 15162 20366 15174 20418
rect 15226 20366 24315 20418
rect 24367 20366 24379 20418
rect 24431 20366 24443 20418
rect 24495 20366 24507 20418
rect 24559 20366 26864 20418
rect 1104 20344 26864 20366
rect 12434 20264 12440 20316
rect 12492 20304 12498 20316
rect 12529 20307 12587 20313
rect 12529 20304 12541 20307
rect 12492 20276 12541 20304
rect 12492 20264 12498 20276
rect 12529 20273 12541 20276
rect 12575 20273 12587 20307
rect 12529 20267 12587 20273
rect 14737 20307 14795 20313
rect 14737 20273 14749 20307
rect 14783 20304 14795 20307
rect 15286 20304 15292 20316
rect 14783 20276 15292 20304
rect 14783 20273 14795 20276
rect 14737 20267 14795 20273
rect 15286 20264 15292 20276
rect 15344 20264 15350 20316
rect 16482 20264 16488 20316
rect 16540 20304 16546 20316
rect 16669 20307 16727 20313
rect 16669 20304 16681 20307
rect 16540 20276 16681 20304
rect 16540 20264 16546 20276
rect 16669 20273 16681 20276
rect 16715 20273 16727 20307
rect 17954 20304 17960 20316
rect 17915 20276 17960 20304
rect 16669 20267 16727 20273
rect 17954 20264 17960 20276
rect 18012 20264 18018 20316
rect 19334 20264 19340 20316
rect 19392 20304 19398 20316
rect 19429 20307 19487 20313
rect 19429 20304 19441 20307
rect 19392 20276 19441 20304
rect 19392 20264 19398 20276
rect 19429 20273 19441 20276
rect 19475 20273 19487 20307
rect 20530 20304 20536 20316
rect 20491 20276 20536 20304
rect 19429 20267 19487 20273
rect 20530 20264 20536 20276
rect 20588 20264 20594 20316
rect 23474 20264 23480 20316
rect 23532 20304 23538 20316
rect 23532 20276 23704 20304
rect 23532 20264 23538 20276
rect 19058 20196 19064 20248
rect 19116 20236 19122 20248
rect 19797 20239 19855 20245
rect 19797 20236 19809 20239
rect 19116 20208 19809 20236
rect 19116 20196 19122 20208
rect 19797 20205 19809 20208
rect 19843 20236 19855 20239
rect 20806 20236 20812 20248
rect 19843 20208 20812 20236
rect 19843 20205 19855 20208
rect 19797 20199 19855 20205
rect 20806 20196 20812 20208
rect 20864 20196 20870 20248
rect 23676 20236 23704 20276
rect 23842 20264 23848 20316
rect 23900 20304 23906 20316
rect 24397 20307 24455 20313
rect 24397 20304 24409 20307
rect 23900 20276 24409 20304
rect 23900 20264 23906 20276
rect 24397 20273 24409 20276
rect 24443 20273 24455 20307
rect 25130 20304 25136 20316
rect 25091 20276 25136 20304
rect 24397 20267 24455 20273
rect 25130 20264 25136 20276
rect 25188 20264 25194 20316
rect 25314 20264 25320 20316
rect 25372 20304 25378 20316
rect 25501 20307 25559 20313
rect 25501 20304 25513 20307
rect 25372 20276 25513 20304
rect 25372 20264 25378 20276
rect 25501 20273 25513 20276
rect 25547 20273 25559 20307
rect 25501 20267 25559 20273
rect 24121 20239 24179 20245
rect 24121 20236 24133 20239
rect 23676 20208 24133 20236
rect 24121 20205 24133 20208
rect 24167 20205 24179 20239
rect 24121 20199 24179 20205
rect 17221 20171 17279 20177
rect 17221 20137 17233 20171
rect 17267 20168 17279 20171
rect 17267 20140 18184 20168
rect 17267 20137 17279 20140
rect 17221 20131 17279 20137
rect 10413 20103 10471 20109
rect 10413 20069 10425 20103
rect 10459 20100 10471 20103
rect 10505 20103 10563 20109
rect 10505 20100 10517 20103
rect 10459 20072 10517 20100
rect 10459 20069 10471 20072
rect 10413 20063 10471 20069
rect 10505 20069 10517 20072
rect 10551 20100 10563 20103
rect 12161 20103 12219 20109
rect 12161 20100 12173 20103
rect 10551 20072 12173 20100
rect 10551 20069 10563 20072
rect 10505 20063 10563 20069
rect 12161 20069 12173 20072
rect 12207 20100 12219 20103
rect 12434 20100 12440 20112
rect 12207 20072 12440 20100
rect 12207 20069 12219 20072
rect 12161 20063 12219 20069
rect 12434 20060 12440 20072
rect 12492 20100 12498 20112
rect 12710 20100 12716 20112
rect 12492 20072 12716 20100
rect 12492 20060 12498 20072
rect 12710 20060 12716 20072
rect 12768 20060 12774 20112
rect 12986 20109 12992 20112
rect 12980 20100 12992 20109
rect 12899 20072 12992 20100
rect 12980 20063 12992 20072
rect 13044 20100 13050 20112
rect 13722 20100 13728 20112
rect 13044 20072 13728 20100
rect 12986 20060 12992 20063
rect 13044 20060 13050 20072
rect 13722 20060 13728 20072
rect 13780 20060 13786 20112
rect 15289 20103 15347 20109
rect 15289 20100 15301 20103
rect 15028 20072 15301 20100
rect 10772 20035 10830 20041
rect 10772 20001 10784 20035
rect 10818 20032 10830 20035
rect 10870 20032 10876 20044
rect 10818 20004 10876 20032
rect 10818 20001 10830 20004
rect 10772 19995 10830 20001
rect 10870 19992 10876 20004
rect 10928 19992 10934 20044
rect 12618 20032 12624 20044
rect 11900 20004 12624 20032
rect 11900 19973 11928 20004
rect 12618 19992 12624 20004
rect 12676 20032 12682 20044
rect 13262 20032 13268 20044
rect 12676 20004 13268 20032
rect 12676 19992 12682 20004
rect 13262 19992 13268 20004
rect 13320 19992 13326 20044
rect 15028 19976 15056 20072
rect 15289 20069 15301 20072
rect 15335 20069 15347 20103
rect 15289 20063 15347 20069
rect 15378 20060 15384 20112
rect 15436 20100 15442 20112
rect 15545 20103 15603 20109
rect 15545 20100 15557 20103
rect 15436 20072 15557 20100
rect 15436 20060 15442 20072
rect 15545 20069 15557 20072
rect 15591 20069 15603 20103
rect 18049 20103 18107 20109
rect 18049 20100 18061 20103
rect 15545 20063 15603 20069
rect 17512 20072 18061 20100
rect 11885 19967 11943 19973
rect 11885 19933 11897 19967
rect 11931 19933 11943 19967
rect 14090 19964 14096 19976
rect 14051 19936 14096 19964
rect 11885 19927 11943 19933
rect 14090 19924 14096 19936
rect 14148 19924 14154 19976
rect 15010 19964 15016 19976
rect 14971 19936 15016 19964
rect 15010 19924 15016 19936
rect 15068 19924 15074 19976
rect 15654 19924 15660 19976
rect 15712 19964 15718 19976
rect 17512 19973 17540 20072
rect 18049 20069 18061 20072
rect 18095 20069 18107 20103
rect 18156 20100 18184 20140
rect 18316 20103 18374 20109
rect 18316 20100 18328 20103
rect 18156 20072 18328 20100
rect 18049 20063 18107 20069
rect 18316 20069 18328 20072
rect 18362 20100 18374 20103
rect 19076 20100 19104 20196
rect 20901 20171 20959 20177
rect 20901 20137 20913 20171
rect 20947 20168 20959 20171
rect 20990 20168 20996 20180
rect 20947 20140 20996 20168
rect 20947 20137 20959 20140
rect 20901 20131 20959 20137
rect 20990 20128 20996 20140
rect 21048 20128 21054 20180
rect 18362 20072 19104 20100
rect 22097 20103 22155 20109
rect 18362 20069 18374 20072
rect 18316 20063 18374 20069
rect 22097 20069 22109 20103
rect 22143 20100 22155 20103
rect 22554 20100 22560 20112
rect 22143 20072 22560 20100
rect 22143 20069 22155 20072
rect 22097 20063 22155 20069
rect 18064 20032 18092 20063
rect 22554 20060 22560 20072
rect 22612 20060 22618 20112
rect 22741 20103 22799 20109
rect 22741 20100 22753 20103
rect 22664 20072 22753 20100
rect 19242 20032 19248 20044
rect 18064 20004 19248 20032
rect 19242 19992 19248 20004
rect 19300 20032 19306 20044
rect 20162 20032 20168 20044
rect 19300 20004 20168 20032
rect 19300 19992 19306 20004
rect 20162 19992 20168 20004
rect 20220 19992 20226 20044
rect 22664 19976 22692 20072
rect 22741 20069 22753 20072
rect 22787 20069 22799 20103
rect 22741 20063 22799 20069
rect 22830 20060 22836 20112
rect 22888 20100 22894 20112
rect 22997 20103 23055 20109
rect 22997 20100 23009 20103
rect 22888 20072 23009 20100
rect 22888 20060 22894 20072
rect 22997 20069 23009 20072
rect 23043 20069 23055 20103
rect 22997 20063 23055 20069
rect 23474 20060 23480 20112
rect 23532 20100 23538 20112
rect 23934 20100 23940 20112
rect 23532 20072 23940 20100
rect 23532 20060 23538 20072
rect 23934 20060 23940 20072
rect 23992 20060 23998 20112
rect 24949 20103 25007 20109
rect 24949 20069 24961 20103
rect 24995 20069 25007 20103
rect 24949 20063 25007 20069
rect 24964 19976 24992 20063
rect 17497 19967 17555 19973
rect 17497 19964 17509 19967
rect 15712 19936 17509 19964
rect 15712 19924 15718 19936
rect 17497 19933 17509 19936
rect 17543 19933 17555 19967
rect 22646 19964 22652 19976
rect 22607 19936 22652 19964
rect 17497 19927 17555 19933
rect 22646 19924 22652 19936
rect 22704 19924 22710 19976
rect 24857 19967 24915 19973
rect 24857 19933 24869 19967
rect 24903 19964 24915 19967
rect 24946 19964 24952 19976
rect 24903 19936 24952 19964
rect 24903 19933 24915 19936
rect 24857 19927 24915 19933
rect 24946 19924 24952 19936
rect 25004 19924 25010 19976
rect 1104 19874 26864 19896
rect 1104 19822 10315 19874
rect 10367 19822 10379 19874
rect 10431 19822 10443 19874
rect 10495 19822 10507 19874
rect 10559 19822 19648 19874
rect 19700 19822 19712 19874
rect 19764 19822 19776 19874
rect 19828 19822 19840 19874
rect 19892 19822 26864 19874
rect 1104 19800 26864 19822
rect 10597 19763 10655 19769
rect 10597 19729 10609 19763
rect 10643 19760 10655 19763
rect 10870 19760 10876 19772
rect 10643 19732 10876 19760
rect 10643 19729 10655 19732
rect 10597 19723 10655 19729
rect 10870 19720 10876 19732
rect 10928 19720 10934 19772
rect 11698 19720 11704 19772
rect 11756 19760 11762 19772
rect 12069 19763 12127 19769
rect 12069 19760 12081 19763
rect 11756 19732 12081 19760
rect 11756 19720 11762 19732
rect 12069 19729 12081 19732
rect 12115 19729 12127 19763
rect 12986 19760 12992 19772
rect 12947 19732 12992 19760
rect 12069 19723 12127 19729
rect 12986 19720 12992 19732
rect 13044 19720 13050 19772
rect 13262 19760 13268 19772
rect 13223 19732 13268 19760
rect 13262 19720 13268 19732
rect 13320 19720 13326 19772
rect 15289 19763 15347 19769
rect 15289 19729 15301 19763
rect 15335 19760 15347 19763
rect 15378 19760 15384 19772
rect 15335 19732 15384 19760
rect 15335 19729 15347 19732
rect 15289 19723 15347 19729
rect 15378 19720 15384 19732
rect 15436 19720 15442 19772
rect 17954 19720 17960 19772
rect 18012 19760 18018 19772
rect 18325 19763 18383 19769
rect 18325 19760 18337 19763
rect 18012 19732 18337 19760
rect 18012 19720 18018 19732
rect 18325 19729 18337 19732
rect 18371 19760 18383 19763
rect 18414 19760 18420 19772
rect 18371 19732 18420 19760
rect 18371 19729 18383 19732
rect 18325 19723 18383 19729
rect 18414 19720 18420 19732
rect 18472 19720 18478 19772
rect 22005 19763 22063 19769
rect 22005 19729 22017 19763
rect 22051 19760 22063 19763
rect 24121 19763 24179 19769
rect 24121 19760 24133 19763
rect 22051 19732 24133 19760
rect 22051 19729 22063 19732
rect 22005 19723 22063 19729
rect 24121 19729 24133 19732
rect 24167 19760 24179 19763
rect 24762 19760 24768 19772
rect 24167 19732 24768 19760
rect 24167 19729 24179 19732
rect 24121 19723 24179 19729
rect 24762 19720 24768 19732
rect 24820 19720 24826 19772
rect 25406 19760 25412 19772
rect 25367 19732 25412 19760
rect 25406 19720 25412 19732
rect 25464 19720 25470 19772
rect 13725 19695 13783 19701
rect 13725 19661 13737 19695
rect 13771 19692 13783 19695
rect 14090 19692 14096 19704
rect 13771 19664 14096 19692
rect 13771 19661 13783 19664
rect 13725 19655 13783 19661
rect 14090 19652 14096 19664
rect 14148 19701 14154 19704
rect 14148 19695 14212 19701
rect 14148 19661 14166 19695
rect 14200 19661 14212 19695
rect 14148 19655 14212 19661
rect 14148 19652 14154 19655
rect 15654 19652 15660 19704
rect 15712 19652 15718 19704
rect 12710 19584 12716 19636
rect 12768 19624 12774 19636
rect 13909 19627 13967 19633
rect 13909 19624 13921 19627
rect 12768 19596 13921 19624
rect 12768 19584 12774 19596
rect 13909 19593 13921 19596
rect 13955 19624 13967 19627
rect 14734 19624 14740 19636
rect 13955 19596 14740 19624
rect 13955 19593 13967 19596
rect 13909 19587 13967 19593
rect 14734 19584 14740 19596
rect 14792 19624 14798 19636
rect 15010 19624 15016 19636
rect 14792 19596 15016 19624
rect 14792 19584 14798 19596
rect 15010 19584 15016 19596
rect 15068 19624 15074 19636
rect 15672 19624 15700 19652
rect 15749 19627 15807 19633
rect 15749 19624 15761 19627
rect 15068 19596 15761 19624
rect 15068 19584 15074 19596
rect 15749 19593 15761 19596
rect 15795 19593 15807 19627
rect 15749 19587 15807 19593
rect 18138 19584 18144 19636
rect 18196 19624 18202 19636
rect 18690 19624 18696 19636
rect 18196 19596 18696 19624
rect 18196 19584 18202 19596
rect 18690 19584 18696 19596
rect 18748 19584 18754 19636
rect 18966 19624 18972 19636
rect 18927 19596 18972 19624
rect 18966 19584 18972 19596
rect 19024 19584 19030 19636
rect 22373 19627 22431 19633
rect 22373 19624 22385 19627
rect 21836 19596 22385 19624
rect 12434 19516 12440 19568
rect 12492 19556 12498 19568
rect 12492 19528 12537 19556
rect 12492 19516 12498 19528
rect 15654 19516 15660 19568
rect 15712 19556 15718 19568
rect 16117 19559 16175 19565
rect 16117 19556 16129 19559
rect 15712 19528 16129 19556
rect 15712 19516 15718 19528
rect 16117 19525 16129 19528
rect 16163 19525 16175 19559
rect 16117 19519 16175 19525
rect 20990 19420 20996 19432
rect 20951 19392 20996 19420
rect 20990 19380 20996 19392
rect 21048 19380 21054 19432
rect 21542 19380 21548 19432
rect 21600 19420 21606 19432
rect 21836 19429 21864 19596
rect 22373 19593 22385 19596
rect 22419 19593 22431 19627
rect 24026 19624 24032 19636
rect 23987 19596 24032 19624
rect 22373 19587 22431 19593
rect 24026 19584 24032 19596
rect 24084 19584 24090 19636
rect 24854 19584 24860 19636
rect 24912 19624 24918 19636
rect 25225 19627 25283 19633
rect 25225 19624 25237 19627
rect 24912 19596 25237 19624
rect 24912 19584 24918 19596
rect 25225 19593 25237 19596
rect 25271 19624 25283 19627
rect 25866 19624 25872 19636
rect 25271 19596 25872 19624
rect 25271 19593 25283 19596
rect 25225 19587 25283 19593
rect 25866 19584 25872 19596
rect 25924 19584 25930 19636
rect 22094 19516 22100 19568
rect 22152 19556 22158 19568
rect 22465 19559 22523 19565
rect 22465 19556 22477 19559
rect 22152 19528 22477 19556
rect 22152 19516 22158 19528
rect 22465 19525 22477 19528
rect 22511 19525 22523 19559
rect 22465 19519 22523 19525
rect 22554 19516 22560 19568
rect 22612 19556 22618 19568
rect 22612 19528 22657 19556
rect 22612 19516 22618 19528
rect 22830 19516 22836 19568
rect 22888 19556 22894 19568
rect 24118 19556 24124 19568
rect 22888 19528 24124 19556
rect 22888 19516 22894 19528
rect 24118 19516 24124 19528
rect 24176 19556 24182 19568
rect 24213 19559 24271 19565
rect 24213 19556 24225 19559
rect 24176 19528 24225 19556
rect 24176 19516 24182 19528
rect 24213 19525 24225 19528
rect 24259 19525 24271 19559
rect 24213 19519 24271 19525
rect 21821 19423 21879 19429
rect 21821 19420 21833 19423
rect 21600 19392 21833 19420
rect 21600 19380 21606 19392
rect 21821 19389 21833 19392
rect 21867 19389 21879 19423
rect 23658 19420 23664 19432
rect 23619 19392 23664 19420
rect 21821 19383 21879 19389
rect 23658 19380 23664 19392
rect 23716 19380 23722 19432
rect 1104 19330 26864 19352
rect 1104 19278 5648 19330
rect 5700 19278 5712 19330
rect 5764 19278 5776 19330
rect 5828 19278 5840 19330
rect 5892 19278 14982 19330
rect 15034 19278 15046 19330
rect 15098 19278 15110 19330
rect 15162 19278 15174 19330
rect 15226 19278 24315 19330
rect 24367 19278 24379 19330
rect 24431 19278 24443 19330
rect 24495 19278 24507 19330
rect 24559 19278 26864 19330
rect 1104 19256 26864 19278
rect 14734 19216 14740 19228
rect 14695 19188 14740 19216
rect 14734 19176 14740 19188
rect 14792 19176 14798 19228
rect 18690 19216 18696 19228
rect 18651 19188 18696 19216
rect 18690 19176 18696 19188
rect 18748 19176 18754 19228
rect 24026 19176 24032 19228
rect 24084 19216 24090 19228
rect 24397 19219 24455 19225
rect 24397 19216 24409 19219
rect 24084 19188 24409 19216
rect 24084 19176 24090 19188
rect 24397 19185 24409 19188
rect 24443 19185 24455 19219
rect 24762 19216 24768 19228
rect 24723 19188 24768 19216
rect 24397 19179 24455 19185
rect 24762 19176 24768 19188
rect 24820 19176 24826 19228
rect 25866 19216 25872 19228
rect 25827 19188 25872 19216
rect 25866 19176 25872 19188
rect 25924 19176 25930 19228
rect 12342 19108 12348 19160
rect 12400 19148 12406 19160
rect 20901 19151 20959 19157
rect 12400 19120 12756 19148
rect 12400 19108 12406 19120
rect 11698 19040 11704 19092
rect 11756 19080 11762 19092
rect 12728 19089 12756 19120
rect 20901 19117 20913 19151
rect 20947 19117 20959 19151
rect 22094 19148 22100 19160
rect 22055 19120 22100 19148
rect 20901 19111 20959 19117
rect 12529 19083 12587 19089
rect 12529 19080 12541 19083
rect 11756 19052 12541 19080
rect 11756 19040 11762 19052
rect 12529 19049 12541 19052
rect 12575 19049 12587 19083
rect 12529 19043 12587 19049
rect 12713 19083 12771 19089
rect 12713 19049 12725 19083
rect 12759 19080 12771 19083
rect 12986 19080 12992 19092
rect 12759 19052 12992 19080
rect 12759 19049 12771 19052
rect 12713 19043 12771 19049
rect 12986 19040 12992 19052
rect 13044 19040 13050 19092
rect 14090 19040 14096 19092
rect 14148 19080 14154 19092
rect 14185 19083 14243 19089
rect 14185 19080 14197 19083
rect 14148 19052 14197 19080
rect 14148 19040 14154 19052
rect 14185 19049 14197 19052
rect 14231 19049 14243 19083
rect 14185 19043 14243 19049
rect 15378 19040 15384 19092
rect 15436 19080 15442 19092
rect 15841 19083 15899 19089
rect 15841 19080 15853 19083
rect 15436 19052 15853 19080
rect 15436 19040 15442 19052
rect 15841 19049 15853 19052
rect 15887 19049 15899 19083
rect 15841 19043 15899 19049
rect 11977 19015 12035 19021
rect 11977 18981 11989 19015
rect 12023 19012 12035 19015
rect 12434 19012 12440 19024
rect 12023 18984 12440 19012
rect 12023 18981 12035 18984
rect 11977 18975 12035 18981
rect 12434 18972 12440 18984
rect 12492 19012 12498 19024
rect 15105 19015 15163 19021
rect 12492 18984 12537 19012
rect 12492 18972 12498 18984
rect 15105 18981 15117 19015
rect 15151 19012 15163 19015
rect 15654 19012 15660 19024
rect 15151 18984 15660 19012
rect 15151 18981 15163 18984
rect 15105 18975 15163 18981
rect 15654 18972 15660 18984
rect 15712 18972 15718 19024
rect 18046 18972 18052 19024
rect 18104 19012 18110 19024
rect 18233 19015 18291 19021
rect 18233 19012 18245 19015
rect 18104 18984 18245 19012
rect 18104 18972 18110 18984
rect 18233 18981 18245 18984
rect 18279 18981 18291 19015
rect 20916 19012 20944 19111
rect 22094 19108 22100 19120
rect 22152 19108 22158 19160
rect 24118 19148 24124 19160
rect 24079 19120 24124 19148
rect 24118 19108 24124 19120
rect 24176 19108 24182 19160
rect 20990 19040 20996 19092
rect 21048 19080 21054 19092
rect 21453 19083 21511 19089
rect 21453 19080 21465 19083
rect 21048 19052 21465 19080
rect 21048 19040 21054 19052
rect 21453 19049 21465 19052
rect 21499 19049 21511 19083
rect 22646 19080 22652 19092
rect 21453 19043 21511 19049
rect 22480 19052 22652 19080
rect 22094 19012 22100 19024
rect 20916 18984 22100 19012
rect 18233 18975 18291 18981
rect 22094 18972 22100 18984
rect 22152 18972 22158 19024
rect 13446 18944 13452 18956
rect 13407 18916 13452 18944
rect 13446 18904 13452 18916
rect 13504 18944 13510 18956
rect 14093 18947 14151 18953
rect 14093 18944 14105 18947
rect 13504 18916 14105 18944
rect 13504 18904 13510 18916
rect 14093 18913 14105 18916
rect 14139 18913 14151 18947
rect 21361 18947 21419 18953
rect 21361 18944 21373 18947
rect 14093 18907 14151 18913
rect 20732 18916 21373 18944
rect 20732 18888 20760 18916
rect 21361 18913 21373 18916
rect 21407 18913 21419 18947
rect 21361 18907 21419 18913
rect 12069 18879 12127 18885
rect 12069 18845 12081 18879
rect 12115 18876 12127 18879
rect 12250 18876 12256 18888
rect 12115 18848 12256 18876
rect 12115 18845 12127 18848
rect 12069 18839 12127 18845
rect 12250 18836 12256 18848
rect 12308 18836 12314 18888
rect 13630 18876 13636 18888
rect 13591 18848 13636 18876
rect 13630 18836 13636 18848
rect 13688 18836 13694 18888
rect 13722 18836 13728 18888
rect 13780 18876 13786 18888
rect 14001 18879 14059 18885
rect 14001 18876 14013 18879
rect 13780 18848 14013 18876
rect 13780 18836 13786 18848
rect 14001 18845 14013 18848
rect 14047 18876 14059 18879
rect 14642 18876 14648 18888
rect 14047 18848 14648 18876
rect 14047 18845 14059 18848
rect 14001 18839 14059 18845
rect 14642 18836 14648 18848
rect 14700 18836 14706 18888
rect 15289 18879 15347 18885
rect 15289 18845 15301 18879
rect 15335 18876 15347 18879
rect 15562 18876 15568 18888
rect 15335 18848 15568 18876
rect 15335 18845 15347 18848
rect 15289 18839 15347 18845
rect 15562 18836 15568 18848
rect 15620 18836 15626 18888
rect 15746 18876 15752 18888
rect 15707 18848 15752 18876
rect 15746 18836 15752 18848
rect 15804 18836 15810 18888
rect 20714 18876 20720 18888
rect 20675 18848 20720 18876
rect 20714 18836 20720 18848
rect 20772 18836 20778 18888
rect 21266 18876 21272 18888
rect 21227 18848 21272 18876
rect 21266 18836 21272 18848
rect 21324 18836 21330 18888
rect 21450 18836 21456 18888
rect 21508 18876 21514 18888
rect 22480 18876 22508 19052
rect 22646 19040 22652 19052
rect 22704 19080 22710 19092
rect 22741 19083 22799 19089
rect 22741 19080 22753 19083
rect 22704 19052 22753 19080
rect 22704 19040 22710 19052
rect 22741 19049 22753 19052
rect 22787 19049 22799 19083
rect 22741 19043 22799 19049
rect 22554 18972 22560 19024
rect 22612 18972 22618 19024
rect 24949 19015 25007 19021
rect 24949 18981 24961 19015
rect 24995 19012 25007 19015
rect 25498 19012 25504 19024
rect 24995 18984 25504 19012
rect 24995 18981 25007 18984
rect 24949 18975 25007 18981
rect 25498 18972 25504 18984
rect 25556 18972 25562 19024
rect 22572 18944 22600 18972
rect 22986 18947 23044 18953
rect 22986 18944 22998 18947
rect 22572 18916 22998 18944
rect 22986 18913 22998 18916
rect 23032 18913 23044 18947
rect 22986 18907 23044 18913
rect 22557 18879 22615 18885
rect 22557 18876 22569 18879
rect 21508 18848 22569 18876
rect 21508 18836 21514 18848
rect 22557 18845 22569 18848
rect 22603 18845 22615 18879
rect 25130 18876 25136 18888
rect 25091 18848 25136 18876
rect 22557 18839 22615 18845
rect 25130 18836 25136 18848
rect 25188 18836 25194 18888
rect 1104 18786 26864 18808
rect 1104 18734 10315 18786
rect 10367 18734 10379 18786
rect 10431 18734 10443 18786
rect 10495 18734 10507 18786
rect 10559 18734 19648 18786
rect 19700 18734 19712 18786
rect 19764 18734 19776 18786
rect 19828 18734 19840 18786
rect 19892 18734 26864 18786
rect 1104 18712 26864 18734
rect 12161 18675 12219 18681
rect 12161 18641 12173 18675
rect 12207 18672 12219 18675
rect 12342 18672 12348 18684
rect 12207 18644 12348 18672
rect 12207 18641 12219 18644
rect 12161 18635 12219 18641
rect 12342 18632 12348 18644
rect 12400 18632 12406 18684
rect 13722 18672 13728 18684
rect 13683 18644 13728 18672
rect 13722 18632 13728 18644
rect 13780 18632 13786 18684
rect 14090 18672 14096 18684
rect 14051 18644 14096 18672
rect 14090 18632 14096 18644
rect 14148 18632 14154 18684
rect 15378 18672 15384 18684
rect 15339 18644 15384 18672
rect 15378 18632 15384 18644
rect 15436 18632 15442 18684
rect 15746 18672 15752 18684
rect 15707 18644 15752 18672
rect 15746 18632 15752 18644
rect 15804 18632 15810 18684
rect 20257 18675 20315 18681
rect 20257 18641 20269 18675
rect 20303 18672 20315 18675
rect 20990 18672 20996 18684
rect 20303 18644 20996 18672
rect 20303 18641 20315 18644
rect 20257 18635 20315 18641
rect 20990 18632 20996 18644
rect 21048 18632 21054 18684
rect 22554 18632 22560 18684
rect 22612 18672 22618 18684
rect 22741 18675 22799 18681
rect 22741 18672 22753 18675
rect 22612 18644 22753 18672
rect 22612 18632 22618 18644
rect 22741 18641 22753 18644
rect 22787 18672 22799 18675
rect 23017 18675 23075 18681
rect 23017 18672 23029 18675
rect 22787 18644 23029 18672
rect 22787 18641 22799 18644
rect 22741 18635 22799 18641
rect 23017 18641 23029 18644
rect 23063 18641 23075 18675
rect 23017 18635 23075 18641
rect 24026 18632 24032 18684
rect 24084 18672 24090 18684
rect 25317 18675 25375 18681
rect 25317 18672 25329 18675
rect 24084 18644 25329 18672
rect 24084 18632 24090 18644
rect 25317 18641 25329 18644
rect 25363 18641 25375 18675
rect 25317 18635 25375 18641
rect 16761 18607 16819 18613
rect 16761 18573 16773 18607
rect 16807 18604 16819 18607
rect 16850 18604 16856 18616
rect 16807 18576 16856 18604
rect 16807 18573 16819 18576
rect 16761 18567 16819 18573
rect 16850 18564 16856 18576
rect 16908 18564 16914 18616
rect 23937 18607 23995 18613
rect 23937 18573 23949 18607
rect 23983 18604 23995 18607
rect 24118 18604 24124 18616
rect 23983 18576 24124 18604
rect 23983 18573 23995 18576
rect 23937 18567 23995 18573
rect 24118 18564 24124 18576
rect 24176 18564 24182 18616
rect 17586 18496 17592 18548
rect 17644 18536 17650 18548
rect 18305 18539 18363 18545
rect 18305 18536 18317 18539
rect 17644 18508 18317 18536
rect 17644 18496 17650 18508
rect 18305 18505 18317 18508
rect 18351 18505 18363 18539
rect 21450 18536 21456 18548
rect 18305 18499 18363 18505
rect 21376 18508 21456 18536
rect 16390 18428 16396 18480
rect 16448 18468 16454 18480
rect 16853 18471 16911 18477
rect 16853 18468 16865 18471
rect 16448 18440 16865 18468
rect 16448 18428 16454 18440
rect 16853 18437 16865 18440
rect 16899 18437 16911 18471
rect 16853 18431 16911 18437
rect 17037 18471 17095 18477
rect 17037 18437 17049 18471
rect 17083 18468 17095 18471
rect 17604 18468 17632 18496
rect 18046 18468 18052 18480
rect 17083 18440 17632 18468
rect 18007 18440 18052 18468
rect 17083 18437 17095 18440
rect 17037 18431 17095 18437
rect 18046 18428 18052 18440
rect 18104 18428 18110 18480
rect 20349 18471 20407 18477
rect 20349 18437 20361 18471
rect 20395 18468 20407 18471
rect 20530 18468 20536 18480
rect 20395 18440 20536 18468
rect 20395 18437 20407 18440
rect 20349 18431 20407 18437
rect 20530 18428 20536 18440
rect 20588 18428 20594 18480
rect 20898 18428 20904 18480
rect 20956 18468 20962 18480
rect 21376 18477 21404 18508
rect 21450 18496 21456 18508
rect 21508 18496 21514 18548
rect 21628 18539 21686 18545
rect 21628 18505 21640 18539
rect 21674 18536 21686 18539
rect 22186 18536 22192 18548
rect 21674 18508 22192 18536
rect 21674 18505 21686 18508
rect 21628 18499 21686 18505
rect 22186 18496 22192 18508
rect 22244 18496 22250 18548
rect 23658 18496 23664 18548
rect 23716 18536 23722 18548
rect 24029 18539 24087 18545
rect 24029 18536 24041 18539
rect 23716 18508 24041 18536
rect 23716 18496 23722 18508
rect 24029 18505 24041 18508
rect 24075 18505 24087 18539
rect 24029 18499 24087 18505
rect 21361 18471 21419 18477
rect 21361 18468 21373 18471
rect 20956 18440 21373 18468
rect 20956 18428 20962 18440
rect 21361 18437 21373 18440
rect 21407 18437 21419 18471
rect 21361 18431 21419 18437
rect 24305 18471 24363 18477
rect 24305 18437 24317 18471
rect 24351 18468 24363 18471
rect 25130 18468 25136 18480
rect 24351 18440 25136 18468
rect 24351 18437 24363 18440
rect 24305 18431 24363 18437
rect 25130 18428 25136 18440
rect 25188 18428 25194 18480
rect 16114 18332 16120 18344
rect 16075 18304 16120 18332
rect 16114 18292 16120 18304
rect 16172 18292 16178 18344
rect 16393 18335 16451 18341
rect 16393 18301 16405 18335
rect 16439 18332 16451 18335
rect 16482 18332 16488 18344
rect 16439 18304 16488 18332
rect 16439 18301 16451 18304
rect 16393 18295 16451 18301
rect 16482 18292 16488 18304
rect 16540 18292 16546 18344
rect 19426 18332 19432 18344
rect 19387 18304 19432 18332
rect 19426 18292 19432 18304
rect 19484 18292 19490 18344
rect 20993 18335 21051 18341
rect 20993 18301 21005 18335
rect 21039 18332 21051 18335
rect 21358 18332 21364 18344
rect 21039 18304 21364 18332
rect 21039 18301 21051 18304
rect 20993 18295 21051 18301
rect 21358 18292 21364 18304
rect 21416 18292 21422 18344
rect 1104 18242 26864 18264
rect 1104 18190 5648 18242
rect 5700 18190 5712 18242
rect 5764 18190 5776 18242
rect 5828 18190 5840 18242
rect 5892 18190 14982 18242
rect 15034 18190 15046 18242
rect 15098 18190 15110 18242
rect 15162 18190 15174 18242
rect 15226 18190 24315 18242
rect 24367 18190 24379 18242
rect 24431 18190 24443 18242
rect 24495 18190 24507 18242
rect 24559 18190 26864 18242
rect 1104 18168 26864 18190
rect 15378 18128 15384 18140
rect 15339 18100 15384 18128
rect 15378 18088 15384 18100
rect 15436 18088 15442 18140
rect 16850 18128 16856 18140
rect 16811 18100 16856 18128
rect 16850 18088 16856 18100
rect 16908 18088 16914 18140
rect 17126 18088 17132 18140
rect 17184 18128 17190 18140
rect 17221 18131 17279 18137
rect 17221 18128 17233 18131
rect 17184 18100 17233 18128
rect 17184 18088 17190 18100
rect 17221 18097 17233 18100
rect 17267 18128 17279 18131
rect 17586 18128 17592 18140
rect 17267 18100 17592 18128
rect 17267 18097 17279 18100
rect 17221 18091 17279 18097
rect 17586 18088 17592 18100
rect 17644 18088 17650 18140
rect 22186 18088 22192 18140
rect 22244 18128 22250 18140
rect 22281 18131 22339 18137
rect 22281 18128 22293 18131
rect 22244 18100 22293 18128
rect 22244 18088 22250 18100
rect 22281 18097 22293 18100
rect 22327 18128 22339 18131
rect 22370 18128 22376 18140
rect 22327 18100 22376 18128
rect 22327 18097 22339 18100
rect 22281 18091 22339 18097
rect 22370 18088 22376 18100
rect 22428 18128 22434 18140
rect 22557 18131 22615 18137
rect 22557 18128 22569 18131
rect 22428 18100 22569 18128
rect 22428 18088 22434 18100
rect 22557 18097 22569 18100
rect 22603 18097 22615 18131
rect 22557 18091 22615 18097
rect 23658 18088 23664 18140
rect 23716 18128 23722 18140
rect 24581 18131 24639 18137
rect 24581 18128 24593 18131
rect 23716 18100 24593 18128
rect 23716 18088 23722 18100
rect 24581 18097 24593 18100
rect 24627 18097 24639 18131
rect 25314 18128 25320 18140
rect 25275 18100 25320 18128
rect 24581 18091 24639 18097
rect 25314 18088 25320 18100
rect 25372 18088 25378 18140
rect 15105 17995 15163 18001
rect 15105 17961 15117 17995
rect 15151 17992 15163 17995
rect 15930 17992 15936 18004
rect 15151 17964 15936 17992
rect 15151 17961 15163 17964
rect 15105 17955 15163 17961
rect 15930 17952 15936 17964
rect 15988 17952 15994 18004
rect 16390 17924 16396 17936
rect 16351 17896 16396 17924
rect 16390 17884 16396 17896
rect 16448 17884 16454 17936
rect 18417 17927 18475 17933
rect 18417 17924 18429 17927
rect 18248 17896 18429 17924
rect 15749 17859 15807 17865
rect 15749 17825 15761 17859
rect 15795 17856 15807 17859
rect 16114 17856 16120 17868
rect 15795 17828 16120 17856
rect 15795 17825 15807 17828
rect 15749 17819 15807 17825
rect 16114 17816 16120 17828
rect 16172 17816 16178 17868
rect 14737 17791 14795 17797
rect 14737 17757 14749 17791
rect 14783 17788 14795 17791
rect 15286 17788 15292 17800
rect 14783 17760 15292 17788
rect 14783 17757 14795 17760
rect 14737 17751 14795 17757
rect 15286 17748 15292 17760
rect 15344 17788 15350 17800
rect 15841 17791 15899 17797
rect 15841 17788 15853 17791
rect 15344 17760 15853 17788
rect 15344 17748 15350 17760
rect 15841 17757 15853 17760
rect 15887 17757 15899 17791
rect 15841 17751 15899 17757
rect 17957 17791 18015 17797
rect 17957 17757 17969 17791
rect 18003 17788 18015 17791
rect 18138 17788 18144 17800
rect 18003 17760 18144 17788
rect 18003 17757 18015 17760
rect 17957 17751 18015 17757
rect 18138 17748 18144 17760
rect 18196 17788 18202 17800
rect 18248 17797 18276 17896
rect 18417 17893 18429 17896
rect 18463 17893 18475 17927
rect 20898 17924 20904 17936
rect 18417 17887 18475 17893
rect 20732 17896 20904 17924
rect 18598 17816 18604 17868
rect 18656 17865 18662 17868
rect 18656 17859 18720 17865
rect 18656 17825 18674 17859
rect 18708 17825 18720 17859
rect 18656 17819 18720 17825
rect 18656 17816 18662 17819
rect 19426 17816 19432 17868
rect 19484 17856 19490 17868
rect 20073 17859 20131 17865
rect 20073 17856 20085 17859
rect 19484 17828 20085 17856
rect 19484 17816 19490 17828
rect 20073 17825 20085 17828
rect 20119 17825 20131 17859
rect 20073 17819 20131 17825
rect 20732 17800 20760 17896
rect 20898 17884 20904 17896
rect 20956 17884 20962 17936
rect 20990 17884 20996 17936
rect 21048 17924 21054 17936
rect 21157 17927 21215 17933
rect 21157 17924 21169 17927
rect 21048 17896 21169 17924
rect 21048 17884 21054 17896
rect 21157 17893 21169 17896
rect 21203 17893 21215 17927
rect 23845 17927 23903 17933
rect 23845 17924 23857 17927
rect 21157 17887 21215 17893
rect 23676 17896 23857 17924
rect 23676 17800 23704 17896
rect 23845 17893 23857 17896
rect 23891 17893 23903 17927
rect 25130 17924 25136 17936
rect 25091 17896 25136 17924
rect 23845 17887 23903 17893
rect 25130 17884 25136 17896
rect 25188 17924 25194 17936
rect 25685 17927 25743 17933
rect 25685 17924 25697 17927
rect 25188 17896 25697 17924
rect 25188 17884 25194 17896
rect 25685 17893 25697 17896
rect 25731 17893 25743 17927
rect 25685 17887 25743 17893
rect 24118 17856 24124 17868
rect 24079 17828 24124 17856
rect 24118 17816 24124 17828
rect 24176 17816 24182 17868
rect 18233 17791 18291 17797
rect 18233 17788 18245 17791
rect 18196 17760 18245 17788
rect 18196 17748 18202 17760
rect 18233 17757 18245 17760
rect 18279 17757 18291 17791
rect 18233 17751 18291 17757
rect 19797 17791 19855 17797
rect 19797 17757 19809 17791
rect 19843 17788 19855 17791
rect 19978 17788 19984 17800
rect 19843 17760 19984 17788
rect 19843 17757 19855 17760
rect 19797 17751 19855 17757
rect 19978 17748 19984 17760
rect 20036 17748 20042 17800
rect 20714 17788 20720 17800
rect 20675 17760 20720 17788
rect 20714 17748 20720 17760
rect 20772 17748 20778 17800
rect 23658 17788 23664 17800
rect 23619 17760 23664 17788
rect 23658 17748 23664 17760
rect 23716 17748 23722 17800
rect 1104 17698 26864 17720
rect 1104 17646 10315 17698
rect 10367 17646 10379 17698
rect 10431 17646 10443 17698
rect 10495 17646 10507 17698
rect 10559 17646 19648 17698
rect 19700 17646 19712 17698
rect 19764 17646 19776 17698
rect 19828 17646 19840 17698
rect 19892 17646 26864 17698
rect 1104 17624 26864 17646
rect 14553 17587 14611 17593
rect 14553 17553 14565 17587
rect 14599 17584 14611 17587
rect 14642 17584 14648 17596
rect 14599 17556 14648 17584
rect 14599 17553 14611 17556
rect 14553 17547 14611 17553
rect 14642 17544 14648 17556
rect 14700 17544 14706 17596
rect 17126 17584 17132 17596
rect 17087 17556 17132 17584
rect 17126 17544 17132 17556
rect 17184 17544 17190 17596
rect 18506 17584 18512 17596
rect 18467 17556 18512 17584
rect 18506 17544 18512 17556
rect 18564 17544 18570 17596
rect 20990 17584 20996 17596
rect 20951 17556 20996 17584
rect 20990 17544 20996 17556
rect 21048 17544 21054 17596
rect 21818 17584 21824 17596
rect 21779 17556 21824 17584
rect 21818 17544 21824 17556
rect 21876 17544 21882 17596
rect 22094 17544 22100 17596
rect 22152 17584 22158 17596
rect 22281 17587 22339 17593
rect 22281 17584 22293 17587
rect 22152 17556 22293 17584
rect 22152 17544 22158 17556
rect 22281 17553 22293 17556
rect 22327 17553 22339 17587
rect 24762 17584 24768 17596
rect 24723 17556 24768 17584
rect 22281 17547 22339 17553
rect 24762 17544 24768 17556
rect 24820 17544 24826 17596
rect 14734 17476 14740 17528
rect 14792 17516 14798 17528
rect 14792 17488 15792 17516
rect 14792 17476 14798 17488
rect 15764 17460 15792 17488
rect 15930 17476 15936 17528
rect 15988 17525 15994 17528
rect 15988 17519 16052 17525
rect 15988 17485 16006 17519
rect 16040 17485 16052 17519
rect 20714 17516 20720 17528
rect 15988 17479 16052 17485
rect 19628 17488 20720 17516
rect 15988 17476 15994 17479
rect 14182 17408 14188 17460
rect 14240 17448 14246 17460
rect 14645 17451 14703 17457
rect 14645 17448 14657 17451
rect 14240 17420 14657 17448
rect 14240 17408 14246 17420
rect 14645 17417 14657 17420
rect 14691 17417 14703 17451
rect 15746 17448 15752 17460
rect 15659 17420 15752 17448
rect 14645 17411 14703 17417
rect 15746 17408 15752 17420
rect 15804 17408 15810 17460
rect 18046 17408 18052 17460
rect 18104 17448 18110 17460
rect 18414 17448 18420 17460
rect 18104 17420 18420 17448
rect 18104 17408 18110 17420
rect 18414 17408 18420 17420
rect 18472 17408 18478 17460
rect 19334 17408 19340 17460
rect 19392 17448 19398 17460
rect 19628 17457 19656 17488
rect 20714 17476 20720 17488
rect 20772 17516 20778 17528
rect 21361 17519 21419 17525
rect 21361 17516 21373 17519
rect 20772 17488 21373 17516
rect 20772 17476 20778 17488
rect 21361 17485 21373 17488
rect 21407 17485 21419 17519
rect 21361 17479 21419 17485
rect 19886 17457 19892 17460
rect 19613 17451 19671 17457
rect 19613 17448 19625 17451
rect 19392 17420 19625 17448
rect 19392 17408 19398 17420
rect 19613 17417 19625 17420
rect 19659 17417 19671 17451
rect 19880 17448 19892 17457
rect 19847 17420 19892 17448
rect 19613 17411 19671 17417
rect 19880 17411 19892 17420
rect 19886 17408 19892 17411
rect 19944 17408 19950 17460
rect 22186 17448 22192 17460
rect 22147 17420 22192 17448
rect 22186 17408 22192 17420
rect 22244 17408 22250 17460
rect 24118 17408 24124 17460
rect 24176 17448 24182 17460
rect 24581 17451 24639 17457
rect 24581 17448 24593 17451
rect 24176 17420 24593 17448
rect 24176 17408 24182 17420
rect 24581 17417 24593 17420
rect 24627 17448 24639 17451
rect 25038 17448 25044 17460
rect 24627 17420 25044 17448
rect 24627 17417 24639 17420
rect 24581 17411 24639 17417
rect 25038 17408 25044 17420
rect 25096 17408 25102 17460
rect 14734 17380 14740 17392
rect 14695 17352 14740 17380
rect 14734 17340 14740 17352
rect 14792 17340 14798 17392
rect 18598 17380 18604 17392
rect 18559 17352 18604 17380
rect 18598 17340 18604 17352
rect 18656 17380 18662 17392
rect 19426 17380 19432 17392
rect 18656 17352 19432 17380
rect 18656 17340 18662 17352
rect 19426 17340 19432 17352
rect 19484 17340 19490 17392
rect 22370 17340 22376 17392
rect 22428 17380 22434 17392
rect 22428 17352 22473 17380
rect 22428 17340 22434 17352
rect 13998 17204 14004 17256
rect 14056 17244 14062 17256
rect 14185 17247 14243 17253
rect 14185 17244 14197 17247
rect 14056 17216 14197 17244
rect 14056 17204 14062 17216
rect 14185 17213 14197 17216
rect 14231 17213 14243 17247
rect 15378 17244 15384 17256
rect 15339 17216 15384 17244
rect 14185 17207 14243 17213
rect 15378 17204 15384 17216
rect 15436 17204 15442 17256
rect 18049 17247 18107 17253
rect 18049 17213 18061 17247
rect 18095 17244 18107 17247
rect 18874 17244 18880 17256
rect 18095 17216 18880 17244
rect 18095 17213 18107 17216
rect 18049 17207 18107 17213
rect 18874 17204 18880 17216
rect 18932 17204 18938 17256
rect 19058 17244 19064 17256
rect 19019 17216 19064 17244
rect 19058 17204 19064 17216
rect 19116 17204 19122 17256
rect 1104 17154 26864 17176
rect 1104 17102 5648 17154
rect 5700 17102 5712 17154
rect 5764 17102 5776 17154
rect 5828 17102 5840 17154
rect 5892 17102 14982 17154
rect 15034 17102 15046 17154
rect 15098 17102 15110 17154
rect 15162 17102 15174 17154
rect 15226 17102 24315 17154
rect 24367 17102 24379 17154
rect 24431 17102 24443 17154
rect 24495 17102 24507 17154
rect 24559 17102 26864 17154
rect 1104 17080 26864 17102
rect 14826 17000 14832 17052
rect 14884 17040 14890 17052
rect 15013 17043 15071 17049
rect 15013 17040 15025 17043
rect 14884 17012 15025 17040
rect 14884 17000 14890 17012
rect 15013 17009 15025 17012
rect 15059 17009 15071 17043
rect 15013 17003 15071 17009
rect 15028 16904 15056 17003
rect 15930 17000 15936 17052
rect 15988 17040 15994 17052
rect 16298 17040 16304 17052
rect 15988 17012 16304 17040
rect 15988 17000 15994 17012
rect 16298 17000 16304 17012
rect 16356 17040 16362 17052
rect 16669 17043 16727 17049
rect 16669 17040 16681 17043
rect 16356 17012 16681 17040
rect 16356 17000 16362 17012
rect 16669 17009 16681 17012
rect 16715 17009 16727 17043
rect 16669 17003 16727 17009
rect 17497 17043 17555 17049
rect 17497 17009 17509 17043
rect 17543 17040 17555 17043
rect 18598 17040 18604 17052
rect 17543 17012 18604 17040
rect 17543 17009 17555 17012
rect 17497 17003 17555 17009
rect 18598 17000 18604 17012
rect 18656 17000 18662 17052
rect 19334 17000 19340 17052
rect 19392 17040 19398 17052
rect 19613 17043 19671 17049
rect 19613 17040 19625 17043
rect 19392 17012 19625 17040
rect 19392 17000 19398 17012
rect 19613 17009 19625 17012
rect 19659 17009 19671 17043
rect 19613 17003 19671 17009
rect 20530 17000 20536 17052
rect 20588 17040 20594 17052
rect 21361 17043 21419 17049
rect 21361 17040 21373 17043
rect 20588 17012 21373 17040
rect 20588 17000 20594 17012
rect 21361 17009 21373 17012
rect 21407 17040 21419 17043
rect 22186 17040 22192 17052
rect 21407 17012 22192 17040
rect 21407 17009 21419 17012
rect 21361 17003 21419 17009
rect 22186 17000 22192 17012
rect 22244 17000 22250 17052
rect 25038 17040 25044 17052
rect 24999 17012 25044 17040
rect 25038 17000 25044 17012
rect 25096 17000 25102 17052
rect 25406 17040 25412 17052
rect 25367 17012 25412 17040
rect 25406 17000 25412 17012
rect 25464 17000 25470 17052
rect 18046 16972 18052 16984
rect 18007 16944 18052 16972
rect 18046 16932 18052 16944
rect 18104 16932 18110 16984
rect 15289 16907 15347 16913
rect 15289 16904 15301 16907
rect 15028 16876 15301 16904
rect 15289 16873 15301 16876
rect 15335 16873 15347 16907
rect 18414 16904 18420 16916
rect 18375 16876 18420 16904
rect 15289 16867 15347 16873
rect 18414 16864 18420 16876
rect 18472 16864 18478 16916
rect 18616 16904 18644 17000
rect 22094 16932 22100 16984
rect 22152 16972 22158 16984
rect 23293 16975 23351 16981
rect 23293 16972 23305 16975
rect 22152 16944 23305 16972
rect 22152 16932 22158 16944
rect 23293 16941 23305 16944
rect 23339 16941 23351 16975
rect 23293 16935 23351 16941
rect 19153 16907 19211 16913
rect 19153 16904 19165 16907
rect 18616 16876 19165 16904
rect 19153 16873 19165 16876
rect 19199 16873 19211 16907
rect 19153 16867 19211 16873
rect 22278 16864 22284 16916
rect 22336 16904 22342 16916
rect 22465 16907 22523 16913
rect 22465 16904 22477 16907
rect 22336 16876 22477 16904
rect 22336 16864 22342 16876
rect 22465 16873 22477 16876
rect 22511 16873 22523 16907
rect 22465 16867 22523 16873
rect 14182 16836 14188 16848
rect 14143 16808 14188 16836
rect 14182 16796 14188 16808
rect 14240 16796 14246 16848
rect 15378 16796 15384 16848
rect 15436 16836 15442 16848
rect 15545 16839 15603 16845
rect 15545 16836 15557 16839
rect 15436 16808 15557 16836
rect 15436 16796 15442 16808
rect 15545 16805 15557 16808
rect 15591 16805 15603 16839
rect 15545 16799 15603 16805
rect 17589 16839 17647 16845
rect 17589 16805 17601 16839
rect 17635 16836 17647 16839
rect 18969 16839 19027 16845
rect 18969 16836 18981 16839
rect 17635 16808 18981 16836
rect 17635 16805 17647 16808
rect 17589 16799 17647 16805
rect 18969 16805 18981 16808
rect 19015 16836 19027 16839
rect 19058 16836 19064 16848
rect 19015 16808 19064 16836
rect 19015 16805 19027 16808
rect 18969 16799 19027 16805
rect 19058 16796 19064 16808
rect 19116 16796 19122 16848
rect 23934 16836 23940 16848
rect 23895 16808 23940 16836
rect 23934 16796 23940 16808
rect 23992 16796 23998 16848
rect 24213 16839 24271 16845
rect 24213 16805 24225 16839
rect 24259 16836 24271 16839
rect 25225 16839 25283 16845
rect 25225 16836 25237 16839
rect 24259 16808 25237 16836
rect 24259 16805 24271 16808
rect 24213 16799 24271 16805
rect 25225 16805 25237 16808
rect 25271 16836 25283 16839
rect 25777 16839 25835 16845
rect 25777 16836 25789 16839
rect 25271 16808 25789 16836
rect 25271 16805 25283 16808
rect 25225 16799 25283 16805
rect 25777 16805 25789 16808
rect 25823 16805 25835 16839
rect 25777 16799 25835 16805
rect 13909 16771 13967 16777
rect 13909 16737 13921 16771
rect 13955 16768 13967 16771
rect 14734 16768 14740 16780
rect 13955 16740 14740 16768
rect 13955 16737 13967 16740
rect 13909 16731 13967 16737
rect 14734 16728 14740 16740
rect 14792 16728 14798 16780
rect 18414 16728 18420 16780
rect 18472 16768 18478 16780
rect 18472 16740 19104 16768
rect 18472 16728 18478 16740
rect 19076 16712 19104 16740
rect 19334 16728 19340 16780
rect 19392 16768 19398 16780
rect 19886 16768 19892 16780
rect 19392 16740 19892 16768
rect 19392 16728 19398 16740
rect 19886 16728 19892 16740
rect 19944 16768 19950 16780
rect 19981 16771 20039 16777
rect 19981 16768 19993 16771
rect 19944 16740 19993 16768
rect 19944 16728 19950 16740
rect 19981 16737 19993 16740
rect 20027 16737 20039 16771
rect 19981 16731 20039 16737
rect 21726 16728 21732 16780
rect 21784 16768 21790 16780
rect 21821 16771 21879 16777
rect 21821 16768 21833 16771
rect 21784 16740 21833 16768
rect 21784 16728 21790 16740
rect 21821 16737 21833 16740
rect 21867 16768 21879 16771
rect 22281 16771 22339 16777
rect 22281 16768 22293 16771
rect 21867 16740 22293 16768
rect 21867 16737 21879 16740
rect 21821 16731 21879 16737
rect 22281 16737 22293 16740
rect 22327 16768 22339 16771
rect 23658 16768 23664 16780
rect 22327 16740 23664 16768
rect 22327 16737 22339 16740
rect 22281 16731 22339 16737
rect 23658 16728 23664 16740
rect 23716 16728 23722 16780
rect 23952 16768 23980 16796
rect 24673 16771 24731 16777
rect 24673 16768 24685 16771
rect 23952 16740 24685 16768
rect 24673 16737 24685 16740
rect 24719 16737 24731 16771
rect 24673 16731 24731 16737
rect 14642 16700 14648 16712
rect 14603 16672 14648 16700
rect 14642 16660 14648 16672
rect 14700 16660 14706 16712
rect 18598 16700 18604 16712
rect 18559 16672 18604 16700
rect 18598 16660 18604 16672
rect 18656 16660 18662 16712
rect 19058 16700 19064 16712
rect 18971 16672 19064 16700
rect 19058 16660 19064 16672
rect 19116 16660 19122 16712
rect 21910 16700 21916 16712
rect 21871 16672 21916 16700
rect 21910 16660 21916 16672
rect 21968 16660 21974 16712
rect 22370 16660 22376 16712
rect 22428 16700 22434 16712
rect 22925 16703 22983 16709
rect 22925 16700 22937 16703
rect 22428 16672 22937 16700
rect 22428 16660 22434 16672
rect 22925 16669 22937 16672
rect 22971 16669 22983 16703
rect 22925 16663 22983 16669
rect 1104 16610 26864 16632
rect 1104 16558 10315 16610
rect 10367 16558 10379 16610
rect 10431 16558 10443 16610
rect 10495 16558 10507 16610
rect 10559 16558 19648 16610
rect 19700 16558 19712 16610
rect 19764 16558 19776 16610
rect 19828 16558 19840 16610
rect 19892 16558 26864 16610
rect 1104 16536 26864 16558
rect 15378 16456 15384 16508
rect 15436 16496 15442 16508
rect 15657 16499 15715 16505
rect 15657 16496 15669 16499
rect 15436 16468 15669 16496
rect 15436 16456 15442 16468
rect 15657 16465 15669 16468
rect 15703 16496 15715 16499
rect 15838 16496 15844 16508
rect 15703 16468 15844 16496
rect 15703 16465 15715 16468
rect 15657 16459 15715 16465
rect 15838 16456 15844 16468
rect 15896 16456 15902 16508
rect 16298 16496 16304 16508
rect 16259 16468 16304 16496
rect 16298 16456 16304 16468
rect 16356 16456 16362 16508
rect 18325 16499 18383 16505
rect 18325 16465 18337 16499
rect 18371 16496 18383 16499
rect 18506 16496 18512 16508
rect 18371 16468 18512 16496
rect 18371 16465 18383 16468
rect 18325 16459 18383 16465
rect 18506 16456 18512 16468
rect 18564 16456 18570 16508
rect 18690 16496 18696 16508
rect 18651 16468 18696 16496
rect 18690 16456 18696 16468
rect 18748 16456 18754 16508
rect 18874 16456 18880 16508
rect 18932 16496 18938 16508
rect 19153 16499 19211 16505
rect 19153 16496 19165 16499
rect 18932 16468 19165 16496
rect 18932 16456 18938 16468
rect 19153 16465 19165 16468
rect 19199 16496 19211 16499
rect 19426 16496 19432 16508
rect 19199 16468 19432 16496
rect 19199 16465 19211 16468
rect 19153 16459 19211 16465
rect 19426 16456 19432 16468
rect 19484 16456 19490 16508
rect 20717 16499 20775 16505
rect 20717 16465 20729 16499
rect 20763 16496 20775 16499
rect 22370 16496 22376 16508
rect 20763 16468 22376 16496
rect 20763 16465 20775 16468
rect 20717 16459 20775 16465
rect 22370 16456 22376 16468
rect 22428 16456 22434 16508
rect 25406 16496 25412 16508
rect 25367 16468 25412 16496
rect 25406 16456 25412 16468
rect 25464 16456 25470 16508
rect 14544 16431 14602 16437
rect 14544 16397 14556 16431
rect 14590 16428 14602 16431
rect 14734 16428 14740 16440
rect 14590 16400 14740 16428
rect 14590 16397 14602 16400
rect 14544 16391 14602 16397
rect 14734 16388 14740 16400
rect 14792 16388 14798 16440
rect 15856 16428 15884 16456
rect 16945 16431 17003 16437
rect 16945 16428 16957 16431
rect 15856 16400 16957 16428
rect 16945 16397 16957 16400
rect 16991 16397 17003 16431
rect 21174 16428 21180 16440
rect 21135 16400 21180 16428
rect 16945 16391 17003 16397
rect 21174 16388 21180 16400
rect 21232 16388 21238 16440
rect 21913 16431 21971 16437
rect 21913 16397 21925 16431
rect 21959 16428 21971 16431
rect 22462 16428 22468 16440
rect 21959 16400 22468 16428
rect 21959 16397 21971 16400
rect 21913 16391 21971 16397
rect 22462 16388 22468 16400
rect 22520 16388 22526 16440
rect 15746 16320 15752 16372
rect 15804 16360 15810 16372
rect 15933 16363 15991 16369
rect 15933 16360 15945 16363
rect 15804 16332 15945 16360
rect 15804 16320 15810 16332
rect 15933 16329 15945 16332
rect 15979 16329 15991 16363
rect 15933 16323 15991 16329
rect 18598 16320 18604 16372
rect 18656 16360 18662 16372
rect 19061 16363 19119 16369
rect 19061 16360 19073 16363
rect 18656 16332 19073 16360
rect 18656 16320 18662 16332
rect 19061 16329 19073 16332
rect 19107 16329 19119 16363
rect 19061 16323 19119 16329
rect 21085 16363 21143 16369
rect 21085 16329 21097 16363
rect 21131 16360 21143 16363
rect 21542 16360 21548 16372
rect 21131 16332 21548 16360
rect 21131 16329 21143 16332
rect 21085 16323 21143 16329
rect 21542 16320 21548 16332
rect 21600 16320 21606 16372
rect 22554 16360 22560 16372
rect 22515 16332 22560 16360
rect 22554 16320 22560 16332
rect 22612 16320 22618 16372
rect 23750 16320 23756 16372
rect 23808 16360 23814 16372
rect 23937 16363 23995 16369
rect 23937 16360 23949 16363
rect 23808 16332 23949 16360
rect 23808 16320 23814 16332
rect 23937 16329 23949 16332
rect 23983 16329 23995 16363
rect 23937 16323 23995 16329
rect 24213 16363 24271 16369
rect 24213 16329 24225 16363
rect 24259 16360 24271 16363
rect 25222 16360 25228 16372
rect 24259 16332 25228 16360
rect 24259 16329 24271 16332
rect 24213 16323 24271 16329
rect 25222 16320 25228 16332
rect 25280 16320 25286 16372
rect 14274 16292 14280 16304
rect 14235 16264 14280 16292
rect 14274 16252 14280 16264
rect 14332 16252 14338 16304
rect 16482 16292 16488 16304
rect 16443 16264 16488 16292
rect 16482 16252 16488 16264
rect 16540 16252 16546 16304
rect 19245 16295 19303 16301
rect 19245 16261 19257 16295
rect 19291 16292 19303 16295
rect 19334 16292 19340 16304
rect 19291 16264 19340 16292
rect 19291 16261 19303 16264
rect 19245 16255 19303 16261
rect 18782 16184 18788 16236
rect 18840 16224 18846 16236
rect 19260 16224 19288 16255
rect 19334 16252 19340 16264
rect 19392 16252 19398 16304
rect 21266 16252 21272 16304
rect 21324 16292 21330 16304
rect 22278 16292 22284 16304
rect 21324 16264 21369 16292
rect 22239 16264 22284 16292
rect 21324 16252 21330 16264
rect 22278 16252 22284 16264
rect 22336 16252 22342 16304
rect 23566 16252 23572 16304
rect 23624 16292 23630 16304
rect 24118 16292 24124 16304
rect 23624 16264 24124 16292
rect 23624 16252 23630 16264
rect 24118 16252 24124 16264
rect 24176 16252 24182 16304
rect 18840 16196 19288 16224
rect 18840 16184 18846 16196
rect 23474 16184 23480 16236
rect 23532 16224 23538 16236
rect 23934 16224 23940 16236
rect 23532 16196 23940 16224
rect 23532 16184 23538 16196
rect 23934 16184 23940 16196
rect 23992 16184 23998 16236
rect 1104 16066 26864 16088
rect 1104 16014 5648 16066
rect 5700 16014 5712 16066
rect 5764 16014 5776 16066
rect 5828 16014 5840 16066
rect 5892 16014 14982 16066
rect 15034 16014 15046 16066
rect 15098 16014 15110 16066
rect 15162 16014 15174 16066
rect 15226 16014 24315 16066
rect 24367 16014 24379 16066
rect 24431 16014 24443 16066
rect 24495 16014 24507 16066
rect 24559 16014 26864 16066
rect 1104 15992 26864 16014
rect 13998 15952 14004 15964
rect 13959 15924 14004 15952
rect 13998 15912 14004 15924
rect 14056 15912 14062 15964
rect 15286 15952 15292 15964
rect 15247 15924 15292 15952
rect 15286 15912 15292 15924
rect 15344 15912 15350 15964
rect 16393 15955 16451 15961
rect 16393 15921 16405 15955
rect 16439 15952 16451 15955
rect 16482 15952 16488 15964
rect 16439 15924 16488 15952
rect 16439 15921 16451 15924
rect 16393 15915 16451 15921
rect 16482 15912 16488 15924
rect 16540 15912 16546 15964
rect 19426 15912 19432 15964
rect 19484 15952 19490 15964
rect 19981 15955 20039 15961
rect 19981 15952 19993 15955
rect 19484 15924 19993 15952
rect 19484 15912 19490 15924
rect 19981 15921 19993 15924
rect 20027 15921 20039 15955
rect 21174 15952 21180 15964
rect 21135 15924 21180 15952
rect 19981 15915 20039 15921
rect 21174 15912 21180 15924
rect 21232 15912 21238 15964
rect 23750 15912 23756 15964
rect 23808 15952 23814 15964
rect 23937 15955 23995 15961
rect 23937 15952 23949 15955
rect 23808 15924 23949 15952
rect 23808 15912 23814 15924
rect 23937 15921 23949 15924
rect 23983 15921 23995 15955
rect 24762 15952 24768 15964
rect 24723 15924 24768 15952
rect 23937 15915 23995 15921
rect 24762 15912 24768 15924
rect 24820 15912 24826 15964
rect 25222 15912 25228 15964
rect 25280 15952 25286 15964
rect 25501 15955 25559 15961
rect 25501 15952 25513 15955
rect 25280 15924 25513 15952
rect 25280 15912 25286 15924
rect 25501 15921 25513 15924
rect 25547 15921 25559 15955
rect 25501 15915 25559 15921
rect 14016 15816 14044 15912
rect 16114 15844 16120 15896
rect 16172 15884 16178 15896
rect 16853 15887 16911 15893
rect 16853 15884 16865 15887
rect 16172 15856 16865 15884
rect 16172 15844 16178 15856
rect 16853 15853 16865 15856
rect 16899 15853 16911 15887
rect 16853 15847 16911 15853
rect 15749 15819 15807 15825
rect 15749 15816 15761 15819
rect 14016 15788 15761 15816
rect 15749 15785 15761 15788
rect 15795 15785 15807 15819
rect 15749 15779 15807 15785
rect 15838 15776 15844 15828
rect 15896 15816 15902 15828
rect 17405 15819 17463 15825
rect 17405 15816 17417 15819
rect 15896 15788 17417 15816
rect 15896 15776 15902 15788
rect 17405 15785 17417 15788
rect 17451 15785 17463 15819
rect 17405 15779 17463 15785
rect 18509 15819 18567 15825
rect 18509 15785 18521 15819
rect 18555 15816 18567 15819
rect 19153 15819 19211 15825
rect 19153 15816 19165 15819
rect 18555 15788 19165 15816
rect 18555 15785 18567 15788
rect 18509 15779 18567 15785
rect 19153 15785 19165 15788
rect 19199 15816 19211 15819
rect 19242 15816 19248 15828
rect 19199 15788 19248 15816
rect 19199 15785 19211 15788
rect 19153 15779 19211 15785
rect 19242 15776 19248 15788
rect 19300 15776 19306 15828
rect 20714 15776 20720 15828
rect 20772 15816 20778 15828
rect 22005 15819 22063 15825
rect 22005 15816 22017 15819
rect 20772 15788 22017 15816
rect 20772 15776 20778 15788
rect 22005 15785 22017 15788
rect 22051 15785 22063 15819
rect 22005 15779 22063 15785
rect 16482 15708 16488 15760
rect 16540 15748 16546 15760
rect 17221 15751 17279 15757
rect 17221 15748 17233 15751
rect 16540 15720 17233 15748
rect 16540 15708 16546 15720
rect 17221 15717 17233 15720
rect 17267 15717 17279 15751
rect 17221 15711 17279 15717
rect 17313 15751 17371 15757
rect 17313 15717 17325 15751
rect 17359 15748 17371 15751
rect 17862 15748 17868 15760
rect 17359 15720 17868 15748
rect 17359 15717 17371 15720
rect 17313 15711 17371 15717
rect 16761 15683 16819 15689
rect 16761 15649 16773 15683
rect 16807 15680 16819 15683
rect 17328 15680 17356 15711
rect 17862 15708 17868 15720
rect 17920 15708 17926 15760
rect 22020 15748 22048 15779
rect 22189 15751 22247 15757
rect 22189 15748 22201 15751
rect 22020 15720 22201 15748
rect 22189 15717 22201 15720
rect 22235 15717 22247 15751
rect 22189 15711 22247 15717
rect 22278 15708 22284 15760
rect 22336 15748 22342 15760
rect 22445 15751 22503 15757
rect 22445 15748 22457 15751
rect 22336 15720 22457 15748
rect 22336 15708 22342 15720
rect 22445 15717 22457 15720
rect 22491 15717 22503 15751
rect 22445 15711 22503 15717
rect 24581 15751 24639 15757
rect 24581 15717 24593 15751
rect 24627 15748 24639 15751
rect 24670 15748 24676 15760
rect 24627 15720 24676 15748
rect 24627 15717 24639 15720
rect 24581 15711 24639 15717
rect 24670 15708 24676 15720
rect 24728 15748 24734 15760
rect 25133 15751 25191 15757
rect 25133 15748 25145 15751
rect 24728 15720 25145 15748
rect 24728 15708 24734 15720
rect 25133 15717 25145 15720
rect 25179 15717 25191 15751
rect 25133 15711 25191 15717
rect 16807 15652 17356 15680
rect 18141 15683 18199 15689
rect 16807 15649 16819 15652
rect 16761 15643 16819 15649
rect 18141 15649 18153 15683
rect 18187 15680 18199 15683
rect 18874 15680 18880 15692
rect 18187 15652 18880 15680
rect 18187 15649 18199 15652
rect 18141 15643 18199 15649
rect 18874 15640 18880 15652
rect 18932 15680 18938 15692
rect 19061 15683 19119 15689
rect 19061 15680 19073 15683
rect 18932 15652 19073 15680
rect 18932 15640 18938 15652
rect 19061 15649 19073 15652
rect 19107 15649 19119 15683
rect 19061 15643 19119 15649
rect 20346 15640 20352 15692
rect 20404 15680 20410 15692
rect 20717 15683 20775 15689
rect 20717 15680 20729 15683
rect 20404 15652 20729 15680
rect 20404 15640 20410 15652
rect 20717 15649 20729 15652
rect 20763 15680 20775 15683
rect 21266 15680 21272 15692
rect 20763 15652 21272 15680
rect 20763 15649 20775 15652
rect 20717 15643 20775 15649
rect 21266 15640 21272 15652
rect 21324 15680 21330 15692
rect 21726 15680 21732 15692
rect 21324 15652 21732 15680
rect 21324 15640 21330 15652
rect 21726 15640 21732 15652
rect 21784 15640 21790 15692
rect 13630 15572 13636 15624
rect 13688 15612 13694 15624
rect 14274 15612 14280 15624
rect 13688 15584 14280 15612
rect 13688 15572 13694 15584
rect 14274 15572 14280 15584
rect 14332 15572 14338 15624
rect 14734 15612 14740 15624
rect 14695 15584 14740 15612
rect 14734 15572 14740 15584
rect 14792 15572 14798 15624
rect 15105 15615 15163 15621
rect 15105 15581 15117 15615
rect 15151 15612 15163 15615
rect 15654 15612 15660 15624
rect 15151 15584 15660 15612
rect 15151 15581 15163 15584
rect 15105 15575 15163 15581
rect 15654 15572 15660 15584
rect 15712 15572 15718 15624
rect 18601 15615 18659 15621
rect 18601 15581 18613 15615
rect 18647 15612 18659 15615
rect 18690 15612 18696 15624
rect 18647 15584 18696 15612
rect 18647 15581 18659 15584
rect 18601 15575 18659 15581
rect 18690 15572 18696 15584
rect 18748 15572 18754 15624
rect 18966 15612 18972 15624
rect 18927 15584 18972 15612
rect 18966 15572 18972 15584
rect 19024 15612 19030 15624
rect 19613 15615 19671 15621
rect 19613 15612 19625 15615
rect 19024 15584 19625 15612
rect 19024 15572 19030 15584
rect 19613 15581 19625 15584
rect 19659 15581 19671 15615
rect 21542 15612 21548 15624
rect 21503 15584 21548 15612
rect 19613 15575 19671 15581
rect 21542 15572 21548 15584
rect 21600 15572 21606 15624
rect 23569 15615 23627 15621
rect 23569 15581 23581 15615
rect 23615 15612 23627 15615
rect 23658 15612 23664 15624
rect 23615 15584 23664 15612
rect 23615 15581 23627 15584
rect 23569 15575 23627 15581
rect 23658 15572 23664 15584
rect 23716 15572 23722 15624
rect 1104 15522 26864 15544
rect 1104 15470 10315 15522
rect 10367 15470 10379 15522
rect 10431 15470 10443 15522
rect 10495 15470 10507 15522
rect 10559 15470 19648 15522
rect 19700 15470 19712 15522
rect 19764 15470 19776 15522
rect 19828 15470 19840 15522
rect 19892 15470 26864 15522
rect 1104 15448 26864 15470
rect 14734 15368 14740 15420
rect 14792 15408 14798 15420
rect 15013 15411 15071 15417
rect 15013 15408 15025 15411
rect 14792 15380 15025 15408
rect 14792 15368 14798 15380
rect 15013 15377 15025 15380
rect 15059 15377 15071 15411
rect 15013 15371 15071 15377
rect 15381 15411 15439 15417
rect 15381 15377 15393 15411
rect 15427 15408 15439 15411
rect 15838 15408 15844 15420
rect 15427 15380 15844 15408
rect 15427 15377 15439 15380
rect 15381 15371 15439 15377
rect 15838 15368 15844 15380
rect 15896 15368 15902 15420
rect 16390 15408 16396 15420
rect 16351 15380 16396 15408
rect 16390 15368 16396 15380
rect 16448 15368 16454 15420
rect 18417 15411 18475 15417
rect 18417 15377 18429 15411
rect 18463 15408 18475 15411
rect 18598 15408 18604 15420
rect 18463 15380 18604 15408
rect 18463 15377 18475 15380
rect 18417 15371 18475 15377
rect 18598 15368 18604 15380
rect 18656 15368 18662 15420
rect 18782 15408 18788 15420
rect 18743 15380 18788 15408
rect 18782 15368 18788 15380
rect 18840 15368 18846 15420
rect 20346 15408 20352 15420
rect 20307 15380 20352 15408
rect 20346 15368 20352 15380
rect 20404 15368 20410 15420
rect 22278 15368 22284 15420
rect 22336 15408 22342 15420
rect 22557 15411 22615 15417
rect 22557 15408 22569 15411
rect 22336 15380 22569 15408
rect 22336 15368 22342 15380
rect 22557 15377 22569 15380
rect 22603 15408 22615 15411
rect 22833 15411 22891 15417
rect 22833 15408 22845 15411
rect 22603 15380 22845 15408
rect 22603 15377 22615 15380
rect 22557 15371 22615 15377
rect 22833 15377 22845 15380
rect 22879 15408 22891 15411
rect 23014 15408 23020 15420
rect 22879 15380 23020 15408
rect 22879 15377 22891 15380
rect 22833 15371 22891 15377
rect 23014 15368 23020 15380
rect 23072 15368 23078 15420
rect 24026 15368 24032 15420
rect 24084 15408 24090 15420
rect 24121 15411 24179 15417
rect 24121 15408 24133 15411
rect 24084 15380 24133 15408
rect 24084 15368 24090 15380
rect 24121 15377 24133 15380
rect 24167 15408 24179 15411
rect 24854 15408 24860 15420
rect 24167 15380 24860 15408
rect 24167 15377 24179 15380
rect 24121 15371 24179 15377
rect 24854 15368 24860 15380
rect 24912 15368 24918 15420
rect 25409 15411 25467 15417
rect 25409 15377 25421 15411
rect 25455 15408 25467 15411
rect 25590 15408 25596 15420
rect 25455 15380 25596 15408
rect 25455 15377 25467 15380
rect 25409 15371 25467 15377
rect 25590 15368 25596 15380
rect 25648 15368 25654 15420
rect 19242 15349 19248 15352
rect 19236 15340 19248 15349
rect 19203 15312 19248 15340
rect 19236 15303 19248 15312
rect 19242 15300 19248 15303
rect 19300 15300 19306 15352
rect 13906 15281 13912 15284
rect 13900 15272 13912 15281
rect 13867 15244 13912 15272
rect 13900 15235 13912 15244
rect 13906 15232 13912 15235
rect 13964 15232 13970 15284
rect 15286 15232 15292 15284
rect 15344 15272 15350 15284
rect 16298 15272 16304 15284
rect 15344 15244 16304 15272
rect 15344 15232 15350 15244
rect 16298 15232 16304 15244
rect 16356 15232 16362 15284
rect 20714 15232 20720 15284
rect 20772 15272 20778 15284
rect 21177 15275 21235 15281
rect 21177 15272 21189 15275
rect 20772 15244 21189 15272
rect 20772 15232 20778 15244
rect 21177 15241 21189 15244
rect 21223 15272 21235 15275
rect 21266 15272 21272 15284
rect 21223 15244 21272 15272
rect 21223 15241 21235 15244
rect 21177 15235 21235 15241
rect 21266 15232 21272 15244
rect 21324 15232 21330 15284
rect 21444 15275 21502 15281
rect 21444 15241 21456 15275
rect 21490 15272 21502 15275
rect 21726 15272 21732 15284
rect 21490 15244 21732 15272
rect 21490 15241 21502 15244
rect 21444 15235 21502 15241
rect 21726 15232 21732 15244
rect 21784 15232 21790 15284
rect 23474 15232 23480 15284
rect 23532 15272 23538 15284
rect 24029 15275 24087 15281
rect 24029 15272 24041 15275
rect 23532 15244 24041 15272
rect 23532 15232 23538 15244
rect 24029 15241 24041 15244
rect 24075 15241 24087 15275
rect 24029 15235 24087 15241
rect 25225 15275 25283 15281
rect 25225 15241 25237 15275
rect 25271 15272 25283 15275
rect 25866 15272 25872 15284
rect 25271 15244 25872 15272
rect 25271 15241 25283 15244
rect 25225 15235 25283 15241
rect 25866 15232 25872 15244
rect 25924 15232 25930 15284
rect 13630 15204 13636 15216
rect 13591 15176 13636 15204
rect 13630 15164 13636 15176
rect 13688 15164 13694 15216
rect 16485 15207 16543 15213
rect 16485 15173 16497 15207
rect 16531 15173 16543 15207
rect 16485 15167 16543 15173
rect 15841 15139 15899 15145
rect 15841 15105 15853 15139
rect 15887 15136 15899 15139
rect 16500 15136 16528 15167
rect 18782 15164 18788 15216
rect 18840 15204 18846 15216
rect 18969 15207 19027 15213
rect 18969 15204 18981 15207
rect 18840 15176 18981 15204
rect 18840 15164 18846 15176
rect 18969 15173 18981 15176
rect 19015 15173 19027 15207
rect 18969 15167 19027 15173
rect 23658 15164 23664 15216
rect 23716 15204 23722 15216
rect 24118 15204 24124 15216
rect 23716 15176 24124 15204
rect 23716 15164 23722 15176
rect 24118 15164 24124 15176
rect 24176 15204 24182 15216
rect 24213 15207 24271 15213
rect 24213 15204 24225 15207
rect 24176 15176 24225 15204
rect 24176 15164 24182 15176
rect 24213 15173 24225 15176
rect 24259 15173 24271 15207
rect 24213 15167 24271 15173
rect 16850 15136 16856 15148
rect 15887 15108 16856 15136
rect 15887 15105 15899 15108
rect 15841 15099 15899 15105
rect 16850 15096 16856 15108
rect 16908 15136 16914 15148
rect 16945 15139 17003 15145
rect 16945 15136 16957 15139
rect 16908 15108 16957 15136
rect 16908 15096 16914 15108
rect 16945 15105 16957 15108
rect 16991 15105 17003 15139
rect 16945 15099 17003 15105
rect 15930 15068 15936 15080
rect 15891 15040 15936 15068
rect 15930 15028 15936 15040
rect 15988 15028 15994 15080
rect 23658 15068 23664 15080
rect 23619 15040 23664 15068
rect 23658 15028 23664 15040
rect 23716 15028 23722 15080
rect 1104 14978 26864 15000
rect 1104 14926 5648 14978
rect 5700 14926 5712 14978
rect 5764 14926 5776 14978
rect 5828 14926 5840 14978
rect 5892 14926 14982 14978
rect 15034 14926 15046 14978
rect 15098 14926 15110 14978
rect 15162 14926 15174 14978
rect 15226 14926 24315 14978
rect 24367 14926 24379 14978
rect 24431 14926 24443 14978
rect 24495 14926 24507 14978
rect 24559 14926 26864 14978
rect 1104 14904 26864 14926
rect 13906 14824 13912 14876
rect 13964 14864 13970 14876
rect 14001 14867 14059 14873
rect 14001 14864 14013 14867
rect 13964 14836 14013 14864
rect 13964 14824 13970 14836
rect 14001 14833 14013 14836
rect 14047 14833 14059 14867
rect 14001 14827 14059 14833
rect 14642 14824 14648 14876
rect 14700 14864 14706 14876
rect 15105 14867 15163 14873
rect 15105 14864 15117 14867
rect 14700 14836 15117 14864
rect 14700 14824 14706 14836
rect 15105 14833 15117 14836
rect 15151 14864 15163 14867
rect 15286 14864 15292 14876
rect 15151 14836 15292 14864
rect 15151 14833 15163 14836
rect 15105 14827 15163 14833
rect 15286 14824 15292 14836
rect 15344 14824 15350 14876
rect 15470 14864 15476 14876
rect 15431 14836 15476 14864
rect 15470 14824 15476 14836
rect 15528 14824 15534 14876
rect 16025 14867 16083 14873
rect 16025 14833 16037 14867
rect 16071 14864 16083 14867
rect 16390 14864 16396 14876
rect 16071 14836 16396 14864
rect 16071 14833 16083 14836
rect 16025 14827 16083 14833
rect 16390 14824 16396 14836
rect 16448 14824 16454 14876
rect 18874 14864 18880 14876
rect 18835 14836 18880 14864
rect 18874 14824 18880 14836
rect 18932 14824 18938 14876
rect 19334 14824 19340 14876
rect 19392 14864 19398 14876
rect 19889 14867 19947 14873
rect 19889 14864 19901 14867
rect 19392 14836 19901 14864
rect 19392 14824 19398 14836
rect 19889 14833 19901 14836
rect 19935 14833 19947 14867
rect 19889 14827 19947 14833
rect 21266 14824 21272 14876
rect 21324 14864 21330 14876
rect 21361 14867 21419 14873
rect 21361 14864 21373 14867
rect 21324 14836 21373 14864
rect 21324 14824 21330 14836
rect 21361 14833 21373 14836
rect 21407 14833 21419 14867
rect 21726 14864 21732 14876
rect 21687 14836 21732 14864
rect 21361 14827 21419 14833
rect 21726 14824 21732 14836
rect 21784 14824 21790 14876
rect 23753 14867 23811 14873
rect 23753 14833 23765 14867
rect 23799 14864 23811 14867
rect 24118 14864 24124 14876
rect 23799 14836 24124 14864
rect 23799 14833 23811 14836
rect 23753 14827 23811 14833
rect 24118 14824 24124 14836
rect 24176 14824 24182 14876
rect 24854 14864 24860 14876
rect 24815 14836 24860 14864
rect 24854 14824 24860 14836
rect 24912 14824 24918 14876
rect 25498 14864 25504 14876
rect 25459 14836 25504 14864
rect 25498 14824 25504 14836
rect 25556 14824 25562 14876
rect 25866 14864 25872 14876
rect 25827 14836 25872 14864
rect 25866 14824 25872 14836
rect 25924 14824 25930 14876
rect 15746 14756 15752 14808
rect 15804 14796 15810 14808
rect 16485 14799 16543 14805
rect 16485 14796 16497 14799
rect 15804 14768 16497 14796
rect 15804 14756 15810 14768
rect 16485 14765 16497 14768
rect 16531 14796 16543 14799
rect 22465 14799 22523 14805
rect 16531 14768 16712 14796
rect 16531 14765 16543 14768
rect 16485 14759 16543 14765
rect 16684 14737 16712 14768
rect 22465 14765 22477 14799
rect 22511 14796 22523 14799
rect 23474 14796 23480 14808
rect 22511 14768 23480 14796
rect 22511 14765 22523 14768
rect 22465 14759 22523 14765
rect 23474 14756 23480 14768
rect 23532 14756 23538 14808
rect 16669 14731 16727 14737
rect 16669 14697 16681 14731
rect 16715 14697 16727 14731
rect 16669 14691 16727 14697
rect 19058 14688 19064 14740
rect 19116 14728 19122 14740
rect 19337 14731 19395 14737
rect 19337 14728 19349 14731
rect 19116 14700 19349 14728
rect 19116 14688 19122 14700
rect 19337 14697 19349 14700
rect 19383 14697 19395 14731
rect 19518 14728 19524 14740
rect 19431 14700 19524 14728
rect 19337 14691 19395 14697
rect 19518 14688 19524 14700
rect 19576 14728 19582 14740
rect 20257 14731 20315 14737
rect 20257 14728 20269 14731
rect 19576 14700 20269 14728
rect 19576 14688 19582 14700
rect 20257 14697 20269 14700
rect 20303 14697 20315 14731
rect 20714 14728 20720 14740
rect 20675 14700 20720 14728
rect 20257 14691 20315 14697
rect 20714 14688 20720 14700
rect 20772 14688 20778 14740
rect 23014 14728 23020 14740
rect 22975 14700 23020 14728
rect 23014 14688 23020 14700
rect 23072 14688 23078 14740
rect 24305 14731 24363 14737
rect 24305 14697 24317 14731
rect 24351 14728 24363 14731
rect 24670 14728 24676 14740
rect 24351 14700 24676 14728
rect 24351 14697 24363 14700
rect 24305 14691 24363 14697
rect 24670 14688 24676 14700
rect 24728 14688 24734 14740
rect 15289 14663 15347 14669
rect 15289 14629 15301 14663
rect 15335 14660 15347 14663
rect 15378 14660 15384 14672
rect 15335 14632 15384 14660
rect 15335 14629 15347 14632
rect 15289 14623 15347 14629
rect 15378 14620 15384 14632
rect 15436 14620 15442 14672
rect 22554 14620 22560 14672
rect 22612 14660 22618 14672
rect 22833 14663 22891 14669
rect 22833 14660 22845 14663
rect 22612 14632 22845 14660
rect 22612 14620 22618 14632
rect 22833 14629 22845 14632
rect 22879 14629 22891 14663
rect 22833 14623 22891 14629
rect 23658 14620 23664 14672
rect 23716 14660 23722 14672
rect 24029 14663 24087 14669
rect 24029 14660 24041 14663
rect 23716 14632 24041 14660
rect 23716 14620 23722 14632
rect 24029 14629 24041 14632
rect 24075 14660 24087 14663
rect 24578 14660 24584 14672
rect 24075 14632 24584 14660
rect 24075 14629 24087 14632
rect 24029 14623 24087 14629
rect 24578 14620 24584 14632
rect 24636 14620 24642 14672
rect 25317 14663 25375 14669
rect 25317 14660 25329 14663
rect 25148 14632 25329 14660
rect 16850 14552 16856 14604
rect 16908 14601 16914 14604
rect 16908 14595 16972 14601
rect 16908 14561 16926 14595
rect 16960 14561 16972 14595
rect 16908 14555 16972 14561
rect 16908 14552 16914 14555
rect 18138 14552 18144 14604
rect 18196 14592 18202 14604
rect 18693 14595 18751 14601
rect 18693 14592 18705 14595
rect 18196 14564 18705 14592
rect 18196 14552 18202 14564
rect 18693 14561 18705 14564
rect 18739 14592 18751 14595
rect 18782 14592 18788 14604
rect 18739 14564 18788 14592
rect 18739 14561 18751 14564
rect 18693 14555 18751 14561
rect 18782 14552 18788 14564
rect 18840 14552 18846 14604
rect 13630 14524 13636 14536
rect 13591 14496 13636 14524
rect 13630 14484 13636 14496
rect 13688 14484 13694 14536
rect 18046 14524 18052 14536
rect 18007 14496 18052 14524
rect 18046 14484 18052 14496
rect 18104 14484 18110 14536
rect 18414 14524 18420 14536
rect 18327 14496 18420 14524
rect 18414 14484 18420 14496
rect 18472 14524 18478 14536
rect 19242 14524 19248 14536
rect 18472 14496 19248 14524
rect 18472 14484 18478 14496
rect 19242 14484 19248 14496
rect 19300 14484 19306 14536
rect 20898 14524 20904 14536
rect 20859 14496 20904 14524
rect 20898 14484 20904 14496
rect 20956 14484 20962 14536
rect 22186 14484 22192 14536
rect 22244 14524 22250 14536
rect 22373 14527 22431 14533
rect 22373 14524 22385 14527
rect 22244 14496 22385 14524
rect 22244 14484 22250 14496
rect 22373 14493 22385 14496
rect 22419 14524 22431 14527
rect 22922 14524 22928 14536
rect 22419 14496 22928 14524
rect 22419 14493 22431 14496
rect 22373 14487 22431 14493
rect 22922 14484 22928 14496
rect 22980 14484 22986 14536
rect 25038 14484 25044 14536
rect 25096 14524 25102 14536
rect 25148 14533 25176 14632
rect 25317 14629 25329 14632
rect 25363 14629 25375 14663
rect 25317 14623 25375 14629
rect 25133 14527 25191 14533
rect 25133 14524 25145 14527
rect 25096 14496 25145 14524
rect 25096 14484 25102 14496
rect 25133 14493 25145 14496
rect 25179 14493 25191 14527
rect 25133 14487 25191 14493
rect 1104 14434 26864 14456
rect 1104 14382 10315 14434
rect 10367 14382 10379 14434
rect 10431 14382 10443 14434
rect 10495 14382 10507 14434
rect 10559 14382 19648 14434
rect 19700 14382 19712 14434
rect 19764 14382 19776 14434
rect 19828 14382 19840 14434
rect 19892 14382 26864 14434
rect 1104 14360 26864 14382
rect 13538 14280 13544 14332
rect 13596 14320 13602 14332
rect 13633 14323 13691 14329
rect 13633 14320 13645 14323
rect 13596 14292 13645 14320
rect 13596 14280 13602 14292
rect 13633 14289 13645 14292
rect 13679 14289 13691 14323
rect 13633 14283 13691 14289
rect 16850 14280 16856 14332
rect 16908 14320 16914 14332
rect 16945 14323 17003 14329
rect 16945 14320 16957 14323
rect 16908 14292 16957 14320
rect 16908 14280 16914 14292
rect 16945 14289 16957 14292
rect 16991 14289 17003 14323
rect 16945 14283 17003 14289
rect 19334 14280 19340 14332
rect 19392 14320 19398 14332
rect 19705 14323 19763 14329
rect 19705 14320 19717 14323
rect 19392 14292 19717 14320
rect 19392 14280 19398 14292
rect 19705 14289 19717 14292
rect 19751 14289 19763 14323
rect 22554 14320 22560 14332
rect 22515 14292 22560 14320
rect 19705 14283 19763 14289
rect 22554 14280 22560 14292
rect 22612 14280 22618 14332
rect 22925 14323 22983 14329
rect 22925 14289 22937 14323
rect 22971 14320 22983 14323
rect 23014 14320 23020 14332
rect 22971 14292 23020 14320
rect 22971 14289 22983 14292
rect 22925 14283 22983 14289
rect 23014 14280 23020 14292
rect 23072 14280 23078 14332
rect 23474 14320 23480 14332
rect 23435 14292 23480 14320
rect 23474 14280 23480 14292
rect 23532 14280 23538 14332
rect 24578 14320 24584 14332
rect 24539 14292 24584 14320
rect 24578 14280 24584 14292
rect 24636 14280 24642 14332
rect 25130 14280 25136 14332
rect 25188 14320 25194 14332
rect 25317 14323 25375 14329
rect 25317 14320 25329 14323
rect 25188 14292 25329 14320
rect 25188 14280 25194 14292
rect 25317 14289 25329 14292
rect 25363 14289 25375 14323
rect 25317 14283 25375 14289
rect 15746 14212 15752 14264
rect 15804 14212 15810 14264
rect 21082 14252 21088 14264
rect 21043 14224 21088 14252
rect 21082 14212 21088 14224
rect 21140 14212 21146 14264
rect 24121 14255 24179 14261
rect 24121 14221 24133 14255
rect 24167 14252 24179 14255
rect 25038 14252 25044 14264
rect 24167 14224 25044 14252
rect 24167 14221 24179 14224
rect 24121 14215 24179 14221
rect 25038 14212 25044 14224
rect 25096 14212 25102 14264
rect 13446 14184 13452 14196
rect 13407 14156 13452 14184
rect 13446 14144 13452 14156
rect 13504 14144 13510 14196
rect 15565 14187 15623 14193
rect 15565 14153 15577 14187
rect 15611 14184 15623 14187
rect 15764 14184 15792 14212
rect 15611 14156 15792 14184
rect 15832 14187 15890 14193
rect 15611 14153 15623 14156
rect 15565 14147 15623 14153
rect 15832 14153 15844 14187
rect 15878 14184 15890 14187
rect 16390 14184 16396 14196
rect 15878 14156 16396 14184
rect 15878 14153 15890 14156
rect 15832 14147 15890 14153
rect 16390 14144 16396 14156
rect 16448 14144 16454 14196
rect 18046 14144 18052 14196
rect 18104 14184 18110 14196
rect 18592 14187 18650 14193
rect 18592 14184 18604 14187
rect 18104 14156 18604 14184
rect 18104 14144 18110 14156
rect 18592 14153 18604 14156
rect 18638 14184 18650 14187
rect 19518 14184 19524 14196
rect 18638 14156 19524 14184
rect 18638 14153 18650 14156
rect 18592 14147 18650 14153
rect 19518 14144 19524 14156
rect 19576 14144 19582 14196
rect 20806 14184 20812 14196
rect 20767 14156 20812 14184
rect 20806 14144 20812 14156
rect 20864 14144 20870 14196
rect 23658 14144 23664 14196
rect 23716 14184 23722 14196
rect 23845 14187 23903 14193
rect 23845 14184 23857 14187
rect 23716 14156 23857 14184
rect 23716 14144 23722 14156
rect 23845 14153 23857 14156
rect 23891 14153 23903 14187
rect 23845 14147 23903 14153
rect 25133 14187 25191 14193
rect 25133 14153 25145 14187
rect 25179 14184 25191 14187
rect 25590 14184 25596 14196
rect 25179 14156 25596 14184
rect 25179 14153 25191 14156
rect 25133 14147 25191 14153
rect 25590 14144 25596 14156
rect 25648 14144 25654 14196
rect 18138 14076 18144 14128
rect 18196 14116 18202 14128
rect 18325 14119 18383 14125
rect 18325 14116 18337 14119
rect 18196 14088 18337 14116
rect 18196 14076 18202 14088
rect 18325 14085 18337 14088
rect 18371 14085 18383 14119
rect 18325 14079 18383 14085
rect 15378 13980 15384 13992
rect 15339 13952 15384 13980
rect 15378 13940 15384 13952
rect 15436 13940 15442 13992
rect 1104 13890 26864 13912
rect 1104 13838 5648 13890
rect 5700 13838 5712 13890
rect 5764 13838 5776 13890
rect 5828 13838 5840 13890
rect 5892 13838 14982 13890
rect 15034 13838 15046 13890
rect 15098 13838 15110 13890
rect 15162 13838 15174 13890
rect 15226 13838 24315 13890
rect 24367 13838 24379 13890
rect 24431 13838 24443 13890
rect 24495 13838 24507 13890
rect 24559 13838 26864 13890
rect 1104 13816 26864 13838
rect 13446 13776 13452 13788
rect 13407 13748 13452 13776
rect 13446 13736 13452 13748
rect 13504 13736 13510 13788
rect 15746 13736 15752 13788
rect 15804 13776 15810 13788
rect 15930 13776 15936 13788
rect 15804 13748 15936 13776
rect 15804 13736 15810 13748
rect 15930 13736 15936 13748
rect 15988 13776 15994 13788
rect 16025 13779 16083 13785
rect 16025 13776 16037 13779
rect 15988 13748 16037 13776
rect 15988 13736 15994 13748
rect 16025 13745 16037 13748
rect 16071 13745 16083 13779
rect 16390 13776 16396 13788
rect 16351 13748 16396 13776
rect 16025 13739 16083 13745
rect 16390 13736 16396 13748
rect 16448 13736 16454 13788
rect 16853 13779 16911 13785
rect 16853 13745 16865 13779
rect 16899 13776 16911 13779
rect 16942 13776 16948 13788
rect 16899 13748 16948 13776
rect 16899 13745 16911 13748
rect 16853 13739 16911 13745
rect 16942 13736 16948 13748
rect 17000 13736 17006 13788
rect 17681 13779 17739 13785
rect 17681 13745 17693 13779
rect 17727 13776 17739 13779
rect 18046 13776 18052 13788
rect 17727 13748 18052 13776
rect 17727 13745 17739 13748
rect 17681 13739 17739 13745
rect 18046 13736 18052 13748
rect 18104 13736 18110 13788
rect 18509 13779 18567 13785
rect 18509 13745 18521 13779
rect 18555 13776 18567 13779
rect 18966 13776 18972 13788
rect 18555 13748 18972 13776
rect 18555 13745 18567 13748
rect 18509 13739 18567 13745
rect 18966 13736 18972 13748
rect 19024 13736 19030 13788
rect 19518 13776 19524 13788
rect 19479 13748 19524 13776
rect 19518 13736 19524 13748
rect 19576 13736 19582 13788
rect 20254 13776 20260 13788
rect 20215 13748 20260 13776
rect 20254 13736 20260 13748
rect 20312 13776 20318 13788
rect 20312 13748 21496 13776
rect 20312 13736 20318 13748
rect 12989 13643 13047 13649
rect 12989 13609 13001 13643
rect 13035 13640 13047 13643
rect 13464 13640 13492 13736
rect 17954 13708 17960 13720
rect 17915 13680 17960 13708
rect 17954 13668 17960 13680
rect 18012 13668 18018 13720
rect 13035 13612 13492 13640
rect 13035 13609 13047 13612
rect 12989 13603 13047 13609
rect 15378 13600 15384 13652
rect 15436 13640 15442 13652
rect 15473 13643 15531 13649
rect 15473 13640 15485 13643
rect 15436 13612 15485 13640
rect 15436 13600 15442 13612
rect 15473 13609 15485 13612
rect 15519 13609 15531 13643
rect 17972 13640 18000 13668
rect 18969 13643 19027 13649
rect 18969 13640 18981 13643
rect 17972 13612 18981 13640
rect 15473 13603 15531 13609
rect 18969 13609 18981 13612
rect 19015 13609 19027 13643
rect 18969 13603 19027 13609
rect 19153 13643 19211 13649
rect 19153 13609 19165 13643
rect 19199 13640 19211 13643
rect 19536 13640 19564 13736
rect 19981 13711 20039 13717
rect 19981 13677 19993 13711
rect 20027 13708 20039 13711
rect 20806 13708 20812 13720
rect 20027 13680 20812 13708
rect 20027 13677 20039 13680
rect 19981 13671 20039 13677
rect 20806 13668 20812 13680
rect 20864 13708 20870 13720
rect 20901 13711 20959 13717
rect 20901 13708 20913 13711
rect 20864 13680 20913 13708
rect 20864 13668 20870 13680
rect 20901 13677 20913 13680
rect 20947 13677 20959 13711
rect 20901 13671 20959 13677
rect 21468 13649 21496 13748
rect 23658 13736 23664 13788
rect 23716 13776 23722 13788
rect 23845 13779 23903 13785
rect 23845 13776 23857 13779
rect 23716 13748 23857 13776
rect 23716 13736 23722 13748
rect 23845 13745 23857 13748
rect 23891 13745 23903 13779
rect 23845 13739 23903 13745
rect 23934 13736 23940 13788
rect 23992 13776 23998 13788
rect 24765 13779 24823 13785
rect 24765 13776 24777 13779
rect 23992 13748 24777 13776
rect 23992 13736 23998 13748
rect 24765 13745 24777 13748
rect 24811 13745 24823 13779
rect 25590 13776 25596 13788
rect 25551 13748 25596 13776
rect 24765 13739 24823 13745
rect 25590 13736 25596 13748
rect 25648 13736 25654 13788
rect 19199 13612 19564 13640
rect 21453 13643 21511 13649
rect 19199 13609 19211 13612
rect 19153 13603 19211 13609
rect 21453 13609 21465 13643
rect 21499 13640 21511 13643
rect 22094 13640 22100 13652
rect 21499 13612 22100 13640
rect 21499 13609 21511 13612
rect 21453 13603 21511 13609
rect 22094 13600 22100 13612
rect 22152 13600 22158 13652
rect 25222 13640 25228 13652
rect 25183 13612 25228 13640
rect 25222 13600 25228 13612
rect 25280 13600 25286 13652
rect 12713 13575 12771 13581
rect 12713 13541 12725 13575
rect 12759 13541 12771 13575
rect 12713 13535 12771 13541
rect 15105 13575 15163 13581
rect 15105 13541 15117 13575
rect 15151 13572 15163 13575
rect 15286 13572 15292 13584
rect 15151 13544 15292 13572
rect 15151 13541 15163 13544
rect 15105 13535 15163 13541
rect 12621 13439 12679 13445
rect 12621 13405 12633 13439
rect 12667 13436 12679 13439
rect 12728 13436 12756 13535
rect 15286 13532 15292 13544
rect 15344 13532 15350 13584
rect 16669 13575 16727 13581
rect 16669 13541 16681 13575
rect 16715 13572 16727 13575
rect 16942 13572 16948 13584
rect 16715 13544 16948 13572
rect 16715 13541 16727 13544
rect 16669 13535 16727 13541
rect 16942 13532 16948 13544
rect 17000 13572 17006 13584
rect 17221 13575 17279 13581
rect 17221 13572 17233 13575
rect 17000 13544 17233 13572
rect 17000 13532 17006 13544
rect 17221 13541 17233 13544
rect 17267 13541 17279 13575
rect 17221 13535 17279 13541
rect 18138 13532 18144 13584
rect 18196 13572 18202 13584
rect 18325 13575 18383 13581
rect 18325 13572 18337 13575
rect 18196 13544 18337 13572
rect 18196 13532 18202 13544
rect 18325 13541 18337 13544
rect 18371 13541 18383 13575
rect 18325 13535 18383 13541
rect 20806 13532 20812 13584
rect 20864 13572 20870 13584
rect 21361 13575 21419 13581
rect 21361 13572 21373 13575
rect 20864 13544 21373 13572
rect 20864 13532 20870 13544
rect 21361 13541 21373 13544
rect 21407 13572 21419 13575
rect 21913 13575 21971 13581
rect 21913 13572 21925 13575
rect 21407 13544 21925 13572
rect 21407 13541 21419 13544
rect 21361 13535 21419 13541
rect 21913 13541 21925 13544
rect 21959 13541 21971 13575
rect 21913 13535 21971 13541
rect 24581 13575 24639 13581
rect 24581 13541 24593 13575
rect 24627 13572 24639 13575
rect 25240 13572 25268 13600
rect 24627 13544 25268 13572
rect 24627 13541 24639 13544
rect 24581 13535 24639 13541
rect 18874 13504 18880 13516
rect 18835 13476 18880 13504
rect 18874 13464 18880 13476
rect 18932 13464 18938 13516
rect 20717 13507 20775 13513
rect 20717 13473 20729 13507
rect 20763 13504 20775 13507
rect 21269 13507 21327 13513
rect 21269 13504 21281 13507
rect 20763 13476 21281 13504
rect 20763 13473 20775 13476
rect 20717 13467 20775 13473
rect 21269 13473 21281 13476
rect 21315 13504 21327 13507
rect 21818 13504 21824 13516
rect 21315 13476 21824 13504
rect 21315 13473 21327 13476
rect 21269 13467 21327 13473
rect 21818 13464 21824 13476
rect 21876 13464 21882 13516
rect 13170 13436 13176 13448
rect 12667 13408 13176 13436
rect 12667 13405 12679 13408
rect 12621 13399 12679 13405
rect 13170 13396 13176 13408
rect 13228 13396 13234 13448
rect 1104 13346 26864 13368
rect 1104 13294 10315 13346
rect 10367 13294 10379 13346
rect 10431 13294 10443 13346
rect 10495 13294 10507 13346
rect 10559 13294 19648 13346
rect 19700 13294 19712 13346
rect 19764 13294 19776 13346
rect 19828 13294 19840 13346
rect 19892 13294 26864 13346
rect 1104 13272 26864 13294
rect 18785 13235 18843 13241
rect 18785 13201 18797 13235
rect 18831 13232 18843 13235
rect 18874 13232 18880 13244
rect 18831 13204 18880 13232
rect 18831 13201 18843 13204
rect 18785 13195 18843 13201
rect 18874 13192 18880 13204
rect 18932 13192 18938 13244
rect 21818 13232 21824 13244
rect 21779 13204 21824 13232
rect 21818 13192 21824 13204
rect 21876 13192 21882 13244
rect 23842 13192 23848 13244
rect 23900 13232 23906 13244
rect 24765 13235 24823 13241
rect 24765 13232 24777 13235
rect 23900 13204 24777 13232
rect 23900 13192 23906 13204
rect 24765 13201 24777 13204
rect 24811 13201 24823 13235
rect 24765 13195 24823 13201
rect 16942 13164 16948 13176
rect 16903 13136 16948 13164
rect 16942 13124 16948 13136
rect 17000 13124 17006 13176
rect 21266 13164 21272 13176
rect 19628 13136 21272 13164
rect 19628 13108 19656 13136
rect 21266 13124 21272 13136
rect 21324 13124 21330 13176
rect 16666 13096 16672 13108
rect 16627 13068 16672 13096
rect 16666 13056 16672 13068
rect 16724 13056 16730 13108
rect 19610 13096 19616 13108
rect 19523 13068 19616 13096
rect 19610 13056 19616 13068
rect 19668 13056 19674 13108
rect 19886 13105 19892 13108
rect 19880 13096 19892 13105
rect 19847 13068 19892 13096
rect 19880 13059 19892 13068
rect 19886 13056 19892 13059
rect 19944 13056 19950 13108
rect 24581 13099 24639 13105
rect 24581 13065 24593 13099
rect 24627 13096 24639 13099
rect 25038 13096 25044 13108
rect 24627 13068 25044 13096
rect 24627 13065 24639 13068
rect 24581 13059 24639 13065
rect 25038 13056 25044 13068
rect 25096 13056 25102 13108
rect 12713 13031 12771 13037
rect 12713 12997 12725 13031
rect 12759 13028 12771 13031
rect 12986 13028 12992 13040
rect 12759 13000 12992 13028
rect 12759 12997 12771 13000
rect 12713 12991 12771 12997
rect 12986 12988 12992 13000
rect 13044 12988 13050 13040
rect 18046 12988 18052 13040
rect 18104 13028 18110 13040
rect 18233 13031 18291 13037
rect 18233 13028 18245 13031
rect 18104 13000 18245 13028
rect 18104 12988 18110 13000
rect 18233 12997 18245 13000
rect 18279 12997 18291 13031
rect 18233 12991 18291 12997
rect 13262 12892 13268 12904
rect 13223 12864 13268 12892
rect 13262 12852 13268 12864
rect 13320 12852 13326 12904
rect 15381 12895 15439 12901
rect 15381 12861 15393 12895
rect 15427 12892 15439 12895
rect 15838 12892 15844 12904
rect 15427 12864 15844 12892
rect 15427 12861 15439 12864
rect 15381 12855 15439 12861
rect 15838 12852 15844 12864
rect 15896 12852 15902 12904
rect 20993 12895 21051 12901
rect 20993 12861 21005 12895
rect 21039 12892 21051 12895
rect 21358 12892 21364 12904
rect 21039 12864 21364 12892
rect 21039 12861 21051 12864
rect 20993 12855 21051 12861
rect 21358 12852 21364 12864
rect 21416 12852 21422 12904
rect 1104 12802 26864 12824
rect 1104 12750 5648 12802
rect 5700 12750 5712 12802
rect 5764 12750 5776 12802
rect 5828 12750 5840 12802
rect 5892 12750 14982 12802
rect 15034 12750 15046 12802
rect 15098 12750 15110 12802
rect 15162 12750 15174 12802
rect 15226 12750 24315 12802
rect 24367 12750 24379 12802
rect 24431 12750 24443 12802
rect 24495 12750 24507 12802
rect 24559 12750 26864 12802
rect 1104 12728 26864 12750
rect 12986 12688 12992 12700
rect 12947 12660 12992 12688
rect 12986 12648 12992 12660
rect 13044 12648 13050 12700
rect 13170 12688 13176 12700
rect 13131 12660 13176 12688
rect 13170 12648 13176 12660
rect 13228 12648 13234 12700
rect 15286 12688 15292 12700
rect 15247 12660 15292 12688
rect 15286 12648 15292 12660
rect 15344 12648 15350 12700
rect 18046 12688 18052 12700
rect 18007 12660 18052 12688
rect 18046 12648 18052 12660
rect 18104 12648 18110 12700
rect 19610 12688 19616 12700
rect 19571 12660 19616 12688
rect 19610 12648 19616 12660
rect 19668 12688 19674 12700
rect 20625 12691 20683 12697
rect 20625 12688 20637 12691
rect 19668 12660 20637 12688
rect 19668 12648 19674 12660
rect 20625 12657 20637 12660
rect 20671 12657 20683 12691
rect 20625 12651 20683 12657
rect 13004 12484 13032 12648
rect 16666 12580 16672 12632
rect 16724 12620 16730 12632
rect 16761 12623 16819 12629
rect 16761 12620 16773 12623
rect 16724 12592 16773 12620
rect 16724 12580 16730 12592
rect 16761 12589 16773 12592
rect 16807 12620 16819 12623
rect 18141 12623 18199 12629
rect 18141 12620 18153 12623
rect 16807 12592 18153 12620
rect 16807 12589 16819 12592
rect 16761 12583 16819 12589
rect 18141 12589 18153 12592
rect 18187 12589 18199 12623
rect 18141 12583 18199 12589
rect 13262 12512 13268 12564
rect 13320 12552 13326 12564
rect 13725 12555 13783 12561
rect 13725 12552 13737 12555
rect 13320 12524 13737 12552
rect 13320 12512 13326 12524
rect 13725 12521 13737 12524
rect 13771 12521 13783 12555
rect 15838 12552 15844 12564
rect 15799 12524 15844 12552
rect 13725 12515 13783 12521
rect 15838 12512 15844 12524
rect 15896 12552 15902 12564
rect 16482 12552 16488 12564
rect 15896 12524 16488 12552
rect 15896 12512 15902 12524
rect 16482 12512 16488 12524
rect 16540 12512 16546 12564
rect 17313 12555 17371 12561
rect 17313 12521 17325 12555
rect 17359 12552 17371 12555
rect 18598 12552 18604 12564
rect 17359 12524 18604 12552
rect 17359 12521 17371 12524
rect 17313 12515 17371 12521
rect 18598 12512 18604 12524
rect 18656 12512 18662 12564
rect 18693 12555 18751 12561
rect 18693 12521 18705 12555
rect 18739 12521 18751 12555
rect 20640 12552 20668 12651
rect 22094 12648 22100 12700
rect 22152 12688 22158 12700
rect 22281 12691 22339 12697
rect 22281 12688 22293 12691
rect 22152 12660 22293 12688
rect 22152 12648 22158 12660
rect 22281 12657 22293 12660
rect 22327 12657 22339 12691
rect 24210 12688 24216 12700
rect 24171 12660 24216 12688
rect 22281 12651 22339 12657
rect 24210 12648 24216 12660
rect 24268 12648 24274 12700
rect 25038 12688 25044 12700
rect 24999 12660 25044 12688
rect 25038 12648 25044 12660
rect 25096 12648 25102 12700
rect 20901 12555 20959 12561
rect 20901 12552 20913 12555
rect 20640 12524 20913 12552
rect 18693 12515 18751 12521
rect 20901 12521 20913 12524
rect 20947 12521 20959 12555
rect 24670 12552 24676 12564
rect 20901 12515 20959 12521
rect 24044 12524 24676 12552
rect 13541 12487 13599 12493
rect 13541 12484 13553 12487
rect 13004 12456 13553 12484
rect 13541 12453 13553 12456
rect 13587 12453 13599 12487
rect 13541 12447 13599 12453
rect 18046 12444 18052 12496
rect 18104 12484 18110 12496
rect 18509 12487 18567 12493
rect 18509 12484 18521 12487
rect 18104 12456 18521 12484
rect 18104 12444 18110 12456
rect 18509 12453 18521 12456
rect 18555 12453 18567 12487
rect 18708 12484 18736 12515
rect 19518 12484 19524 12496
rect 18509 12447 18567 12453
rect 18616 12456 19524 12484
rect 12713 12419 12771 12425
rect 12713 12385 12725 12419
rect 12759 12416 12771 12419
rect 13078 12416 13084 12428
rect 12759 12388 13084 12416
rect 12759 12385 12771 12388
rect 12713 12379 12771 12385
rect 13078 12376 13084 12388
rect 13136 12416 13142 12428
rect 13633 12419 13691 12425
rect 13633 12416 13645 12419
rect 13136 12388 13645 12416
rect 13136 12376 13142 12388
rect 13633 12385 13645 12388
rect 13679 12385 13691 12419
rect 13633 12379 13691 12385
rect 15105 12419 15163 12425
rect 15105 12385 15117 12419
rect 15151 12416 15163 12419
rect 15378 12416 15384 12428
rect 15151 12388 15384 12416
rect 15151 12385 15163 12388
rect 15105 12379 15163 12385
rect 15378 12376 15384 12388
rect 15436 12416 15442 12428
rect 15657 12419 15715 12425
rect 15657 12416 15669 12419
rect 15436 12388 15669 12416
rect 15436 12376 15442 12388
rect 15657 12385 15669 12388
rect 15703 12385 15715 12419
rect 15657 12379 15715 12385
rect 14737 12351 14795 12357
rect 14737 12317 14749 12351
rect 14783 12348 14795 12351
rect 15562 12348 15568 12360
rect 14783 12320 15568 12348
rect 14783 12317 14795 12320
rect 14737 12311 14795 12317
rect 15562 12308 15568 12320
rect 15620 12348 15626 12360
rect 15749 12351 15807 12357
rect 15749 12348 15761 12351
rect 15620 12320 15761 12348
rect 15620 12308 15626 12320
rect 15749 12317 15761 12320
rect 15795 12317 15807 12351
rect 15749 12311 15807 12317
rect 17681 12351 17739 12357
rect 17681 12317 17693 12351
rect 17727 12348 17739 12351
rect 18616 12348 18644 12456
rect 19518 12444 19524 12456
rect 19576 12484 19582 12496
rect 19886 12484 19892 12496
rect 19576 12456 19892 12484
rect 19576 12444 19582 12456
rect 19886 12444 19892 12456
rect 19944 12484 19950 12496
rect 24044 12493 24072 12524
rect 24670 12512 24676 12524
rect 24728 12512 24734 12564
rect 19981 12487 20039 12493
rect 19981 12484 19993 12487
rect 19944 12456 19993 12484
rect 19944 12444 19950 12456
rect 19981 12453 19993 12456
rect 20027 12453 20039 12487
rect 19981 12447 20039 12453
rect 24029 12487 24087 12493
rect 24029 12453 24041 12487
rect 24075 12453 24087 12487
rect 24029 12447 24087 12453
rect 21168 12419 21226 12425
rect 21168 12385 21180 12419
rect 21214 12416 21226 12419
rect 21358 12416 21364 12428
rect 21214 12388 21364 12416
rect 21214 12385 21226 12388
rect 21168 12379 21226 12385
rect 21358 12376 21364 12388
rect 21416 12376 21422 12428
rect 17727 12320 18644 12348
rect 17727 12317 17739 12320
rect 17681 12311 17739 12317
rect 1104 12258 26864 12280
rect 1104 12206 10315 12258
rect 10367 12206 10379 12258
rect 10431 12206 10443 12258
rect 10495 12206 10507 12258
rect 10559 12206 19648 12258
rect 19700 12206 19712 12258
rect 19764 12206 19776 12258
rect 19828 12206 19840 12258
rect 19892 12206 26864 12258
rect 1104 12184 26864 12206
rect 16482 12104 16488 12156
rect 16540 12144 16546 12156
rect 16577 12147 16635 12153
rect 16577 12144 16589 12147
rect 16540 12116 16589 12144
rect 16540 12104 16546 12116
rect 16577 12113 16589 12116
rect 16623 12144 16635 12147
rect 16758 12144 16764 12156
rect 16623 12116 16764 12144
rect 16623 12113 16635 12116
rect 16577 12107 16635 12113
rect 16758 12104 16764 12116
rect 16816 12104 16822 12156
rect 19518 12144 19524 12156
rect 19479 12116 19524 12144
rect 19518 12104 19524 12116
rect 19576 12104 19582 12156
rect 20806 12144 20812 12156
rect 20767 12116 20812 12144
rect 20806 12104 20812 12116
rect 20864 12104 20870 12156
rect 24026 12104 24032 12156
rect 24084 12144 24090 12156
rect 24765 12147 24823 12153
rect 24765 12144 24777 12147
rect 24084 12116 24777 12144
rect 24084 12104 24090 12116
rect 24765 12113 24777 12116
rect 24811 12113 24823 12147
rect 24765 12107 24823 12113
rect 13262 12085 13268 12088
rect 13256 12076 13268 12085
rect 13223 12048 13268 12076
rect 13256 12039 13268 12048
rect 13262 12036 13268 12039
rect 13320 12036 13326 12088
rect 13630 12036 13636 12088
rect 13688 12076 13694 12088
rect 15930 12076 15936 12088
rect 13688 12048 15936 12076
rect 13688 12036 13694 12048
rect 12526 11968 12532 12020
rect 12584 12008 12590 12020
rect 12989 12011 13047 12017
rect 12989 12008 13001 12011
rect 12584 11980 13001 12008
rect 12584 11968 12590 11980
rect 12989 11977 13001 11980
rect 13035 12008 13047 12011
rect 13648 12008 13676 12036
rect 15212 12017 15240 12048
rect 15930 12036 15936 12048
rect 15988 12036 15994 12088
rect 13035 11980 13676 12008
rect 15197 12011 15255 12017
rect 13035 11977 13047 11980
rect 12989 11971 13047 11977
rect 15197 11977 15209 12011
rect 15243 11977 15255 12011
rect 15197 11971 15255 11977
rect 15286 11968 15292 12020
rect 15344 12008 15350 12020
rect 15453 12011 15511 12017
rect 15453 12008 15465 12011
rect 15344 11980 15465 12008
rect 15344 11968 15350 11980
rect 15453 11977 15465 11980
rect 15499 11977 15511 12011
rect 15453 11971 15511 11977
rect 18046 11968 18052 12020
rect 18104 12008 18110 12020
rect 18397 12011 18455 12017
rect 18397 12008 18409 12011
rect 18104 11980 18409 12008
rect 18104 11968 18110 11980
rect 18397 11977 18409 11980
rect 18443 11977 18455 12011
rect 21174 12008 21180 12020
rect 21135 11980 21180 12008
rect 18397 11971 18455 11977
rect 21174 11968 21180 11980
rect 21232 11968 21238 12020
rect 21269 12011 21327 12017
rect 21269 11977 21281 12011
rect 21315 12008 21327 12011
rect 21450 12008 21456 12020
rect 21315 11980 21456 12008
rect 21315 11977 21327 11980
rect 21269 11971 21327 11977
rect 21450 11968 21456 11980
rect 21508 11968 21514 12020
rect 24578 12008 24584 12020
rect 24539 11980 24584 12008
rect 24578 11968 24584 11980
rect 24636 11968 24642 12020
rect 18138 11940 18144 11952
rect 18099 11912 18144 11940
rect 18138 11900 18144 11912
rect 18196 11900 18202 11952
rect 21358 11940 21364 11952
rect 21319 11912 21364 11940
rect 21358 11900 21364 11912
rect 21416 11900 21422 11952
rect 14366 11804 14372 11816
rect 14327 11776 14372 11804
rect 14366 11764 14372 11776
rect 14424 11764 14430 11816
rect 1104 11714 26864 11736
rect 1104 11662 5648 11714
rect 5700 11662 5712 11714
rect 5764 11662 5776 11714
rect 5828 11662 5840 11714
rect 5892 11662 14982 11714
rect 15034 11662 15046 11714
rect 15098 11662 15110 11714
rect 15162 11662 15174 11714
rect 15226 11662 24315 11714
rect 24367 11662 24379 11714
rect 24431 11662 24443 11714
rect 24495 11662 24507 11714
rect 24559 11662 26864 11714
rect 1104 11640 26864 11662
rect 13262 11560 13268 11612
rect 13320 11600 13326 11612
rect 13909 11603 13967 11609
rect 13909 11600 13921 11603
rect 13320 11572 13921 11600
rect 13320 11560 13326 11572
rect 13909 11569 13921 11572
rect 13955 11600 13967 11603
rect 14185 11603 14243 11609
rect 14185 11600 14197 11603
rect 13955 11572 14197 11600
rect 13955 11569 13967 11572
rect 13909 11563 13967 11569
rect 14185 11569 14197 11572
rect 14231 11569 14243 11603
rect 14185 11563 14243 11569
rect 14366 11560 14372 11612
rect 14424 11600 14430 11612
rect 15013 11603 15071 11609
rect 15013 11600 15025 11603
rect 14424 11572 15025 11600
rect 14424 11560 14430 11572
rect 15013 11569 15025 11572
rect 15059 11600 15071 11603
rect 15286 11600 15292 11612
rect 15059 11572 15292 11600
rect 15059 11569 15071 11572
rect 15013 11563 15071 11569
rect 15286 11560 15292 11572
rect 15344 11560 15350 11612
rect 15930 11600 15936 11612
rect 15843 11572 15936 11600
rect 15930 11560 15936 11572
rect 15988 11600 15994 11612
rect 16577 11603 16635 11609
rect 16577 11600 16589 11603
rect 15988 11572 16589 11600
rect 15988 11560 15994 11572
rect 16577 11569 16589 11572
rect 16623 11600 16635 11603
rect 18138 11600 18144 11612
rect 16623 11572 18144 11600
rect 16623 11569 16635 11572
rect 16577 11563 16635 11569
rect 12526 11464 12532 11476
rect 12487 11436 12532 11464
rect 12526 11424 12532 11436
rect 12584 11424 12590 11476
rect 15378 11464 15384 11476
rect 15339 11436 15384 11464
rect 15378 11424 15384 11436
rect 15436 11424 15442 11476
rect 16684 11473 16712 11572
rect 18138 11560 18144 11572
rect 18196 11600 18202 11612
rect 18325 11603 18383 11609
rect 18325 11600 18337 11603
rect 18196 11572 18337 11600
rect 18196 11560 18202 11572
rect 18325 11569 18337 11572
rect 18371 11569 18383 11603
rect 18325 11563 18383 11569
rect 18598 11560 18604 11612
rect 18656 11600 18662 11612
rect 18877 11603 18935 11609
rect 18877 11600 18889 11603
rect 18656 11572 18889 11600
rect 18656 11560 18662 11572
rect 18877 11569 18889 11572
rect 18923 11569 18935 11603
rect 18877 11563 18935 11569
rect 20717 11603 20775 11609
rect 20717 11569 20729 11603
rect 20763 11600 20775 11603
rect 21358 11600 21364 11612
rect 20763 11572 21364 11600
rect 20763 11569 20775 11572
rect 20717 11563 20775 11569
rect 21358 11560 21364 11572
rect 21416 11560 21422 11612
rect 21450 11560 21456 11612
rect 21508 11600 21514 11612
rect 24670 11600 24676 11612
rect 21508 11572 21553 11600
rect 24631 11572 24676 11600
rect 21508 11560 21514 11572
rect 24670 11560 24676 11572
rect 24728 11560 24734 11612
rect 16669 11467 16727 11473
rect 16669 11433 16681 11467
rect 16715 11433 16727 11467
rect 19426 11464 19432 11476
rect 19387 11436 19432 11464
rect 16669 11427 16727 11433
rect 19426 11424 19432 11436
rect 19484 11424 19490 11476
rect 10042 11356 10048 11408
rect 10100 11396 10106 11408
rect 10321 11399 10379 11405
rect 10321 11396 10333 11399
rect 10100 11368 10333 11396
rect 10100 11356 10106 11368
rect 10321 11365 10333 11368
rect 10367 11396 10379 11399
rect 11977 11399 12035 11405
rect 11977 11396 11989 11399
rect 10367 11368 11989 11396
rect 10367 11365 10379 11368
rect 10321 11359 10379 11365
rect 11977 11365 11989 11368
rect 12023 11396 12035 11399
rect 12345 11399 12403 11405
rect 12345 11396 12357 11399
rect 12023 11368 12357 11396
rect 12023 11365 12035 11368
rect 11977 11359 12035 11365
rect 12345 11365 12357 11368
rect 12391 11396 12403 11399
rect 12544 11396 12572 11424
rect 12391 11368 12572 11396
rect 12391 11365 12403 11368
rect 12345 11359 12403 11365
rect 16758 11356 16764 11408
rect 16816 11396 16822 11408
rect 16925 11399 16983 11405
rect 16925 11396 16937 11399
rect 16816 11368 16937 11396
rect 16816 11356 16822 11368
rect 16925 11365 16937 11368
rect 16971 11365 16983 11399
rect 16925 11359 16983 11365
rect 18966 11356 18972 11408
rect 19024 11396 19030 11408
rect 19242 11396 19248 11408
rect 19024 11368 19248 11396
rect 19024 11356 19030 11368
rect 19242 11356 19248 11368
rect 19300 11396 19306 11408
rect 19337 11399 19395 11405
rect 19337 11396 19349 11399
rect 19300 11368 19349 11396
rect 19300 11356 19306 11368
rect 19337 11365 19349 11368
rect 19383 11365 19395 11399
rect 21174 11396 21180 11408
rect 21135 11368 21180 11396
rect 19337 11359 19395 11365
rect 21174 11356 21180 11368
rect 21232 11356 21238 11408
rect 10134 11328 10140 11340
rect 10095 11300 10140 11328
rect 10134 11288 10140 11300
rect 10192 11328 10198 11340
rect 12802 11337 12808 11340
rect 10566 11331 10624 11337
rect 10566 11328 10578 11331
rect 10192 11300 10578 11328
rect 10192 11288 10198 11300
rect 10566 11297 10578 11300
rect 10612 11297 10624 11331
rect 12796 11328 12808 11337
rect 10566 11291 10624 11297
rect 11716 11300 12808 11328
rect 11716 11269 11744 11300
rect 12796 11291 12808 11300
rect 12802 11288 12808 11291
rect 12860 11288 12866 11340
rect 11701 11263 11759 11269
rect 11701 11229 11713 11263
rect 11747 11229 11759 11263
rect 18046 11260 18052 11272
rect 18007 11232 18052 11260
rect 11701 11223 11759 11229
rect 18046 11220 18052 11232
rect 18104 11220 18110 11272
rect 18785 11263 18843 11269
rect 18785 11229 18797 11263
rect 18831 11260 18843 11263
rect 19242 11260 19248 11272
rect 18831 11232 19248 11260
rect 18831 11229 18843 11232
rect 18785 11223 18843 11229
rect 19242 11220 19248 11232
rect 19300 11220 19306 11272
rect 1104 11170 26864 11192
rect 1104 11118 10315 11170
rect 10367 11118 10379 11170
rect 10431 11118 10443 11170
rect 10495 11118 10507 11170
rect 10559 11118 19648 11170
rect 19700 11118 19712 11170
rect 19764 11118 19776 11170
rect 19828 11118 19840 11170
rect 19892 11118 26864 11170
rect 1104 11096 26864 11118
rect 10042 11016 10048 11068
rect 10100 11056 10106 11068
rect 10321 11059 10379 11065
rect 10321 11056 10333 11059
rect 10100 11028 10333 11056
rect 10100 11016 10106 11028
rect 10321 11025 10333 11028
rect 10367 11025 10379 11059
rect 13078 11056 13084 11068
rect 13039 11028 13084 11056
rect 10321 11019 10379 11025
rect 13078 11016 13084 11028
rect 13136 11016 13142 11068
rect 15562 11056 15568 11068
rect 15523 11028 15568 11056
rect 15562 11016 15568 11028
rect 15620 11016 15626 11068
rect 16758 11056 16764 11068
rect 16719 11028 16764 11056
rect 16758 11016 16764 11028
rect 16816 11016 16822 11068
rect 18046 11016 18052 11068
rect 18104 11056 18110 11068
rect 18325 11059 18383 11065
rect 18325 11056 18337 11059
rect 18104 11028 18337 11056
rect 18104 11016 18110 11028
rect 18325 11025 18337 11028
rect 18371 11056 18383 11059
rect 19337 11059 19395 11065
rect 19337 11056 19349 11059
rect 18371 11028 19349 11056
rect 18371 11025 18383 11028
rect 18325 11019 18383 11025
rect 19337 11025 19349 11028
rect 19383 11056 19395 11059
rect 19426 11056 19432 11068
rect 19383 11028 19432 11056
rect 19383 11025 19395 11028
rect 19337 11019 19395 11025
rect 19426 11016 19432 11028
rect 19484 11016 19490 11068
rect 24762 11056 24768 11068
rect 24723 11028 24768 11056
rect 24762 11016 24768 11028
rect 24820 11016 24826 11068
rect 16022 10988 16028 11000
rect 15935 10960 16028 10988
rect 16022 10948 16028 10960
rect 16080 10988 16086 11000
rect 18966 10988 18972 11000
rect 16080 10960 18972 10988
rect 16080 10948 16086 10960
rect 18966 10948 18972 10960
rect 19024 10948 19030 11000
rect 13170 10880 13176 10932
rect 13228 10920 13234 10932
rect 13449 10923 13507 10929
rect 13449 10920 13461 10923
rect 13228 10892 13461 10920
rect 13228 10880 13234 10892
rect 13449 10889 13461 10892
rect 13495 10889 13507 10923
rect 13449 10883 13507 10889
rect 15654 10880 15660 10932
rect 15712 10920 15718 10932
rect 15933 10923 15991 10929
rect 15933 10920 15945 10923
rect 15712 10892 15945 10920
rect 15712 10880 15718 10892
rect 15933 10889 15945 10892
rect 15979 10889 15991 10923
rect 15933 10883 15991 10889
rect 24581 10923 24639 10929
rect 24581 10889 24593 10923
rect 24627 10920 24639 10923
rect 24670 10920 24676 10932
rect 24627 10892 24676 10920
rect 24627 10889 24639 10892
rect 24581 10883 24639 10889
rect 24670 10880 24676 10892
rect 24728 10880 24734 10932
rect 13538 10852 13544 10864
rect 13499 10824 13544 10852
rect 13538 10812 13544 10824
rect 13596 10812 13602 10864
rect 13722 10852 13728 10864
rect 13683 10824 13728 10852
rect 13722 10812 13728 10824
rect 13780 10812 13786 10864
rect 16117 10855 16175 10861
rect 16117 10821 16129 10855
rect 16163 10821 16175 10855
rect 16117 10815 16175 10821
rect 12713 10787 12771 10793
rect 12713 10753 12725 10787
rect 12759 10784 12771 10787
rect 12802 10784 12808 10796
rect 12759 10756 12808 10784
rect 12759 10753 12771 10756
rect 12713 10747 12771 10753
rect 12802 10744 12808 10756
rect 12860 10784 12866 10796
rect 13740 10784 13768 10812
rect 12860 10756 13768 10784
rect 12860 10744 12866 10756
rect 15286 10744 15292 10796
rect 15344 10784 15350 10796
rect 16132 10784 16160 10815
rect 16298 10784 16304 10796
rect 15344 10756 16304 10784
rect 15344 10744 15350 10756
rect 16298 10744 16304 10756
rect 16356 10744 16362 10796
rect 1104 10626 26864 10648
rect 1104 10574 5648 10626
rect 5700 10574 5712 10626
rect 5764 10574 5776 10626
rect 5828 10574 5840 10626
rect 5892 10574 14982 10626
rect 15034 10574 15046 10626
rect 15098 10574 15110 10626
rect 15162 10574 15174 10626
rect 15226 10574 24315 10626
rect 24367 10574 24379 10626
rect 24431 10574 24443 10626
rect 24495 10574 24507 10626
rect 24559 10574 26864 10626
rect 1104 10552 26864 10574
rect 13814 10512 13820 10524
rect 13775 10484 13820 10512
rect 13814 10472 13820 10484
rect 13872 10472 13878 10524
rect 16022 10512 16028 10524
rect 15983 10484 16028 10512
rect 16022 10472 16028 10484
rect 16080 10472 16086 10524
rect 16298 10512 16304 10524
rect 16259 10484 16304 10512
rect 16298 10472 16304 10484
rect 16356 10472 16362 10524
rect 24489 10515 24547 10521
rect 24489 10481 24501 10515
rect 24535 10512 24547 10515
rect 24670 10512 24676 10524
rect 24535 10484 24676 10512
rect 24535 10481 24547 10484
rect 24489 10475 24547 10481
rect 24670 10472 24676 10484
rect 24728 10472 24734 10524
rect 13538 10444 13544 10456
rect 13451 10416 13544 10444
rect 13538 10404 13544 10416
rect 13596 10444 13602 10456
rect 16040 10444 16068 10472
rect 13596 10416 16068 10444
rect 13596 10404 13602 10416
rect 24118 10404 24124 10456
rect 24176 10444 24182 10456
rect 24765 10447 24823 10453
rect 24765 10444 24777 10447
rect 24176 10416 24777 10444
rect 24176 10404 24182 10416
rect 24765 10413 24777 10416
rect 24811 10413 24823 10447
rect 24765 10407 24823 10413
rect 23934 10268 23940 10320
rect 23992 10308 23998 10320
rect 24118 10308 24124 10320
rect 23992 10280 24124 10308
rect 23992 10268 23998 10280
rect 24118 10268 24124 10280
rect 24176 10268 24182 10320
rect 24581 10311 24639 10317
rect 24581 10277 24593 10311
rect 24627 10308 24639 10311
rect 24627 10280 25268 10308
rect 24627 10277 24639 10280
rect 24581 10271 24639 10277
rect 25240 10184 25268 10280
rect 13170 10172 13176 10184
rect 13131 10144 13176 10172
rect 13170 10132 13176 10144
rect 13228 10132 13234 10184
rect 15654 10172 15660 10184
rect 15615 10144 15660 10172
rect 15654 10132 15660 10144
rect 15712 10132 15718 10184
rect 25222 10172 25228 10184
rect 25183 10144 25228 10172
rect 25222 10132 25228 10144
rect 25280 10132 25286 10184
rect 1104 10082 26864 10104
rect 1104 10030 10315 10082
rect 10367 10030 10379 10082
rect 10431 10030 10443 10082
rect 10495 10030 10507 10082
rect 10559 10030 19648 10082
rect 19700 10030 19712 10082
rect 19764 10030 19776 10082
rect 19828 10030 19840 10082
rect 19892 10030 26864 10082
rect 1104 10008 26864 10030
rect 23290 9928 23296 9980
rect 23348 9968 23354 9980
rect 24765 9971 24823 9977
rect 24765 9968 24777 9971
rect 23348 9940 24777 9968
rect 23348 9928 23354 9940
rect 24765 9937 24777 9940
rect 24811 9937 24823 9971
rect 24765 9931 24823 9937
rect 24581 9835 24639 9841
rect 24581 9801 24593 9835
rect 24627 9832 24639 9835
rect 24670 9832 24676 9844
rect 24627 9804 24676 9832
rect 24627 9801 24639 9804
rect 24581 9795 24639 9801
rect 24670 9792 24676 9804
rect 24728 9792 24734 9844
rect 1104 9538 26864 9560
rect 1104 9486 5648 9538
rect 5700 9486 5712 9538
rect 5764 9486 5776 9538
rect 5828 9486 5840 9538
rect 5892 9486 14982 9538
rect 15034 9486 15046 9538
rect 15098 9486 15110 9538
rect 15162 9486 15174 9538
rect 15226 9486 24315 9538
rect 24367 9486 24379 9538
rect 24431 9486 24443 9538
rect 24495 9486 24507 9538
rect 24559 9486 26864 9538
rect 1104 9464 26864 9486
rect 24762 9356 24768 9368
rect 24723 9328 24768 9356
rect 24762 9316 24768 9328
rect 24820 9316 24826 9368
rect 25222 9356 25228 9368
rect 25183 9328 25228 9356
rect 25222 9316 25228 9328
rect 25280 9316 25286 9368
rect 24581 9223 24639 9229
rect 24581 9220 24593 9223
rect 24504 9192 24593 9220
rect 24504 9096 24532 9192
rect 24581 9189 24593 9192
rect 24627 9189 24639 9223
rect 24581 9183 24639 9189
rect 24486 9084 24492 9096
rect 24447 9056 24492 9084
rect 24486 9044 24492 9056
rect 24544 9044 24550 9096
rect 1104 8994 26864 9016
rect 1104 8942 10315 8994
rect 10367 8942 10379 8994
rect 10431 8942 10443 8994
rect 10495 8942 10507 8994
rect 10559 8942 19648 8994
rect 19700 8942 19712 8994
rect 19764 8942 19776 8994
rect 19828 8942 19840 8994
rect 19892 8942 26864 8994
rect 1104 8920 26864 8942
rect 24762 8880 24768 8892
rect 24723 8852 24768 8880
rect 24762 8840 24768 8852
rect 24820 8840 24826 8892
rect 24581 8747 24639 8753
rect 24581 8713 24593 8747
rect 24627 8744 24639 8747
rect 24670 8744 24676 8756
rect 24627 8716 24676 8744
rect 24627 8713 24639 8716
rect 24581 8707 24639 8713
rect 24670 8704 24676 8716
rect 24728 8704 24734 8756
rect 1104 8450 26864 8472
rect 1104 8398 5648 8450
rect 5700 8398 5712 8450
rect 5764 8398 5776 8450
rect 5828 8398 5840 8450
rect 5892 8398 14982 8450
rect 15034 8398 15046 8450
rect 15098 8398 15110 8450
rect 15162 8398 15174 8450
rect 15226 8398 24315 8450
rect 24367 8398 24379 8450
rect 24431 8398 24443 8450
rect 24495 8398 24507 8450
rect 24559 8398 26864 8450
rect 1104 8376 26864 8398
rect 24670 8336 24676 8348
rect 24631 8308 24676 8336
rect 24670 8296 24676 8308
rect 24728 8296 24734 8348
rect 1104 7906 26864 7928
rect 1104 7854 10315 7906
rect 10367 7854 10379 7906
rect 10431 7854 10443 7906
rect 10495 7854 10507 7906
rect 10559 7854 19648 7906
rect 19700 7854 19712 7906
rect 19764 7854 19776 7906
rect 19828 7854 19840 7906
rect 19892 7854 26864 7906
rect 1104 7832 26864 7854
rect 24578 7656 24584 7668
rect 24539 7628 24584 7656
rect 24578 7616 24584 7628
rect 24636 7616 24642 7668
rect 24762 7520 24768 7532
rect 24723 7492 24768 7520
rect 24762 7480 24768 7492
rect 24820 7480 24826 7532
rect 1104 7362 26864 7384
rect 1104 7310 5648 7362
rect 5700 7310 5712 7362
rect 5764 7310 5776 7362
rect 5828 7310 5840 7362
rect 5892 7310 14982 7362
rect 15034 7310 15046 7362
rect 15098 7310 15110 7362
rect 15162 7310 15174 7362
rect 15226 7310 24315 7362
rect 24367 7310 24379 7362
rect 24431 7310 24443 7362
rect 24495 7310 24507 7362
rect 24559 7310 26864 7362
rect 1104 7288 26864 7310
rect 17770 7248 17776 7260
rect 17731 7220 17776 7248
rect 17770 7208 17776 7220
rect 17828 7208 17834 7260
rect 24670 7248 24676 7260
rect 24631 7220 24676 7248
rect 24670 7208 24676 7220
rect 24728 7208 24734 7260
rect 18230 7112 18236 7124
rect 17604 7084 18236 7112
rect 17604 7053 17632 7084
rect 18230 7072 18236 7084
rect 18288 7072 18294 7124
rect 17589 7047 17647 7053
rect 17589 7013 17601 7047
rect 17635 7013 17647 7047
rect 17589 7007 17647 7013
rect 1104 6818 26864 6840
rect 1104 6766 10315 6818
rect 10367 6766 10379 6818
rect 10431 6766 10443 6818
rect 10495 6766 10507 6818
rect 10559 6766 19648 6818
rect 19700 6766 19712 6818
rect 19764 6766 19776 6818
rect 19828 6766 19840 6818
rect 19892 6766 26864 6818
rect 1104 6744 26864 6766
rect 1104 6274 26864 6296
rect 1104 6222 5648 6274
rect 5700 6222 5712 6274
rect 5764 6222 5776 6274
rect 5828 6222 5840 6274
rect 5892 6222 14982 6274
rect 15034 6222 15046 6274
rect 15098 6222 15110 6274
rect 15162 6222 15174 6274
rect 15226 6222 24315 6274
rect 24367 6222 24379 6274
rect 24431 6222 24443 6274
rect 24495 6222 24507 6274
rect 24559 6222 26864 6274
rect 1104 6200 26864 6222
rect 16393 6163 16451 6169
rect 16393 6129 16405 6163
rect 16439 6160 16451 6163
rect 16482 6160 16488 6172
rect 16439 6132 16488 6160
rect 16439 6129 16451 6132
rect 16393 6123 16451 6129
rect 16482 6120 16488 6132
rect 16540 6120 16546 6172
rect 16209 5959 16267 5965
rect 16209 5925 16221 5959
rect 16255 5925 16267 5959
rect 16209 5919 16267 5925
rect 16224 5888 16252 5919
rect 16850 5888 16856 5900
rect 16224 5860 16856 5888
rect 16850 5848 16856 5860
rect 16908 5848 16914 5900
rect 1104 5730 26864 5752
rect 1104 5678 10315 5730
rect 10367 5678 10379 5730
rect 10431 5678 10443 5730
rect 10495 5678 10507 5730
rect 10559 5678 19648 5730
rect 19700 5678 19712 5730
rect 19764 5678 19776 5730
rect 19828 5678 19840 5730
rect 19892 5678 26864 5730
rect 1104 5656 26864 5678
rect 1104 5186 26864 5208
rect 1104 5134 5648 5186
rect 5700 5134 5712 5186
rect 5764 5134 5776 5186
rect 5828 5134 5840 5186
rect 5892 5134 14982 5186
rect 15034 5134 15046 5186
rect 15098 5134 15110 5186
rect 15162 5134 15174 5186
rect 15226 5134 24315 5186
rect 24367 5134 24379 5186
rect 24431 5134 24443 5186
rect 24495 5134 24507 5186
rect 24559 5134 26864 5186
rect 1104 5112 26864 5134
rect 15473 5075 15531 5081
rect 15473 5041 15485 5075
rect 15519 5072 15531 5075
rect 16206 5072 16212 5084
rect 15519 5044 16212 5072
rect 15519 5041 15531 5044
rect 15473 5035 15531 5041
rect 16206 5032 16212 5044
rect 16264 5032 16270 5084
rect 15289 4871 15347 4877
rect 15289 4837 15301 4871
rect 15335 4837 15347 4871
rect 15289 4831 15347 4837
rect 15304 4800 15332 4831
rect 15930 4800 15936 4812
rect 15304 4772 15936 4800
rect 15930 4760 15936 4772
rect 15988 4760 15994 4812
rect 1104 4642 26864 4664
rect 1104 4590 10315 4642
rect 10367 4590 10379 4642
rect 10431 4590 10443 4642
rect 10495 4590 10507 4642
rect 10559 4590 19648 4642
rect 19700 4590 19712 4642
rect 19764 4590 19776 4642
rect 19828 4590 19840 4642
rect 19892 4590 26864 4642
rect 1104 4568 26864 4590
rect 1104 4098 26864 4120
rect 1104 4046 5648 4098
rect 5700 4046 5712 4098
rect 5764 4046 5776 4098
rect 5828 4046 5840 4098
rect 5892 4046 14982 4098
rect 15034 4046 15046 4098
rect 15098 4046 15110 4098
rect 15162 4046 15174 4098
rect 15226 4046 24315 4098
rect 24367 4046 24379 4098
rect 24431 4046 24443 4098
rect 24495 4046 24507 4098
rect 24559 4046 26864 4098
rect 1104 4024 26864 4046
rect 24581 3783 24639 3789
rect 24581 3749 24593 3783
rect 24627 3780 24639 3783
rect 24627 3752 25268 3780
rect 24627 3749 24639 3752
rect 24581 3743 24639 3749
rect 25240 3656 25268 3752
rect 24762 3644 24768 3656
rect 24723 3616 24768 3644
rect 24762 3604 24768 3616
rect 24820 3604 24826 3656
rect 25222 3644 25228 3656
rect 25183 3616 25228 3644
rect 25222 3604 25228 3616
rect 25280 3604 25286 3656
rect 1104 3554 26864 3576
rect 1104 3502 10315 3554
rect 10367 3502 10379 3554
rect 10431 3502 10443 3554
rect 10495 3502 10507 3554
rect 10559 3502 19648 3554
rect 19700 3502 19712 3554
rect 19764 3502 19776 3554
rect 19828 3502 19840 3554
rect 19892 3502 26864 3554
rect 1104 3480 26864 3502
rect 1104 3010 26864 3032
rect 1104 2958 5648 3010
rect 5700 2958 5712 3010
rect 5764 2958 5776 3010
rect 5828 2958 5840 3010
rect 5892 2958 14982 3010
rect 15034 2958 15046 3010
rect 15098 2958 15110 3010
rect 15162 2958 15174 3010
rect 15226 2958 24315 3010
rect 24367 2958 24379 3010
rect 24431 2958 24443 3010
rect 24495 2958 24507 3010
rect 24559 2958 26864 3010
rect 1104 2936 26864 2958
rect 1104 2466 26864 2488
rect 1104 2414 10315 2466
rect 10367 2414 10379 2466
rect 10431 2414 10443 2466
rect 10495 2414 10507 2466
rect 10559 2414 19648 2466
rect 19700 2414 19712 2466
rect 19764 2414 19776 2466
rect 19828 2414 19840 2466
rect 19892 2414 26864 2466
rect 1104 2392 26864 2414
rect 1104 1922 26864 1944
rect 1104 1870 5648 1922
rect 5700 1870 5712 1922
rect 5764 1870 5776 1922
rect 5828 1870 5840 1922
rect 5892 1870 14982 1922
rect 15034 1870 15046 1922
rect 15098 1870 15110 1922
rect 15162 1870 15174 1922
rect 15226 1870 24315 1922
rect 24367 1870 24379 1922
rect 24431 1870 24443 1922
rect 24495 1870 24507 1922
rect 24559 1870 26864 1922
rect 1104 1848 26864 1870
<< via1 >>
rect 296 27132 348 27184
rect 480 27132 532 27184
rect 10315 25262 10367 25314
rect 10379 25262 10431 25314
rect 10443 25262 10495 25314
rect 10507 25262 10559 25314
rect 19648 25262 19700 25314
rect 19712 25262 19764 25314
rect 19776 25262 19828 25314
rect 19840 25262 19892 25314
rect 23572 25160 23624 25212
rect 24768 25203 24820 25212
rect 24768 25169 24777 25203
rect 24777 25169 24811 25203
rect 24811 25169 24820 25203
rect 24768 25160 24820 25169
rect 22836 25067 22888 25076
rect 22836 25033 22845 25067
rect 22845 25033 22879 25067
rect 22879 25033 22888 25067
rect 22836 25024 22888 25033
rect 24768 24956 24820 25008
rect 11428 24863 11480 24872
rect 11428 24829 11437 24863
rect 11437 24829 11471 24863
rect 11471 24829 11480 24863
rect 11428 24820 11480 24829
rect 5648 24718 5700 24770
rect 5712 24718 5764 24770
rect 5776 24718 5828 24770
rect 5840 24718 5892 24770
rect 14982 24718 15034 24770
rect 15046 24718 15098 24770
rect 15110 24718 15162 24770
rect 15174 24718 15226 24770
rect 24315 24718 24367 24770
rect 24379 24718 24431 24770
rect 24443 24718 24495 24770
rect 24507 24718 24559 24770
rect 22836 24548 22888 24600
rect 11244 24480 11296 24532
rect 15292 24480 15344 24532
rect 16212 24480 16264 24532
rect 18696 24480 18748 24532
rect 19156 24480 19208 24532
rect 21364 24480 21416 24532
rect 22008 24480 22060 24532
rect 23756 24480 23808 24532
rect 24676 24480 24728 24532
rect 11060 24412 11112 24464
rect 11428 24412 11480 24464
rect 20720 24412 20772 24464
rect 21640 24412 21692 24464
rect 22560 24455 22612 24464
rect 22560 24421 22569 24455
rect 22569 24421 22603 24455
rect 22603 24421 22612 24455
rect 22560 24412 22612 24421
rect 23848 24412 23900 24464
rect 24216 24412 24268 24464
rect 11244 24319 11296 24328
rect 11244 24285 11253 24319
rect 11253 24285 11287 24319
rect 11287 24285 11296 24319
rect 11244 24276 11296 24285
rect 12348 24344 12400 24396
rect 24676 24344 24728 24396
rect 11796 24319 11848 24328
rect 11796 24285 11805 24319
rect 11805 24285 11839 24319
rect 11839 24285 11848 24319
rect 11796 24276 11848 24285
rect 16856 24276 16908 24328
rect 17408 24319 17460 24328
rect 17408 24285 17417 24319
rect 17417 24285 17451 24319
rect 17451 24285 17460 24319
rect 17408 24276 17460 24285
rect 23388 24276 23440 24328
rect 23848 24276 23900 24328
rect 24768 24319 24820 24328
rect 24768 24285 24777 24319
rect 24777 24285 24811 24319
rect 24811 24285 24820 24319
rect 24768 24276 24820 24285
rect 25136 24319 25188 24328
rect 25136 24285 25145 24319
rect 25145 24285 25179 24319
rect 25179 24285 25188 24319
rect 25136 24276 25188 24285
rect 10315 24174 10367 24226
rect 10379 24174 10431 24226
rect 10443 24174 10495 24226
rect 10507 24174 10559 24226
rect 19648 24174 19700 24226
rect 19712 24174 19764 24226
rect 19776 24174 19828 24226
rect 19840 24174 19892 24226
rect 22744 24072 22796 24124
rect 24216 24004 24268 24056
rect 13176 23936 13228 23988
rect 15108 23936 15160 23988
rect 15476 23936 15528 23988
rect 15936 23936 15988 23988
rect 18144 23936 18196 23988
rect 19248 23979 19300 23988
rect 19248 23945 19257 23979
rect 19257 23945 19291 23979
rect 19291 23945 19300 23979
rect 19248 23936 19300 23945
rect 21088 23936 21140 23988
rect 22284 23936 22336 23988
rect 23664 23979 23716 23988
rect 23664 23945 23673 23979
rect 23673 23945 23707 23979
rect 23707 23945 23716 23979
rect 23664 23936 23716 23945
rect 24676 23936 24728 23988
rect 13820 23868 13872 23920
rect 16120 23868 16172 23920
rect 16856 23911 16908 23920
rect 16856 23877 16865 23911
rect 16865 23877 16899 23911
rect 16899 23877 16908 23911
rect 16856 23868 16908 23877
rect 18420 23868 18472 23920
rect 19432 23800 19484 23852
rect 19984 23800 20036 23852
rect 21456 23800 21508 23852
rect 23296 23800 23348 23852
rect 25136 23843 25188 23852
rect 25136 23809 25145 23843
rect 25145 23809 25179 23843
rect 25179 23809 25188 23843
rect 25136 23800 25188 23809
rect 25228 23800 25280 23852
rect 26148 23800 26200 23852
rect 11060 23732 11112 23784
rect 11796 23732 11848 23784
rect 14280 23732 14332 23784
rect 16304 23775 16356 23784
rect 16304 23741 16313 23775
rect 16313 23741 16347 23775
rect 16347 23741 16356 23775
rect 16304 23732 16356 23741
rect 18328 23775 18380 23784
rect 18328 23741 18337 23775
rect 18337 23741 18371 23775
rect 18371 23741 18380 23775
rect 18328 23732 18380 23741
rect 18696 23775 18748 23784
rect 18696 23741 18705 23775
rect 18705 23741 18739 23775
rect 18739 23741 18748 23775
rect 18696 23732 18748 23741
rect 20536 23775 20588 23784
rect 20536 23741 20545 23775
rect 20545 23741 20579 23775
rect 20579 23741 20588 23775
rect 20536 23732 20588 23741
rect 24216 23732 24268 23784
rect 5648 23630 5700 23682
rect 5712 23630 5764 23682
rect 5776 23630 5828 23682
rect 5840 23630 5892 23682
rect 14982 23630 15034 23682
rect 15046 23630 15098 23682
rect 15110 23630 15162 23682
rect 15174 23630 15226 23682
rect 24315 23630 24367 23682
rect 24379 23630 24431 23682
rect 24443 23630 24495 23682
rect 24507 23630 24559 23682
rect 13176 23571 13228 23580
rect 13176 23537 13185 23571
rect 13185 23537 13219 23571
rect 13219 23537 13228 23571
rect 13176 23528 13228 23537
rect 13452 23571 13504 23580
rect 13452 23537 13461 23571
rect 13461 23537 13495 23571
rect 13495 23537 13504 23571
rect 13452 23528 13504 23537
rect 16120 23528 16172 23580
rect 18144 23571 18196 23580
rect 18144 23537 18153 23571
rect 18153 23537 18187 23571
rect 18187 23537 18196 23571
rect 18144 23528 18196 23537
rect 18420 23571 18472 23580
rect 18420 23537 18429 23571
rect 18429 23537 18463 23571
rect 18463 23537 18472 23571
rect 18420 23528 18472 23537
rect 19984 23571 20036 23580
rect 19984 23537 19993 23571
rect 19993 23537 20027 23571
rect 20027 23537 20036 23571
rect 19984 23528 20036 23537
rect 23664 23571 23716 23580
rect 23664 23537 23673 23571
rect 23673 23537 23707 23571
rect 23707 23537 23716 23571
rect 23664 23528 23716 23537
rect 24676 23528 24728 23580
rect 22100 23503 22152 23512
rect 22100 23469 22109 23503
rect 22109 23469 22143 23503
rect 22143 23469 22152 23503
rect 22100 23460 22152 23469
rect 14280 23435 14332 23444
rect 14280 23401 14289 23435
rect 14289 23401 14323 23435
rect 14323 23401 14332 23435
rect 14280 23392 14332 23401
rect 20536 23392 20588 23444
rect 21456 23435 21508 23444
rect 21456 23401 21465 23435
rect 21465 23401 21499 23435
rect 21499 23401 21508 23435
rect 21456 23392 21508 23401
rect 11336 23367 11388 23376
rect 11336 23333 11345 23367
rect 11345 23333 11379 23367
rect 11379 23333 11388 23367
rect 11336 23324 11388 23333
rect 12164 23256 12216 23308
rect 13820 23324 13872 23376
rect 18144 23324 18196 23376
rect 18696 23324 18748 23376
rect 19432 23324 19484 23376
rect 22836 23392 22888 23444
rect 24768 23392 24820 23444
rect 23664 23324 23716 23376
rect 24216 23324 24268 23376
rect 15936 23299 15988 23308
rect 15936 23265 15945 23299
rect 15945 23265 15979 23299
rect 15979 23265 15988 23299
rect 15936 23256 15988 23265
rect 16856 23256 16908 23308
rect 17316 23256 17368 23308
rect 18328 23256 18380 23308
rect 19340 23256 19392 23308
rect 20536 23256 20588 23308
rect 22376 23299 22428 23308
rect 22376 23265 22385 23299
rect 22385 23265 22419 23299
rect 22419 23265 22428 23299
rect 22376 23256 22428 23265
rect 12256 23188 12308 23240
rect 13820 23188 13872 23240
rect 14004 23231 14056 23240
rect 14004 23197 14013 23231
rect 14013 23197 14047 23231
rect 14047 23197 14056 23231
rect 14004 23188 14056 23197
rect 15292 23231 15344 23240
rect 15292 23197 15301 23231
rect 15301 23197 15335 23231
rect 15335 23197 15344 23231
rect 15292 23188 15344 23197
rect 17224 23188 17276 23240
rect 20720 23231 20772 23240
rect 20720 23197 20729 23231
rect 20729 23197 20763 23231
rect 20763 23197 20772 23231
rect 20720 23188 20772 23197
rect 23572 23188 23624 23240
rect 10315 23086 10367 23138
rect 10379 23086 10431 23138
rect 10443 23086 10495 23138
rect 10507 23086 10559 23138
rect 19648 23086 19700 23138
rect 19712 23086 19764 23138
rect 19776 23086 19828 23138
rect 19840 23086 19892 23138
rect 10968 22984 11020 23036
rect 11060 22984 11112 23036
rect 11888 22984 11940 23036
rect 15200 22984 15252 23036
rect 17408 22984 17460 23036
rect 19432 23027 19484 23036
rect 19432 22993 19441 23027
rect 19441 22993 19475 23027
rect 19475 22993 19484 23027
rect 19432 22984 19484 22993
rect 23572 22984 23624 23036
rect 24124 23027 24176 23036
rect 24124 22993 24133 23027
rect 24133 22993 24167 23027
rect 24167 22993 24176 23027
rect 24124 22984 24176 22993
rect 25412 23027 25464 23036
rect 25412 22993 25421 23027
rect 25421 22993 25455 23027
rect 25455 22993 25464 23027
rect 25412 22984 25464 22993
rect 14280 22916 14332 22968
rect 16304 22916 16356 22968
rect 19340 22916 19392 22968
rect 21180 22916 21232 22968
rect 24216 22916 24268 22968
rect 11152 22891 11204 22900
rect 11152 22857 11161 22891
rect 11161 22857 11195 22891
rect 11195 22857 11204 22891
rect 11152 22848 11204 22857
rect 12440 22891 12492 22900
rect 12440 22857 12449 22891
rect 12449 22857 12483 22891
rect 12483 22857 12492 22891
rect 12440 22848 12492 22857
rect 12992 22848 13044 22900
rect 18328 22891 18380 22900
rect 18328 22857 18351 22891
rect 18351 22857 18380 22891
rect 18328 22848 18380 22857
rect 20352 22848 20404 22900
rect 21364 22891 21416 22900
rect 21364 22857 21387 22891
rect 21387 22857 21416 22891
rect 21364 22848 21416 22857
rect 25688 22848 25740 22900
rect 11612 22780 11664 22832
rect 12256 22780 12308 22832
rect 13728 22780 13780 22832
rect 10876 22712 10928 22764
rect 13728 22687 13780 22696
rect 13728 22653 13737 22687
rect 13737 22653 13771 22687
rect 13771 22653 13780 22687
rect 13728 22644 13780 22653
rect 17224 22780 17276 22832
rect 18052 22823 18104 22832
rect 18052 22789 18061 22823
rect 18061 22789 18095 22823
rect 18095 22789 18104 22823
rect 18052 22780 18104 22789
rect 20996 22780 21048 22832
rect 23940 22780 23992 22832
rect 16396 22755 16448 22764
rect 16396 22721 16405 22755
rect 16405 22721 16439 22755
rect 16439 22721 16448 22755
rect 16396 22712 16448 22721
rect 14096 22644 14148 22696
rect 16028 22687 16080 22696
rect 16028 22653 16037 22687
rect 16037 22653 16071 22687
rect 16071 22653 16080 22687
rect 16028 22644 16080 22653
rect 20444 22644 20496 22696
rect 22468 22687 22520 22696
rect 22468 22653 22477 22687
rect 22477 22653 22511 22687
rect 22511 22653 22520 22687
rect 22468 22644 22520 22653
rect 22836 22687 22888 22696
rect 22836 22653 22845 22687
rect 22845 22653 22879 22687
rect 22879 22653 22888 22687
rect 22836 22644 22888 22653
rect 24860 22644 24912 22696
rect 5648 22542 5700 22594
rect 5712 22542 5764 22594
rect 5776 22542 5828 22594
rect 5840 22542 5892 22594
rect 14982 22542 15034 22594
rect 15046 22542 15098 22594
rect 15110 22542 15162 22594
rect 15174 22542 15226 22594
rect 24315 22542 24367 22594
rect 24379 22542 24431 22594
rect 24443 22542 24495 22594
rect 24507 22542 24559 22594
rect 11060 22440 11112 22492
rect 12716 22483 12768 22492
rect 12716 22449 12725 22483
rect 12725 22449 12759 22483
rect 12759 22449 12768 22483
rect 12716 22440 12768 22449
rect 12992 22483 13044 22492
rect 12992 22449 13001 22483
rect 13001 22449 13035 22483
rect 13035 22449 13044 22483
rect 12992 22440 13044 22449
rect 14280 22483 14332 22492
rect 14280 22449 14289 22483
rect 14289 22449 14323 22483
rect 14323 22449 14332 22483
rect 14280 22440 14332 22449
rect 17316 22483 17368 22492
rect 17316 22449 17325 22483
rect 17325 22449 17359 22483
rect 17359 22449 17368 22483
rect 17316 22440 17368 22449
rect 17408 22440 17460 22492
rect 18144 22483 18196 22492
rect 18144 22449 18153 22483
rect 18153 22449 18187 22483
rect 18187 22449 18196 22483
rect 18144 22440 18196 22449
rect 18328 22440 18380 22492
rect 20352 22483 20404 22492
rect 20352 22449 20361 22483
rect 20361 22449 20395 22483
rect 20395 22449 20404 22483
rect 20352 22440 20404 22449
rect 20996 22440 21048 22492
rect 11336 22347 11388 22356
rect 11336 22313 11345 22347
rect 11345 22313 11379 22347
rect 11379 22313 11388 22347
rect 11336 22304 11388 22313
rect 14096 22304 14148 22356
rect 15384 22304 15436 22356
rect 15936 22347 15988 22356
rect 15936 22313 15945 22347
rect 15945 22313 15979 22347
rect 15979 22313 15988 22347
rect 15936 22304 15988 22313
rect 20628 22304 20680 22356
rect 11152 22236 11204 22288
rect 11612 22279 11664 22288
rect 11612 22245 11646 22279
rect 11646 22245 11664 22279
rect 11612 22236 11664 22245
rect 16028 22236 16080 22288
rect 16488 22236 16540 22288
rect 20444 22236 20496 22288
rect 22468 22304 22520 22356
rect 23204 22440 23256 22492
rect 23940 22483 23992 22492
rect 23940 22449 23949 22483
rect 23949 22449 23983 22483
rect 23983 22449 23992 22483
rect 23940 22440 23992 22449
rect 24124 22440 24176 22492
rect 24768 22279 24820 22288
rect 24768 22245 24777 22279
rect 24777 22245 24811 22279
rect 24811 22245 24820 22279
rect 24768 22236 24820 22245
rect 11796 22168 11848 22220
rect 15568 22168 15620 22220
rect 20720 22211 20772 22220
rect 20720 22177 20729 22211
rect 20729 22177 20763 22211
rect 20763 22177 20772 22211
rect 20720 22168 20772 22177
rect 22836 22211 22888 22220
rect 22836 22177 22870 22211
rect 22870 22177 22888 22211
rect 22836 22168 22888 22177
rect 23388 22168 23440 22220
rect 20904 22143 20956 22152
rect 20904 22109 20913 22143
rect 20913 22109 20947 22143
rect 20947 22109 20956 22143
rect 20904 22100 20956 22109
rect 21180 22100 21232 22152
rect 21732 22100 21784 22152
rect 24216 22143 24268 22152
rect 24216 22109 24225 22143
rect 24225 22109 24259 22143
rect 24259 22109 24268 22143
rect 24216 22100 24268 22109
rect 24952 22143 25004 22152
rect 24952 22109 24961 22143
rect 24961 22109 24995 22143
rect 24995 22109 25004 22143
rect 24952 22100 25004 22109
rect 25688 22143 25740 22152
rect 25688 22109 25697 22143
rect 25697 22109 25731 22143
rect 25731 22109 25740 22143
rect 25688 22100 25740 22109
rect 10315 21998 10367 22050
rect 10379 21998 10431 22050
rect 10443 21998 10495 22050
rect 10507 21998 10559 22050
rect 19648 21998 19700 22050
rect 19712 21998 19764 22050
rect 19776 21998 19828 22050
rect 19840 21998 19892 22050
rect 480 21828 532 21880
rect 11612 21896 11664 21948
rect 14372 21896 14424 21948
rect 15108 21896 15160 21948
rect 17224 21939 17276 21948
rect 17224 21905 17233 21939
rect 17233 21905 17267 21939
rect 17267 21905 17276 21939
rect 17224 21896 17276 21905
rect 24216 21896 24268 21948
rect 19984 21828 20036 21880
rect 20444 21828 20496 21880
rect 23940 21871 23992 21880
rect 23940 21837 23949 21871
rect 23949 21837 23983 21871
rect 23983 21837 23992 21871
rect 23940 21828 23992 21837
rect 13820 21760 13872 21812
rect 17040 21760 17092 21812
rect 18328 21803 18380 21812
rect 480 21692 532 21744
rect 14832 21735 14884 21744
rect 14832 21701 14841 21735
rect 14841 21701 14875 21735
rect 14875 21701 14884 21735
rect 14832 21692 14884 21701
rect 16028 21692 16080 21744
rect 16856 21735 16908 21744
rect 16856 21701 16865 21735
rect 16865 21701 16899 21735
rect 16899 21701 16908 21735
rect 16856 21692 16908 21701
rect 14280 21667 14332 21676
rect 14280 21633 14289 21667
rect 14289 21633 14323 21667
rect 14323 21633 14332 21667
rect 14280 21624 14332 21633
rect 18328 21769 18337 21803
rect 18337 21769 18371 21803
rect 18371 21769 18380 21803
rect 18328 21760 18380 21769
rect 24124 21760 24176 21812
rect 20168 21692 20220 21744
rect 12624 21556 12676 21608
rect 15752 21599 15804 21608
rect 15752 21565 15761 21599
rect 15761 21565 15795 21599
rect 15795 21565 15804 21599
rect 15752 21556 15804 21565
rect 16396 21556 16448 21608
rect 16488 21556 16540 21608
rect 16856 21556 16908 21608
rect 21548 21556 21600 21608
rect 23388 21556 23440 21608
rect 24768 21599 24820 21608
rect 24768 21565 24777 21599
rect 24777 21565 24811 21599
rect 24811 21565 24820 21599
rect 24768 21556 24820 21565
rect 5648 21454 5700 21506
rect 5712 21454 5764 21506
rect 5776 21454 5828 21506
rect 5840 21454 5892 21506
rect 14982 21454 15034 21506
rect 15046 21454 15098 21506
rect 15110 21454 15162 21506
rect 15174 21454 15226 21506
rect 24315 21454 24367 21506
rect 24379 21454 24431 21506
rect 24443 21454 24495 21506
rect 24507 21454 24559 21506
rect 11520 21395 11572 21404
rect 11520 21361 11529 21395
rect 11529 21361 11563 21395
rect 11563 21361 11572 21395
rect 14372 21395 14424 21404
rect 11520 21352 11572 21361
rect 14372 21361 14381 21395
rect 14381 21361 14415 21395
rect 14415 21361 14424 21395
rect 14372 21352 14424 21361
rect 14832 21352 14884 21404
rect 15568 21395 15620 21404
rect 15568 21361 15577 21395
rect 15577 21361 15611 21395
rect 15611 21361 15620 21395
rect 15568 21352 15620 21361
rect 16028 21395 16080 21404
rect 16028 21361 16037 21395
rect 16037 21361 16071 21395
rect 16071 21361 16080 21395
rect 16028 21352 16080 21361
rect 19984 21395 20036 21404
rect 19984 21361 19993 21395
rect 19993 21361 20027 21395
rect 20027 21361 20036 21395
rect 19984 21352 20036 21361
rect 22928 21395 22980 21404
rect 22928 21361 22937 21395
rect 22937 21361 22971 21395
rect 22971 21361 22980 21395
rect 22928 21352 22980 21361
rect 24124 21352 24176 21404
rect 12624 21216 12676 21268
rect 16488 21216 16540 21268
rect 17592 21216 17644 21268
rect 19248 21216 19300 21268
rect 20536 21216 20588 21268
rect 21548 21216 21600 21268
rect 11704 21055 11756 21064
rect 11704 21021 11713 21055
rect 11713 21021 11747 21055
rect 11747 21021 11756 21055
rect 11704 21012 11756 21021
rect 11796 21012 11848 21064
rect 12440 21012 12492 21064
rect 20904 21148 20956 21200
rect 13544 21123 13596 21132
rect 13544 21089 13553 21123
rect 13553 21089 13587 21123
rect 13587 21089 13596 21123
rect 13544 21080 13596 21089
rect 20996 21080 21048 21132
rect 25136 21191 25188 21200
rect 25136 21157 25145 21191
rect 25145 21157 25179 21191
rect 25179 21157 25188 21191
rect 25136 21148 25188 21157
rect 26240 21080 26292 21132
rect 27528 21080 27580 21132
rect 15844 21055 15896 21064
rect 15844 21021 15853 21055
rect 15853 21021 15887 21055
rect 15887 21021 15896 21055
rect 15844 21012 15896 21021
rect 16396 21055 16448 21064
rect 16396 21021 16405 21055
rect 16405 21021 16439 21055
rect 16439 21021 16448 21055
rect 16396 21012 16448 21021
rect 17040 21055 17092 21064
rect 17040 21021 17049 21055
rect 17049 21021 17083 21055
rect 17083 21021 17092 21055
rect 17040 21012 17092 21021
rect 17592 21055 17644 21064
rect 17592 21021 17601 21055
rect 17601 21021 17635 21055
rect 17635 21021 17644 21055
rect 17592 21012 17644 21021
rect 18052 21055 18104 21064
rect 18052 21021 18061 21055
rect 18061 21021 18095 21055
rect 18095 21021 18104 21055
rect 18052 21012 18104 21021
rect 18144 21055 18196 21064
rect 18144 21021 18153 21055
rect 18153 21021 18187 21055
rect 18187 21021 18196 21055
rect 18144 21012 18196 21021
rect 18604 21055 18656 21064
rect 18604 21021 18613 21055
rect 18613 21021 18647 21055
rect 18647 21021 18656 21055
rect 18604 21012 18656 21021
rect 20168 21012 20220 21064
rect 20904 21055 20956 21064
rect 20904 21021 20913 21055
rect 20913 21021 20947 21055
rect 20947 21021 20956 21055
rect 20904 21012 20956 21021
rect 23664 21055 23716 21064
rect 23664 21021 23673 21055
rect 23673 21021 23707 21055
rect 23707 21021 23716 21055
rect 23664 21012 23716 21021
rect 25320 21055 25372 21064
rect 25320 21021 25329 21055
rect 25329 21021 25363 21055
rect 25363 21021 25372 21055
rect 25320 21012 25372 21021
rect 10315 20910 10367 20962
rect 10379 20910 10431 20962
rect 10443 20910 10495 20962
rect 10507 20910 10559 20962
rect 19648 20910 19700 20962
rect 19712 20910 19764 20962
rect 19776 20910 19828 20962
rect 19840 20910 19892 20962
rect 13820 20808 13872 20860
rect 14648 20851 14700 20860
rect 14648 20817 14657 20851
rect 14657 20817 14691 20851
rect 14691 20817 14700 20851
rect 14648 20808 14700 20817
rect 16856 20808 16908 20860
rect 18604 20808 18656 20860
rect 22192 20808 22244 20860
rect 24676 20808 24728 20860
rect 12624 20740 12676 20792
rect 18420 20783 18472 20792
rect 18420 20749 18429 20783
rect 18429 20749 18463 20783
rect 18463 20749 18472 20783
rect 18420 20740 18472 20749
rect 20536 20740 20588 20792
rect 24860 20740 24912 20792
rect 15292 20672 15344 20724
rect 15752 20672 15804 20724
rect 16488 20672 16540 20724
rect 23848 20715 23900 20724
rect 23848 20681 23857 20715
rect 23857 20681 23891 20715
rect 23891 20681 23900 20715
rect 23848 20672 23900 20681
rect 25320 20672 25372 20724
rect 12440 20647 12492 20656
rect 12440 20613 12449 20647
rect 12449 20613 12483 20647
rect 12483 20613 12492 20647
rect 12440 20604 12492 20613
rect 15384 20604 15436 20656
rect 15660 20647 15712 20656
rect 15660 20613 15669 20647
rect 15669 20613 15703 20647
rect 15703 20613 15712 20647
rect 15660 20604 15712 20613
rect 17960 20604 18012 20656
rect 19064 20604 19116 20656
rect 20168 20647 20220 20656
rect 20168 20613 20177 20647
rect 20177 20613 20211 20647
rect 20211 20613 20220 20647
rect 20168 20604 20220 20613
rect 24860 20604 24912 20656
rect 25504 20604 25556 20656
rect 11796 20511 11848 20520
rect 11796 20477 11805 20511
rect 11805 20477 11839 20511
rect 11839 20477 11848 20511
rect 11796 20468 11848 20477
rect 13820 20511 13872 20520
rect 13820 20477 13829 20511
rect 13829 20477 13863 20511
rect 13863 20477 13872 20511
rect 13820 20468 13872 20477
rect 15384 20511 15436 20520
rect 15384 20477 15393 20511
rect 15393 20477 15427 20511
rect 15427 20477 15436 20511
rect 15384 20468 15436 20477
rect 20812 20468 20864 20520
rect 22836 20511 22888 20520
rect 22836 20477 22845 20511
rect 22845 20477 22879 20511
rect 22879 20477 22888 20511
rect 22836 20468 22888 20477
rect 5648 20366 5700 20418
rect 5712 20366 5764 20418
rect 5776 20366 5828 20418
rect 5840 20366 5892 20418
rect 14982 20366 15034 20418
rect 15046 20366 15098 20418
rect 15110 20366 15162 20418
rect 15174 20366 15226 20418
rect 24315 20366 24367 20418
rect 24379 20366 24431 20418
rect 24443 20366 24495 20418
rect 24507 20366 24559 20418
rect 12440 20264 12492 20316
rect 15292 20264 15344 20316
rect 16488 20264 16540 20316
rect 17960 20307 18012 20316
rect 17960 20273 17969 20307
rect 17969 20273 18003 20307
rect 18003 20273 18012 20307
rect 17960 20264 18012 20273
rect 19340 20264 19392 20316
rect 20536 20307 20588 20316
rect 20536 20273 20545 20307
rect 20545 20273 20579 20307
rect 20579 20273 20588 20307
rect 20536 20264 20588 20273
rect 23480 20264 23532 20316
rect 19064 20196 19116 20248
rect 20812 20196 20864 20248
rect 23848 20264 23900 20316
rect 25136 20307 25188 20316
rect 25136 20273 25145 20307
rect 25145 20273 25179 20307
rect 25179 20273 25188 20307
rect 25136 20264 25188 20273
rect 25320 20264 25372 20316
rect 12440 20060 12492 20112
rect 12716 20103 12768 20112
rect 12716 20069 12725 20103
rect 12725 20069 12759 20103
rect 12759 20069 12768 20103
rect 12716 20060 12768 20069
rect 12992 20103 13044 20112
rect 12992 20069 13026 20103
rect 13026 20069 13044 20103
rect 12992 20060 13044 20069
rect 13728 20060 13780 20112
rect 10876 19992 10928 20044
rect 12624 19992 12676 20044
rect 13268 19992 13320 20044
rect 15384 20060 15436 20112
rect 14096 19967 14148 19976
rect 14096 19933 14105 19967
rect 14105 19933 14139 19967
rect 14139 19933 14148 19967
rect 14096 19924 14148 19933
rect 15016 19967 15068 19976
rect 15016 19933 15025 19967
rect 15025 19933 15059 19967
rect 15059 19933 15068 19967
rect 15016 19924 15068 19933
rect 15660 19924 15712 19976
rect 20996 20128 21048 20180
rect 22560 20060 22612 20112
rect 19248 19992 19300 20044
rect 20168 20035 20220 20044
rect 20168 20001 20177 20035
rect 20177 20001 20211 20035
rect 20211 20001 20220 20035
rect 20168 19992 20220 20001
rect 22836 20060 22888 20112
rect 23480 20060 23532 20112
rect 23940 20060 23992 20112
rect 22652 19967 22704 19976
rect 22652 19933 22661 19967
rect 22661 19933 22695 19967
rect 22695 19933 22704 19967
rect 22652 19924 22704 19933
rect 24952 19924 25004 19976
rect 10315 19822 10367 19874
rect 10379 19822 10431 19874
rect 10443 19822 10495 19874
rect 10507 19822 10559 19874
rect 19648 19822 19700 19874
rect 19712 19822 19764 19874
rect 19776 19822 19828 19874
rect 19840 19822 19892 19874
rect 10876 19720 10928 19772
rect 11704 19720 11756 19772
rect 12992 19763 13044 19772
rect 12992 19729 13001 19763
rect 13001 19729 13035 19763
rect 13035 19729 13044 19763
rect 12992 19720 13044 19729
rect 13268 19763 13320 19772
rect 13268 19729 13277 19763
rect 13277 19729 13311 19763
rect 13311 19729 13320 19763
rect 13268 19720 13320 19729
rect 15384 19720 15436 19772
rect 17960 19720 18012 19772
rect 18420 19720 18472 19772
rect 24768 19720 24820 19772
rect 25412 19763 25464 19772
rect 25412 19729 25421 19763
rect 25421 19729 25455 19763
rect 25455 19729 25464 19763
rect 25412 19720 25464 19729
rect 14096 19652 14148 19704
rect 15660 19652 15712 19704
rect 12716 19584 12768 19636
rect 14740 19584 14792 19636
rect 15016 19584 15068 19636
rect 18144 19584 18196 19636
rect 18696 19627 18748 19636
rect 18696 19593 18705 19627
rect 18705 19593 18739 19627
rect 18739 19593 18748 19627
rect 18696 19584 18748 19593
rect 18972 19627 19024 19636
rect 18972 19593 18981 19627
rect 18981 19593 19015 19627
rect 19015 19593 19024 19627
rect 18972 19584 19024 19593
rect 12440 19559 12492 19568
rect 12440 19525 12449 19559
rect 12449 19525 12483 19559
rect 12483 19525 12492 19559
rect 12440 19516 12492 19525
rect 15660 19516 15712 19568
rect 20996 19423 21048 19432
rect 20996 19389 21005 19423
rect 21005 19389 21039 19423
rect 21039 19389 21048 19423
rect 20996 19380 21048 19389
rect 21548 19380 21600 19432
rect 24032 19627 24084 19636
rect 24032 19593 24041 19627
rect 24041 19593 24075 19627
rect 24075 19593 24084 19627
rect 24032 19584 24084 19593
rect 24860 19584 24912 19636
rect 25872 19584 25924 19636
rect 22100 19516 22152 19568
rect 22560 19559 22612 19568
rect 22560 19525 22569 19559
rect 22569 19525 22603 19559
rect 22603 19525 22612 19559
rect 22560 19516 22612 19525
rect 22836 19516 22888 19568
rect 24124 19516 24176 19568
rect 23664 19423 23716 19432
rect 23664 19389 23673 19423
rect 23673 19389 23707 19423
rect 23707 19389 23716 19423
rect 23664 19380 23716 19389
rect 5648 19278 5700 19330
rect 5712 19278 5764 19330
rect 5776 19278 5828 19330
rect 5840 19278 5892 19330
rect 14982 19278 15034 19330
rect 15046 19278 15098 19330
rect 15110 19278 15162 19330
rect 15174 19278 15226 19330
rect 24315 19278 24367 19330
rect 24379 19278 24431 19330
rect 24443 19278 24495 19330
rect 24507 19278 24559 19330
rect 14740 19219 14792 19228
rect 14740 19185 14749 19219
rect 14749 19185 14783 19219
rect 14783 19185 14792 19219
rect 14740 19176 14792 19185
rect 18696 19219 18748 19228
rect 18696 19185 18705 19219
rect 18705 19185 18739 19219
rect 18739 19185 18748 19219
rect 18696 19176 18748 19185
rect 24032 19176 24084 19228
rect 24768 19219 24820 19228
rect 24768 19185 24777 19219
rect 24777 19185 24811 19219
rect 24811 19185 24820 19219
rect 24768 19176 24820 19185
rect 25872 19219 25924 19228
rect 25872 19185 25881 19219
rect 25881 19185 25915 19219
rect 25915 19185 25924 19219
rect 25872 19176 25924 19185
rect 12348 19108 12400 19160
rect 11704 19040 11756 19092
rect 22100 19151 22152 19160
rect 12992 19040 13044 19092
rect 14096 19040 14148 19092
rect 15384 19040 15436 19092
rect 12440 19015 12492 19024
rect 12440 18981 12449 19015
rect 12449 18981 12483 19015
rect 12483 18981 12492 19015
rect 12440 18972 12492 18981
rect 15660 19015 15712 19024
rect 15660 18981 15669 19015
rect 15669 18981 15703 19015
rect 15703 18981 15712 19015
rect 15660 18972 15712 18981
rect 18052 18972 18104 19024
rect 22100 19117 22109 19151
rect 22109 19117 22143 19151
rect 22143 19117 22152 19151
rect 22100 19108 22152 19117
rect 24124 19151 24176 19160
rect 24124 19117 24133 19151
rect 24133 19117 24167 19151
rect 24167 19117 24176 19151
rect 24124 19108 24176 19117
rect 20996 19040 21048 19092
rect 22100 18972 22152 19024
rect 13452 18947 13504 18956
rect 13452 18913 13461 18947
rect 13461 18913 13495 18947
rect 13495 18913 13504 18947
rect 13452 18904 13504 18913
rect 12256 18836 12308 18888
rect 13636 18879 13688 18888
rect 13636 18845 13645 18879
rect 13645 18845 13679 18879
rect 13679 18845 13688 18879
rect 13636 18836 13688 18845
rect 13728 18836 13780 18888
rect 14648 18836 14700 18888
rect 15568 18836 15620 18888
rect 15752 18879 15804 18888
rect 15752 18845 15761 18879
rect 15761 18845 15795 18879
rect 15795 18845 15804 18879
rect 15752 18836 15804 18845
rect 20720 18879 20772 18888
rect 20720 18845 20729 18879
rect 20729 18845 20763 18879
rect 20763 18845 20772 18879
rect 20720 18836 20772 18845
rect 21272 18879 21324 18888
rect 21272 18845 21281 18879
rect 21281 18845 21315 18879
rect 21315 18845 21324 18879
rect 21272 18836 21324 18845
rect 21456 18836 21508 18888
rect 22652 19040 22704 19092
rect 22560 18972 22612 19024
rect 25504 19015 25556 19024
rect 25504 18981 25513 19015
rect 25513 18981 25547 19015
rect 25547 18981 25556 19015
rect 25504 18972 25556 18981
rect 25136 18879 25188 18888
rect 25136 18845 25145 18879
rect 25145 18845 25179 18879
rect 25179 18845 25188 18879
rect 25136 18836 25188 18845
rect 10315 18734 10367 18786
rect 10379 18734 10431 18786
rect 10443 18734 10495 18786
rect 10507 18734 10559 18786
rect 19648 18734 19700 18786
rect 19712 18734 19764 18786
rect 19776 18734 19828 18786
rect 19840 18734 19892 18786
rect 12348 18632 12400 18684
rect 13728 18675 13780 18684
rect 13728 18641 13737 18675
rect 13737 18641 13771 18675
rect 13771 18641 13780 18675
rect 13728 18632 13780 18641
rect 14096 18675 14148 18684
rect 14096 18641 14105 18675
rect 14105 18641 14139 18675
rect 14139 18641 14148 18675
rect 14096 18632 14148 18641
rect 15384 18675 15436 18684
rect 15384 18641 15393 18675
rect 15393 18641 15427 18675
rect 15427 18641 15436 18675
rect 15384 18632 15436 18641
rect 15752 18675 15804 18684
rect 15752 18641 15761 18675
rect 15761 18641 15795 18675
rect 15795 18641 15804 18675
rect 15752 18632 15804 18641
rect 20996 18632 21048 18684
rect 22560 18632 22612 18684
rect 24032 18632 24084 18684
rect 16856 18564 16908 18616
rect 24124 18564 24176 18616
rect 17592 18496 17644 18548
rect 16396 18428 16448 18480
rect 18052 18471 18104 18480
rect 18052 18437 18061 18471
rect 18061 18437 18095 18471
rect 18095 18437 18104 18471
rect 18052 18428 18104 18437
rect 20536 18428 20588 18480
rect 20904 18428 20956 18480
rect 21456 18496 21508 18548
rect 22192 18496 22244 18548
rect 23664 18496 23716 18548
rect 25136 18428 25188 18480
rect 16120 18335 16172 18344
rect 16120 18301 16129 18335
rect 16129 18301 16163 18335
rect 16163 18301 16172 18335
rect 16120 18292 16172 18301
rect 16488 18292 16540 18344
rect 19432 18335 19484 18344
rect 19432 18301 19441 18335
rect 19441 18301 19475 18335
rect 19475 18301 19484 18335
rect 19432 18292 19484 18301
rect 21364 18292 21416 18344
rect 5648 18190 5700 18242
rect 5712 18190 5764 18242
rect 5776 18190 5828 18242
rect 5840 18190 5892 18242
rect 14982 18190 15034 18242
rect 15046 18190 15098 18242
rect 15110 18190 15162 18242
rect 15174 18190 15226 18242
rect 24315 18190 24367 18242
rect 24379 18190 24431 18242
rect 24443 18190 24495 18242
rect 24507 18190 24559 18242
rect 15384 18131 15436 18140
rect 15384 18097 15393 18131
rect 15393 18097 15427 18131
rect 15427 18097 15436 18131
rect 15384 18088 15436 18097
rect 16856 18131 16908 18140
rect 16856 18097 16865 18131
rect 16865 18097 16899 18131
rect 16899 18097 16908 18131
rect 16856 18088 16908 18097
rect 17132 18088 17184 18140
rect 17592 18131 17644 18140
rect 17592 18097 17601 18131
rect 17601 18097 17635 18131
rect 17635 18097 17644 18131
rect 17592 18088 17644 18097
rect 22192 18088 22244 18140
rect 22376 18088 22428 18140
rect 23664 18088 23716 18140
rect 25320 18131 25372 18140
rect 25320 18097 25329 18131
rect 25329 18097 25363 18131
rect 25363 18097 25372 18131
rect 25320 18088 25372 18097
rect 15936 17995 15988 18004
rect 15936 17961 15945 17995
rect 15945 17961 15979 17995
rect 15979 17961 15988 17995
rect 15936 17952 15988 17961
rect 16396 17927 16448 17936
rect 16396 17893 16405 17927
rect 16405 17893 16439 17927
rect 16439 17893 16448 17927
rect 16396 17884 16448 17893
rect 16120 17816 16172 17868
rect 15292 17748 15344 17800
rect 18144 17748 18196 17800
rect 20904 17927 20956 17936
rect 18604 17816 18656 17868
rect 19432 17816 19484 17868
rect 20904 17893 20913 17927
rect 20913 17893 20947 17927
rect 20947 17893 20956 17927
rect 20904 17884 20956 17893
rect 20996 17884 21048 17936
rect 25136 17927 25188 17936
rect 25136 17893 25145 17927
rect 25145 17893 25179 17927
rect 25179 17893 25188 17927
rect 25136 17884 25188 17893
rect 24124 17859 24176 17868
rect 24124 17825 24133 17859
rect 24133 17825 24167 17859
rect 24167 17825 24176 17859
rect 24124 17816 24176 17825
rect 19984 17748 20036 17800
rect 20720 17791 20772 17800
rect 20720 17757 20729 17791
rect 20729 17757 20763 17791
rect 20763 17757 20772 17791
rect 20720 17748 20772 17757
rect 23664 17791 23716 17800
rect 23664 17757 23673 17791
rect 23673 17757 23707 17791
rect 23707 17757 23716 17791
rect 23664 17748 23716 17757
rect 10315 17646 10367 17698
rect 10379 17646 10431 17698
rect 10443 17646 10495 17698
rect 10507 17646 10559 17698
rect 19648 17646 19700 17698
rect 19712 17646 19764 17698
rect 19776 17646 19828 17698
rect 19840 17646 19892 17698
rect 14648 17544 14700 17596
rect 17132 17587 17184 17596
rect 17132 17553 17141 17587
rect 17141 17553 17175 17587
rect 17175 17553 17184 17587
rect 17132 17544 17184 17553
rect 18512 17587 18564 17596
rect 18512 17553 18521 17587
rect 18521 17553 18555 17587
rect 18555 17553 18564 17587
rect 18512 17544 18564 17553
rect 20996 17587 21048 17596
rect 20996 17553 21005 17587
rect 21005 17553 21039 17587
rect 21039 17553 21048 17587
rect 20996 17544 21048 17553
rect 21824 17587 21876 17596
rect 21824 17553 21833 17587
rect 21833 17553 21867 17587
rect 21867 17553 21876 17587
rect 21824 17544 21876 17553
rect 22100 17544 22152 17596
rect 24768 17587 24820 17596
rect 24768 17553 24777 17587
rect 24777 17553 24811 17587
rect 24811 17553 24820 17587
rect 24768 17544 24820 17553
rect 14740 17476 14792 17528
rect 15936 17476 15988 17528
rect 14188 17408 14240 17460
rect 15752 17451 15804 17460
rect 15752 17417 15761 17451
rect 15761 17417 15795 17451
rect 15795 17417 15804 17451
rect 15752 17408 15804 17417
rect 18052 17408 18104 17460
rect 18420 17451 18472 17460
rect 18420 17417 18429 17451
rect 18429 17417 18463 17451
rect 18463 17417 18472 17451
rect 18420 17408 18472 17417
rect 19340 17408 19392 17460
rect 20720 17476 20772 17528
rect 19892 17451 19944 17460
rect 19892 17417 19926 17451
rect 19926 17417 19944 17451
rect 19892 17408 19944 17417
rect 22192 17451 22244 17460
rect 22192 17417 22201 17451
rect 22201 17417 22235 17451
rect 22235 17417 22244 17451
rect 22192 17408 22244 17417
rect 24124 17408 24176 17460
rect 25044 17408 25096 17460
rect 14740 17383 14792 17392
rect 14740 17349 14749 17383
rect 14749 17349 14783 17383
rect 14783 17349 14792 17383
rect 14740 17340 14792 17349
rect 18604 17383 18656 17392
rect 18604 17349 18613 17383
rect 18613 17349 18647 17383
rect 18647 17349 18656 17383
rect 19432 17383 19484 17392
rect 18604 17340 18656 17349
rect 19432 17349 19441 17383
rect 19441 17349 19475 17383
rect 19475 17349 19484 17383
rect 19432 17340 19484 17349
rect 22376 17383 22428 17392
rect 22376 17349 22385 17383
rect 22385 17349 22419 17383
rect 22419 17349 22428 17383
rect 22376 17340 22428 17349
rect 14004 17204 14056 17256
rect 15384 17247 15436 17256
rect 15384 17213 15393 17247
rect 15393 17213 15427 17247
rect 15427 17213 15436 17247
rect 15384 17204 15436 17213
rect 18880 17204 18932 17256
rect 19064 17247 19116 17256
rect 19064 17213 19073 17247
rect 19073 17213 19107 17247
rect 19107 17213 19116 17247
rect 19064 17204 19116 17213
rect 5648 17102 5700 17154
rect 5712 17102 5764 17154
rect 5776 17102 5828 17154
rect 5840 17102 5892 17154
rect 14982 17102 15034 17154
rect 15046 17102 15098 17154
rect 15110 17102 15162 17154
rect 15174 17102 15226 17154
rect 24315 17102 24367 17154
rect 24379 17102 24431 17154
rect 24443 17102 24495 17154
rect 24507 17102 24559 17154
rect 14832 17000 14884 17052
rect 15936 17000 15988 17052
rect 16304 17000 16356 17052
rect 18604 17000 18656 17052
rect 19340 17000 19392 17052
rect 20536 17000 20588 17052
rect 22192 17000 22244 17052
rect 25044 17043 25096 17052
rect 25044 17009 25053 17043
rect 25053 17009 25087 17043
rect 25087 17009 25096 17043
rect 25044 17000 25096 17009
rect 25412 17043 25464 17052
rect 25412 17009 25421 17043
rect 25421 17009 25455 17043
rect 25455 17009 25464 17043
rect 25412 17000 25464 17009
rect 18052 16975 18104 16984
rect 18052 16941 18061 16975
rect 18061 16941 18095 16975
rect 18095 16941 18104 16975
rect 18052 16932 18104 16941
rect 18420 16907 18472 16916
rect 18420 16873 18429 16907
rect 18429 16873 18463 16907
rect 18463 16873 18472 16907
rect 18420 16864 18472 16873
rect 22100 16932 22152 16984
rect 22284 16864 22336 16916
rect 14188 16839 14240 16848
rect 14188 16805 14197 16839
rect 14197 16805 14231 16839
rect 14231 16805 14240 16839
rect 14188 16796 14240 16805
rect 15384 16796 15436 16848
rect 19064 16796 19116 16848
rect 23940 16839 23992 16848
rect 23940 16805 23949 16839
rect 23949 16805 23983 16839
rect 23983 16805 23992 16839
rect 23940 16796 23992 16805
rect 14740 16728 14792 16780
rect 18420 16728 18472 16780
rect 19340 16728 19392 16780
rect 19892 16728 19944 16780
rect 21732 16728 21784 16780
rect 23664 16728 23716 16780
rect 14648 16703 14700 16712
rect 14648 16669 14657 16703
rect 14657 16669 14691 16703
rect 14691 16669 14700 16703
rect 14648 16660 14700 16669
rect 18604 16703 18656 16712
rect 18604 16669 18613 16703
rect 18613 16669 18647 16703
rect 18647 16669 18656 16703
rect 18604 16660 18656 16669
rect 19064 16703 19116 16712
rect 19064 16669 19073 16703
rect 19073 16669 19107 16703
rect 19107 16669 19116 16703
rect 19064 16660 19116 16669
rect 21916 16703 21968 16712
rect 21916 16669 21925 16703
rect 21925 16669 21959 16703
rect 21959 16669 21968 16703
rect 21916 16660 21968 16669
rect 22376 16703 22428 16712
rect 22376 16669 22385 16703
rect 22385 16669 22419 16703
rect 22419 16669 22428 16703
rect 22376 16660 22428 16669
rect 10315 16558 10367 16610
rect 10379 16558 10431 16610
rect 10443 16558 10495 16610
rect 10507 16558 10559 16610
rect 19648 16558 19700 16610
rect 19712 16558 19764 16610
rect 19776 16558 19828 16610
rect 19840 16558 19892 16610
rect 15384 16456 15436 16508
rect 15844 16456 15896 16508
rect 16304 16499 16356 16508
rect 16304 16465 16313 16499
rect 16313 16465 16347 16499
rect 16347 16465 16356 16499
rect 16304 16456 16356 16465
rect 18512 16456 18564 16508
rect 18696 16499 18748 16508
rect 18696 16465 18705 16499
rect 18705 16465 18739 16499
rect 18739 16465 18748 16499
rect 18696 16456 18748 16465
rect 18880 16456 18932 16508
rect 19432 16456 19484 16508
rect 22376 16456 22428 16508
rect 25412 16499 25464 16508
rect 25412 16465 25421 16499
rect 25421 16465 25455 16499
rect 25455 16465 25464 16499
rect 25412 16456 25464 16465
rect 14740 16388 14792 16440
rect 21180 16431 21232 16440
rect 21180 16397 21189 16431
rect 21189 16397 21223 16431
rect 21223 16397 21232 16431
rect 21180 16388 21232 16397
rect 22468 16388 22520 16440
rect 15752 16320 15804 16372
rect 18604 16320 18656 16372
rect 21548 16320 21600 16372
rect 22560 16363 22612 16372
rect 22560 16329 22569 16363
rect 22569 16329 22603 16363
rect 22603 16329 22612 16363
rect 22560 16320 22612 16329
rect 23756 16320 23808 16372
rect 25228 16363 25280 16372
rect 25228 16329 25237 16363
rect 25237 16329 25271 16363
rect 25271 16329 25280 16363
rect 25228 16320 25280 16329
rect 14280 16295 14332 16304
rect 14280 16261 14289 16295
rect 14289 16261 14323 16295
rect 14323 16261 14332 16295
rect 14280 16252 14332 16261
rect 16488 16295 16540 16304
rect 16488 16261 16497 16295
rect 16497 16261 16531 16295
rect 16531 16261 16540 16295
rect 16488 16252 16540 16261
rect 18788 16184 18840 16236
rect 19340 16252 19392 16304
rect 21272 16295 21324 16304
rect 21272 16261 21281 16295
rect 21281 16261 21315 16295
rect 21315 16261 21324 16295
rect 22284 16295 22336 16304
rect 21272 16252 21324 16261
rect 22284 16261 22293 16295
rect 22293 16261 22327 16295
rect 22327 16261 22336 16295
rect 22284 16252 22336 16261
rect 23572 16252 23624 16304
rect 24124 16252 24176 16304
rect 23480 16184 23532 16236
rect 23940 16184 23992 16236
rect 5648 16014 5700 16066
rect 5712 16014 5764 16066
rect 5776 16014 5828 16066
rect 5840 16014 5892 16066
rect 14982 16014 15034 16066
rect 15046 16014 15098 16066
rect 15110 16014 15162 16066
rect 15174 16014 15226 16066
rect 24315 16014 24367 16066
rect 24379 16014 24431 16066
rect 24443 16014 24495 16066
rect 24507 16014 24559 16066
rect 14004 15955 14056 15964
rect 14004 15921 14013 15955
rect 14013 15921 14047 15955
rect 14047 15921 14056 15955
rect 14004 15912 14056 15921
rect 15292 15955 15344 15964
rect 15292 15921 15301 15955
rect 15301 15921 15335 15955
rect 15335 15921 15344 15955
rect 15292 15912 15344 15921
rect 16488 15912 16540 15964
rect 19432 15912 19484 15964
rect 21180 15955 21232 15964
rect 21180 15921 21189 15955
rect 21189 15921 21223 15955
rect 21223 15921 21232 15955
rect 21180 15912 21232 15921
rect 23756 15912 23808 15964
rect 24768 15955 24820 15964
rect 24768 15921 24777 15955
rect 24777 15921 24811 15955
rect 24811 15921 24820 15955
rect 24768 15912 24820 15921
rect 25228 15912 25280 15964
rect 16120 15844 16172 15896
rect 15844 15819 15896 15828
rect 15844 15785 15853 15819
rect 15853 15785 15887 15819
rect 15887 15785 15896 15819
rect 15844 15776 15896 15785
rect 19248 15776 19300 15828
rect 20720 15776 20772 15828
rect 16488 15708 16540 15760
rect 17868 15708 17920 15760
rect 22284 15708 22336 15760
rect 24676 15708 24728 15760
rect 18880 15640 18932 15692
rect 20352 15640 20404 15692
rect 21272 15640 21324 15692
rect 21732 15640 21784 15692
rect 13636 15572 13688 15624
rect 14280 15615 14332 15624
rect 14280 15581 14289 15615
rect 14289 15581 14323 15615
rect 14323 15581 14332 15615
rect 14280 15572 14332 15581
rect 14740 15615 14792 15624
rect 14740 15581 14749 15615
rect 14749 15581 14783 15615
rect 14783 15581 14792 15615
rect 14740 15572 14792 15581
rect 15660 15615 15712 15624
rect 15660 15581 15669 15615
rect 15669 15581 15703 15615
rect 15703 15581 15712 15615
rect 15660 15572 15712 15581
rect 18696 15572 18748 15624
rect 18972 15615 19024 15624
rect 18972 15581 18981 15615
rect 18981 15581 19015 15615
rect 19015 15581 19024 15615
rect 18972 15572 19024 15581
rect 21548 15615 21600 15624
rect 21548 15581 21557 15615
rect 21557 15581 21591 15615
rect 21591 15581 21600 15615
rect 21548 15572 21600 15581
rect 23664 15572 23716 15624
rect 10315 15470 10367 15522
rect 10379 15470 10431 15522
rect 10443 15470 10495 15522
rect 10507 15470 10559 15522
rect 19648 15470 19700 15522
rect 19712 15470 19764 15522
rect 19776 15470 19828 15522
rect 19840 15470 19892 15522
rect 14740 15368 14792 15420
rect 15844 15368 15896 15420
rect 16396 15411 16448 15420
rect 16396 15377 16405 15411
rect 16405 15377 16439 15411
rect 16439 15377 16448 15411
rect 16396 15368 16448 15377
rect 18604 15368 18656 15420
rect 18788 15411 18840 15420
rect 18788 15377 18797 15411
rect 18797 15377 18831 15411
rect 18831 15377 18840 15411
rect 18788 15368 18840 15377
rect 20352 15411 20404 15420
rect 20352 15377 20361 15411
rect 20361 15377 20395 15411
rect 20395 15377 20404 15411
rect 20352 15368 20404 15377
rect 22284 15368 22336 15420
rect 23020 15368 23072 15420
rect 24032 15368 24084 15420
rect 24860 15368 24912 15420
rect 25596 15368 25648 15420
rect 19248 15343 19300 15352
rect 19248 15309 19282 15343
rect 19282 15309 19300 15343
rect 19248 15300 19300 15309
rect 13912 15275 13964 15284
rect 13912 15241 13946 15275
rect 13946 15241 13964 15275
rect 13912 15232 13964 15241
rect 15292 15232 15344 15284
rect 16304 15275 16356 15284
rect 16304 15241 16313 15275
rect 16313 15241 16347 15275
rect 16347 15241 16356 15275
rect 16304 15232 16356 15241
rect 20720 15232 20772 15284
rect 21272 15232 21324 15284
rect 21732 15232 21784 15284
rect 23480 15232 23532 15284
rect 25872 15232 25924 15284
rect 13636 15207 13688 15216
rect 13636 15173 13645 15207
rect 13645 15173 13679 15207
rect 13679 15173 13688 15207
rect 13636 15164 13688 15173
rect 18788 15164 18840 15216
rect 23664 15164 23716 15216
rect 24124 15164 24176 15216
rect 16856 15096 16908 15148
rect 15936 15071 15988 15080
rect 15936 15037 15945 15071
rect 15945 15037 15979 15071
rect 15979 15037 15988 15071
rect 15936 15028 15988 15037
rect 23664 15071 23716 15080
rect 23664 15037 23673 15071
rect 23673 15037 23707 15071
rect 23707 15037 23716 15071
rect 23664 15028 23716 15037
rect 5648 14926 5700 14978
rect 5712 14926 5764 14978
rect 5776 14926 5828 14978
rect 5840 14926 5892 14978
rect 14982 14926 15034 14978
rect 15046 14926 15098 14978
rect 15110 14926 15162 14978
rect 15174 14926 15226 14978
rect 24315 14926 24367 14978
rect 24379 14926 24431 14978
rect 24443 14926 24495 14978
rect 24507 14926 24559 14978
rect 13912 14824 13964 14876
rect 14648 14824 14700 14876
rect 15292 14824 15344 14876
rect 15476 14867 15528 14876
rect 15476 14833 15485 14867
rect 15485 14833 15519 14867
rect 15519 14833 15528 14867
rect 15476 14824 15528 14833
rect 16396 14824 16448 14876
rect 18880 14867 18932 14876
rect 18880 14833 18889 14867
rect 18889 14833 18923 14867
rect 18923 14833 18932 14867
rect 18880 14824 18932 14833
rect 19340 14824 19392 14876
rect 21272 14824 21324 14876
rect 21732 14867 21784 14876
rect 21732 14833 21741 14867
rect 21741 14833 21775 14867
rect 21775 14833 21784 14867
rect 21732 14824 21784 14833
rect 24124 14824 24176 14876
rect 24860 14867 24912 14876
rect 24860 14833 24869 14867
rect 24869 14833 24903 14867
rect 24903 14833 24912 14867
rect 24860 14824 24912 14833
rect 25504 14867 25556 14876
rect 25504 14833 25513 14867
rect 25513 14833 25547 14867
rect 25547 14833 25556 14867
rect 25504 14824 25556 14833
rect 25872 14867 25924 14876
rect 25872 14833 25881 14867
rect 25881 14833 25915 14867
rect 25915 14833 25924 14867
rect 25872 14824 25924 14833
rect 15752 14756 15804 14808
rect 23480 14756 23532 14808
rect 19064 14688 19116 14740
rect 19524 14731 19576 14740
rect 19524 14697 19533 14731
rect 19533 14697 19567 14731
rect 19567 14697 19576 14731
rect 19524 14688 19576 14697
rect 20720 14731 20772 14740
rect 20720 14697 20729 14731
rect 20729 14697 20763 14731
rect 20763 14697 20772 14731
rect 20720 14688 20772 14697
rect 23020 14731 23072 14740
rect 23020 14697 23029 14731
rect 23029 14697 23063 14731
rect 23063 14697 23072 14731
rect 23020 14688 23072 14697
rect 24676 14688 24728 14740
rect 15384 14620 15436 14672
rect 22560 14620 22612 14672
rect 23664 14620 23716 14672
rect 24584 14620 24636 14672
rect 16856 14552 16908 14604
rect 18144 14552 18196 14604
rect 18788 14552 18840 14604
rect 13636 14527 13688 14536
rect 13636 14493 13645 14527
rect 13645 14493 13679 14527
rect 13679 14493 13688 14527
rect 13636 14484 13688 14493
rect 18052 14527 18104 14536
rect 18052 14493 18061 14527
rect 18061 14493 18095 14527
rect 18095 14493 18104 14527
rect 18052 14484 18104 14493
rect 18420 14527 18472 14536
rect 18420 14493 18429 14527
rect 18429 14493 18463 14527
rect 18463 14493 18472 14527
rect 19248 14527 19300 14536
rect 18420 14484 18472 14493
rect 19248 14493 19257 14527
rect 19257 14493 19291 14527
rect 19291 14493 19300 14527
rect 19248 14484 19300 14493
rect 20904 14527 20956 14536
rect 20904 14493 20913 14527
rect 20913 14493 20947 14527
rect 20947 14493 20956 14527
rect 20904 14484 20956 14493
rect 22192 14484 22244 14536
rect 22928 14527 22980 14536
rect 22928 14493 22937 14527
rect 22937 14493 22971 14527
rect 22971 14493 22980 14527
rect 22928 14484 22980 14493
rect 25044 14484 25096 14536
rect 10315 14382 10367 14434
rect 10379 14382 10431 14434
rect 10443 14382 10495 14434
rect 10507 14382 10559 14434
rect 19648 14382 19700 14434
rect 19712 14382 19764 14434
rect 19776 14382 19828 14434
rect 19840 14382 19892 14434
rect 13544 14280 13596 14332
rect 16856 14280 16908 14332
rect 19340 14280 19392 14332
rect 22560 14323 22612 14332
rect 22560 14289 22569 14323
rect 22569 14289 22603 14323
rect 22603 14289 22612 14323
rect 22560 14280 22612 14289
rect 23020 14280 23072 14332
rect 23480 14323 23532 14332
rect 23480 14289 23489 14323
rect 23489 14289 23523 14323
rect 23523 14289 23532 14323
rect 23480 14280 23532 14289
rect 24584 14323 24636 14332
rect 24584 14289 24593 14323
rect 24593 14289 24627 14323
rect 24627 14289 24636 14323
rect 24584 14280 24636 14289
rect 25136 14280 25188 14332
rect 15752 14212 15804 14264
rect 21088 14255 21140 14264
rect 21088 14221 21097 14255
rect 21097 14221 21131 14255
rect 21131 14221 21140 14255
rect 21088 14212 21140 14221
rect 25044 14212 25096 14264
rect 13452 14187 13504 14196
rect 13452 14153 13461 14187
rect 13461 14153 13495 14187
rect 13495 14153 13504 14187
rect 13452 14144 13504 14153
rect 16396 14144 16448 14196
rect 18052 14144 18104 14196
rect 19524 14144 19576 14196
rect 20812 14187 20864 14196
rect 20812 14153 20821 14187
rect 20821 14153 20855 14187
rect 20855 14153 20864 14187
rect 20812 14144 20864 14153
rect 23664 14144 23716 14196
rect 25596 14144 25648 14196
rect 18144 14076 18196 14128
rect 15384 13983 15436 13992
rect 15384 13949 15393 13983
rect 15393 13949 15427 13983
rect 15427 13949 15436 13983
rect 15384 13940 15436 13949
rect 5648 13838 5700 13890
rect 5712 13838 5764 13890
rect 5776 13838 5828 13890
rect 5840 13838 5892 13890
rect 14982 13838 15034 13890
rect 15046 13838 15098 13890
rect 15110 13838 15162 13890
rect 15174 13838 15226 13890
rect 24315 13838 24367 13890
rect 24379 13838 24431 13890
rect 24443 13838 24495 13890
rect 24507 13838 24559 13890
rect 13452 13779 13504 13788
rect 13452 13745 13461 13779
rect 13461 13745 13495 13779
rect 13495 13745 13504 13779
rect 13452 13736 13504 13745
rect 15752 13736 15804 13788
rect 15936 13736 15988 13788
rect 16396 13779 16448 13788
rect 16396 13745 16405 13779
rect 16405 13745 16439 13779
rect 16439 13745 16448 13779
rect 16396 13736 16448 13745
rect 16948 13736 17000 13788
rect 18052 13736 18104 13788
rect 18972 13736 19024 13788
rect 19524 13779 19576 13788
rect 19524 13745 19533 13779
rect 19533 13745 19567 13779
rect 19567 13745 19576 13779
rect 19524 13736 19576 13745
rect 20260 13779 20312 13788
rect 20260 13745 20269 13779
rect 20269 13745 20303 13779
rect 20303 13745 20312 13779
rect 20260 13736 20312 13745
rect 17960 13711 18012 13720
rect 17960 13677 17969 13711
rect 17969 13677 18003 13711
rect 18003 13677 18012 13711
rect 17960 13668 18012 13677
rect 15384 13600 15436 13652
rect 20812 13668 20864 13720
rect 23664 13736 23716 13788
rect 23940 13736 23992 13788
rect 25596 13779 25648 13788
rect 25596 13745 25605 13779
rect 25605 13745 25639 13779
rect 25639 13745 25648 13779
rect 25596 13736 25648 13745
rect 22100 13600 22152 13652
rect 25228 13643 25280 13652
rect 25228 13609 25237 13643
rect 25237 13609 25271 13643
rect 25271 13609 25280 13643
rect 25228 13600 25280 13609
rect 15292 13575 15344 13584
rect 15292 13541 15301 13575
rect 15301 13541 15335 13575
rect 15335 13541 15344 13575
rect 15292 13532 15344 13541
rect 16948 13532 17000 13584
rect 18144 13532 18196 13584
rect 20812 13532 20864 13584
rect 18880 13507 18932 13516
rect 18880 13473 18889 13507
rect 18889 13473 18923 13507
rect 18923 13473 18932 13507
rect 18880 13464 18932 13473
rect 21824 13464 21876 13516
rect 13176 13396 13228 13448
rect 10315 13294 10367 13346
rect 10379 13294 10431 13346
rect 10443 13294 10495 13346
rect 10507 13294 10559 13346
rect 19648 13294 19700 13346
rect 19712 13294 19764 13346
rect 19776 13294 19828 13346
rect 19840 13294 19892 13346
rect 18880 13192 18932 13244
rect 21824 13235 21876 13244
rect 21824 13201 21833 13235
rect 21833 13201 21867 13235
rect 21867 13201 21876 13235
rect 21824 13192 21876 13201
rect 23848 13192 23900 13244
rect 16948 13167 17000 13176
rect 16948 13133 16957 13167
rect 16957 13133 16991 13167
rect 16991 13133 17000 13167
rect 16948 13124 17000 13133
rect 21272 13124 21324 13176
rect 16672 13099 16724 13108
rect 16672 13065 16681 13099
rect 16681 13065 16715 13099
rect 16715 13065 16724 13099
rect 16672 13056 16724 13065
rect 19616 13099 19668 13108
rect 19616 13065 19625 13099
rect 19625 13065 19659 13099
rect 19659 13065 19668 13099
rect 19616 13056 19668 13065
rect 19892 13099 19944 13108
rect 19892 13065 19926 13099
rect 19926 13065 19944 13099
rect 19892 13056 19944 13065
rect 25044 13056 25096 13108
rect 12992 12988 13044 13040
rect 18052 12988 18104 13040
rect 13268 12895 13320 12904
rect 13268 12861 13277 12895
rect 13277 12861 13311 12895
rect 13311 12861 13320 12895
rect 13268 12852 13320 12861
rect 15844 12852 15896 12904
rect 21364 12895 21416 12904
rect 21364 12861 21373 12895
rect 21373 12861 21407 12895
rect 21407 12861 21416 12895
rect 21364 12852 21416 12861
rect 5648 12750 5700 12802
rect 5712 12750 5764 12802
rect 5776 12750 5828 12802
rect 5840 12750 5892 12802
rect 14982 12750 15034 12802
rect 15046 12750 15098 12802
rect 15110 12750 15162 12802
rect 15174 12750 15226 12802
rect 24315 12750 24367 12802
rect 24379 12750 24431 12802
rect 24443 12750 24495 12802
rect 24507 12750 24559 12802
rect 12992 12691 13044 12700
rect 12992 12657 13001 12691
rect 13001 12657 13035 12691
rect 13035 12657 13044 12691
rect 12992 12648 13044 12657
rect 13176 12691 13228 12700
rect 13176 12657 13185 12691
rect 13185 12657 13219 12691
rect 13219 12657 13228 12691
rect 13176 12648 13228 12657
rect 15292 12691 15344 12700
rect 15292 12657 15301 12691
rect 15301 12657 15335 12691
rect 15335 12657 15344 12691
rect 15292 12648 15344 12657
rect 18052 12691 18104 12700
rect 18052 12657 18061 12691
rect 18061 12657 18095 12691
rect 18095 12657 18104 12691
rect 18052 12648 18104 12657
rect 19616 12691 19668 12700
rect 19616 12657 19625 12691
rect 19625 12657 19659 12691
rect 19659 12657 19668 12691
rect 19616 12648 19668 12657
rect 16672 12580 16724 12632
rect 13268 12512 13320 12564
rect 15844 12555 15896 12564
rect 15844 12521 15853 12555
rect 15853 12521 15887 12555
rect 15887 12521 15896 12555
rect 15844 12512 15896 12521
rect 16488 12512 16540 12564
rect 18604 12555 18656 12564
rect 18604 12521 18613 12555
rect 18613 12521 18647 12555
rect 18647 12521 18656 12555
rect 18604 12512 18656 12521
rect 22100 12648 22152 12700
rect 24216 12691 24268 12700
rect 24216 12657 24225 12691
rect 24225 12657 24259 12691
rect 24259 12657 24268 12691
rect 24216 12648 24268 12657
rect 25044 12691 25096 12700
rect 25044 12657 25053 12691
rect 25053 12657 25087 12691
rect 25087 12657 25096 12691
rect 25044 12648 25096 12657
rect 24676 12555 24728 12564
rect 18052 12444 18104 12496
rect 13084 12376 13136 12428
rect 15384 12376 15436 12428
rect 15568 12308 15620 12360
rect 19524 12444 19576 12496
rect 19892 12444 19944 12496
rect 24676 12521 24685 12555
rect 24685 12521 24719 12555
rect 24719 12521 24728 12555
rect 24676 12512 24728 12521
rect 21364 12376 21416 12428
rect 10315 12206 10367 12258
rect 10379 12206 10431 12258
rect 10443 12206 10495 12258
rect 10507 12206 10559 12258
rect 19648 12206 19700 12258
rect 19712 12206 19764 12258
rect 19776 12206 19828 12258
rect 19840 12206 19892 12258
rect 16488 12104 16540 12156
rect 16764 12104 16816 12156
rect 19524 12147 19576 12156
rect 19524 12113 19533 12147
rect 19533 12113 19567 12147
rect 19567 12113 19576 12147
rect 19524 12104 19576 12113
rect 20812 12147 20864 12156
rect 20812 12113 20821 12147
rect 20821 12113 20855 12147
rect 20855 12113 20864 12147
rect 20812 12104 20864 12113
rect 24032 12104 24084 12156
rect 13268 12079 13320 12088
rect 13268 12045 13302 12079
rect 13302 12045 13320 12079
rect 13268 12036 13320 12045
rect 13636 12036 13688 12088
rect 12532 11968 12584 12020
rect 15936 12036 15988 12088
rect 15292 11968 15344 12020
rect 18052 11968 18104 12020
rect 21180 12011 21232 12020
rect 21180 11977 21189 12011
rect 21189 11977 21223 12011
rect 21223 11977 21232 12011
rect 21180 11968 21232 11977
rect 21456 11968 21508 12020
rect 24584 12011 24636 12020
rect 24584 11977 24593 12011
rect 24593 11977 24627 12011
rect 24627 11977 24636 12011
rect 24584 11968 24636 11977
rect 18144 11943 18196 11952
rect 18144 11909 18153 11943
rect 18153 11909 18187 11943
rect 18187 11909 18196 11943
rect 18144 11900 18196 11909
rect 21364 11943 21416 11952
rect 21364 11909 21373 11943
rect 21373 11909 21407 11943
rect 21407 11909 21416 11943
rect 21364 11900 21416 11909
rect 14372 11807 14424 11816
rect 14372 11773 14381 11807
rect 14381 11773 14415 11807
rect 14415 11773 14424 11807
rect 14372 11764 14424 11773
rect 5648 11662 5700 11714
rect 5712 11662 5764 11714
rect 5776 11662 5828 11714
rect 5840 11662 5892 11714
rect 14982 11662 15034 11714
rect 15046 11662 15098 11714
rect 15110 11662 15162 11714
rect 15174 11662 15226 11714
rect 24315 11662 24367 11714
rect 24379 11662 24431 11714
rect 24443 11662 24495 11714
rect 24507 11662 24559 11714
rect 13268 11560 13320 11612
rect 14372 11560 14424 11612
rect 15292 11560 15344 11612
rect 15936 11603 15988 11612
rect 15936 11569 15945 11603
rect 15945 11569 15979 11603
rect 15979 11569 15988 11603
rect 15936 11560 15988 11569
rect 12532 11467 12584 11476
rect 12532 11433 12541 11467
rect 12541 11433 12575 11467
rect 12575 11433 12584 11467
rect 12532 11424 12584 11433
rect 15384 11467 15436 11476
rect 15384 11433 15393 11467
rect 15393 11433 15427 11467
rect 15427 11433 15436 11467
rect 15384 11424 15436 11433
rect 18144 11560 18196 11612
rect 18604 11560 18656 11612
rect 21364 11560 21416 11612
rect 21456 11603 21508 11612
rect 21456 11569 21465 11603
rect 21465 11569 21499 11603
rect 21499 11569 21508 11603
rect 24676 11603 24728 11612
rect 21456 11560 21508 11569
rect 24676 11569 24685 11603
rect 24685 11569 24719 11603
rect 24719 11569 24728 11603
rect 24676 11560 24728 11569
rect 19432 11467 19484 11476
rect 19432 11433 19441 11467
rect 19441 11433 19475 11467
rect 19475 11433 19484 11467
rect 19432 11424 19484 11433
rect 10048 11356 10100 11408
rect 16764 11356 16816 11408
rect 18972 11356 19024 11408
rect 19248 11356 19300 11408
rect 21180 11399 21232 11408
rect 21180 11365 21189 11399
rect 21189 11365 21223 11399
rect 21223 11365 21232 11399
rect 21180 11356 21232 11365
rect 10140 11331 10192 11340
rect 10140 11297 10149 11331
rect 10149 11297 10183 11331
rect 10183 11297 10192 11331
rect 10140 11288 10192 11297
rect 12808 11331 12860 11340
rect 12808 11297 12842 11331
rect 12842 11297 12860 11331
rect 12808 11288 12860 11297
rect 18052 11263 18104 11272
rect 18052 11229 18061 11263
rect 18061 11229 18095 11263
rect 18095 11229 18104 11263
rect 18052 11220 18104 11229
rect 19248 11263 19300 11272
rect 19248 11229 19257 11263
rect 19257 11229 19291 11263
rect 19291 11229 19300 11263
rect 19248 11220 19300 11229
rect 10315 11118 10367 11170
rect 10379 11118 10431 11170
rect 10443 11118 10495 11170
rect 10507 11118 10559 11170
rect 19648 11118 19700 11170
rect 19712 11118 19764 11170
rect 19776 11118 19828 11170
rect 19840 11118 19892 11170
rect 10048 11016 10100 11068
rect 13084 11059 13136 11068
rect 13084 11025 13093 11059
rect 13093 11025 13127 11059
rect 13127 11025 13136 11059
rect 13084 11016 13136 11025
rect 15568 11059 15620 11068
rect 15568 11025 15577 11059
rect 15577 11025 15611 11059
rect 15611 11025 15620 11059
rect 15568 11016 15620 11025
rect 16764 11059 16816 11068
rect 16764 11025 16773 11059
rect 16773 11025 16807 11059
rect 16807 11025 16816 11059
rect 16764 11016 16816 11025
rect 18052 11016 18104 11068
rect 19432 11016 19484 11068
rect 24768 11059 24820 11068
rect 24768 11025 24777 11059
rect 24777 11025 24811 11059
rect 24811 11025 24820 11059
rect 24768 11016 24820 11025
rect 16028 10991 16080 11000
rect 16028 10957 16037 10991
rect 16037 10957 16071 10991
rect 16071 10957 16080 10991
rect 18972 10991 19024 11000
rect 16028 10948 16080 10957
rect 18972 10957 18981 10991
rect 18981 10957 19015 10991
rect 19015 10957 19024 10991
rect 18972 10948 19024 10957
rect 13176 10880 13228 10932
rect 15660 10880 15712 10932
rect 24676 10880 24728 10932
rect 13544 10855 13596 10864
rect 13544 10821 13553 10855
rect 13553 10821 13587 10855
rect 13587 10821 13596 10855
rect 13544 10812 13596 10821
rect 13728 10855 13780 10864
rect 13728 10821 13737 10855
rect 13737 10821 13771 10855
rect 13771 10821 13780 10855
rect 13728 10812 13780 10821
rect 12808 10744 12860 10796
rect 15292 10744 15344 10796
rect 16304 10744 16356 10796
rect 5648 10574 5700 10626
rect 5712 10574 5764 10626
rect 5776 10574 5828 10626
rect 5840 10574 5892 10626
rect 14982 10574 15034 10626
rect 15046 10574 15098 10626
rect 15110 10574 15162 10626
rect 15174 10574 15226 10626
rect 24315 10574 24367 10626
rect 24379 10574 24431 10626
rect 24443 10574 24495 10626
rect 24507 10574 24559 10626
rect 13820 10515 13872 10524
rect 13820 10481 13829 10515
rect 13829 10481 13863 10515
rect 13863 10481 13872 10515
rect 13820 10472 13872 10481
rect 16028 10515 16080 10524
rect 16028 10481 16037 10515
rect 16037 10481 16071 10515
rect 16071 10481 16080 10515
rect 16028 10472 16080 10481
rect 16304 10515 16356 10524
rect 16304 10481 16313 10515
rect 16313 10481 16347 10515
rect 16347 10481 16356 10515
rect 16304 10472 16356 10481
rect 24676 10472 24728 10524
rect 13544 10447 13596 10456
rect 13544 10413 13553 10447
rect 13553 10413 13587 10447
rect 13587 10413 13596 10447
rect 13544 10404 13596 10413
rect 24124 10404 24176 10456
rect 23940 10268 23992 10320
rect 24124 10268 24176 10320
rect 13176 10175 13228 10184
rect 13176 10141 13185 10175
rect 13185 10141 13219 10175
rect 13219 10141 13228 10175
rect 13176 10132 13228 10141
rect 15660 10175 15712 10184
rect 15660 10141 15669 10175
rect 15669 10141 15703 10175
rect 15703 10141 15712 10175
rect 15660 10132 15712 10141
rect 25228 10175 25280 10184
rect 25228 10141 25237 10175
rect 25237 10141 25271 10175
rect 25271 10141 25280 10175
rect 25228 10132 25280 10141
rect 10315 10030 10367 10082
rect 10379 10030 10431 10082
rect 10443 10030 10495 10082
rect 10507 10030 10559 10082
rect 19648 10030 19700 10082
rect 19712 10030 19764 10082
rect 19776 10030 19828 10082
rect 19840 10030 19892 10082
rect 23296 9928 23348 9980
rect 24676 9792 24728 9844
rect 5648 9486 5700 9538
rect 5712 9486 5764 9538
rect 5776 9486 5828 9538
rect 5840 9486 5892 9538
rect 14982 9486 15034 9538
rect 15046 9486 15098 9538
rect 15110 9486 15162 9538
rect 15174 9486 15226 9538
rect 24315 9486 24367 9538
rect 24379 9486 24431 9538
rect 24443 9486 24495 9538
rect 24507 9486 24559 9538
rect 24768 9359 24820 9368
rect 24768 9325 24777 9359
rect 24777 9325 24811 9359
rect 24811 9325 24820 9359
rect 24768 9316 24820 9325
rect 25228 9359 25280 9368
rect 25228 9325 25237 9359
rect 25237 9325 25271 9359
rect 25271 9325 25280 9359
rect 25228 9316 25280 9325
rect 24492 9087 24544 9096
rect 24492 9053 24501 9087
rect 24501 9053 24535 9087
rect 24535 9053 24544 9087
rect 24492 9044 24544 9053
rect 10315 8942 10367 8994
rect 10379 8942 10431 8994
rect 10443 8942 10495 8994
rect 10507 8942 10559 8994
rect 19648 8942 19700 8994
rect 19712 8942 19764 8994
rect 19776 8942 19828 8994
rect 19840 8942 19892 8994
rect 24768 8883 24820 8892
rect 24768 8849 24777 8883
rect 24777 8849 24811 8883
rect 24811 8849 24820 8883
rect 24768 8840 24820 8849
rect 24676 8704 24728 8756
rect 5648 8398 5700 8450
rect 5712 8398 5764 8450
rect 5776 8398 5828 8450
rect 5840 8398 5892 8450
rect 14982 8398 15034 8450
rect 15046 8398 15098 8450
rect 15110 8398 15162 8450
rect 15174 8398 15226 8450
rect 24315 8398 24367 8450
rect 24379 8398 24431 8450
rect 24443 8398 24495 8450
rect 24507 8398 24559 8450
rect 24676 8339 24728 8348
rect 24676 8305 24685 8339
rect 24685 8305 24719 8339
rect 24719 8305 24728 8339
rect 24676 8296 24728 8305
rect 10315 7854 10367 7906
rect 10379 7854 10431 7906
rect 10443 7854 10495 7906
rect 10507 7854 10559 7906
rect 19648 7854 19700 7906
rect 19712 7854 19764 7906
rect 19776 7854 19828 7906
rect 19840 7854 19892 7906
rect 24584 7659 24636 7668
rect 24584 7625 24593 7659
rect 24593 7625 24627 7659
rect 24627 7625 24636 7659
rect 24584 7616 24636 7625
rect 24768 7523 24820 7532
rect 24768 7489 24777 7523
rect 24777 7489 24811 7523
rect 24811 7489 24820 7523
rect 24768 7480 24820 7489
rect 5648 7310 5700 7362
rect 5712 7310 5764 7362
rect 5776 7310 5828 7362
rect 5840 7310 5892 7362
rect 14982 7310 15034 7362
rect 15046 7310 15098 7362
rect 15110 7310 15162 7362
rect 15174 7310 15226 7362
rect 24315 7310 24367 7362
rect 24379 7310 24431 7362
rect 24443 7310 24495 7362
rect 24507 7310 24559 7362
rect 17776 7251 17828 7260
rect 17776 7217 17785 7251
rect 17785 7217 17819 7251
rect 17819 7217 17828 7251
rect 17776 7208 17828 7217
rect 24676 7251 24728 7260
rect 24676 7217 24685 7251
rect 24685 7217 24719 7251
rect 24719 7217 24728 7251
rect 24676 7208 24728 7217
rect 18236 7115 18288 7124
rect 18236 7081 18245 7115
rect 18245 7081 18279 7115
rect 18279 7081 18288 7115
rect 18236 7072 18288 7081
rect 10315 6766 10367 6818
rect 10379 6766 10431 6818
rect 10443 6766 10495 6818
rect 10507 6766 10559 6818
rect 19648 6766 19700 6818
rect 19712 6766 19764 6818
rect 19776 6766 19828 6818
rect 19840 6766 19892 6818
rect 5648 6222 5700 6274
rect 5712 6222 5764 6274
rect 5776 6222 5828 6274
rect 5840 6222 5892 6274
rect 14982 6222 15034 6274
rect 15046 6222 15098 6274
rect 15110 6222 15162 6274
rect 15174 6222 15226 6274
rect 24315 6222 24367 6274
rect 24379 6222 24431 6274
rect 24443 6222 24495 6274
rect 24507 6222 24559 6274
rect 16488 6120 16540 6172
rect 16856 5891 16908 5900
rect 16856 5857 16865 5891
rect 16865 5857 16899 5891
rect 16899 5857 16908 5891
rect 16856 5848 16908 5857
rect 10315 5678 10367 5730
rect 10379 5678 10431 5730
rect 10443 5678 10495 5730
rect 10507 5678 10559 5730
rect 19648 5678 19700 5730
rect 19712 5678 19764 5730
rect 19776 5678 19828 5730
rect 19840 5678 19892 5730
rect 5648 5134 5700 5186
rect 5712 5134 5764 5186
rect 5776 5134 5828 5186
rect 5840 5134 5892 5186
rect 14982 5134 15034 5186
rect 15046 5134 15098 5186
rect 15110 5134 15162 5186
rect 15174 5134 15226 5186
rect 24315 5134 24367 5186
rect 24379 5134 24431 5186
rect 24443 5134 24495 5186
rect 24507 5134 24559 5186
rect 16212 5032 16264 5084
rect 15936 4803 15988 4812
rect 15936 4769 15945 4803
rect 15945 4769 15979 4803
rect 15979 4769 15988 4803
rect 15936 4760 15988 4769
rect 10315 4590 10367 4642
rect 10379 4590 10431 4642
rect 10443 4590 10495 4642
rect 10507 4590 10559 4642
rect 19648 4590 19700 4642
rect 19712 4590 19764 4642
rect 19776 4590 19828 4642
rect 19840 4590 19892 4642
rect 5648 4046 5700 4098
rect 5712 4046 5764 4098
rect 5776 4046 5828 4098
rect 5840 4046 5892 4098
rect 14982 4046 15034 4098
rect 15046 4046 15098 4098
rect 15110 4046 15162 4098
rect 15174 4046 15226 4098
rect 24315 4046 24367 4098
rect 24379 4046 24431 4098
rect 24443 4046 24495 4098
rect 24507 4046 24559 4098
rect 24768 3647 24820 3656
rect 24768 3613 24777 3647
rect 24777 3613 24811 3647
rect 24811 3613 24820 3647
rect 24768 3604 24820 3613
rect 25228 3647 25280 3656
rect 25228 3613 25237 3647
rect 25237 3613 25271 3647
rect 25271 3613 25280 3647
rect 25228 3604 25280 3613
rect 10315 3502 10367 3554
rect 10379 3502 10431 3554
rect 10443 3502 10495 3554
rect 10507 3502 10559 3554
rect 19648 3502 19700 3554
rect 19712 3502 19764 3554
rect 19776 3502 19828 3554
rect 19840 3502 19892 3554
rect 5648 2958 5700 3010
rect 5712 2958 5764 3010
rect 5776 2958 5828 3010
rect 5840 2958 5892 3010
rect 14982 2958 15034 3010
rect 15046 2958 15098 3010
rect 15110 2958 15162 3010
rect 15174 2958 15226 3010
rect 24315 2958 24367 3010
rect 24379 2958 24431 3010
rect 24443 2958 24495 3010
rect 24507 2958 24559 3010
rect 10315 2414 10367 2466
rect 10379 2414 10431 2466
rect 10443 2414 10495 2466
rect 10507 2414 10559 2466
rect 19648 2414 19700 2466
rect 19712 2414 19764 2466
rect 19776 2414 19828 2466
rect 19840 2414 19892 2466
rect 5648 1870 5700 1922
rect 5712 1870 5764 1922
rect 5776 1870 5828 1922
rect 5840 1870 5892 1922
rect 14982 1870 15034 1922
rect 15046 1870 15098 1922
rect 15110 1870 15162 1922
rect 15174 1870 15226 1922
rect 24315 1870 24367 1922
rect 24379 1870 24431 1922
rect 24443 1870 24495 1922
rect 24507 1870 24559 1922
<< metal2 >>
rect 294 27240 350 27720
rect 938 27240 994 27720
rect 1582 27240 1638 27720
rect 2318 27240 2374 27720
rect 2962 27240 3018 27720
rect 3698 27240 3754 27720
rect 4342 27240 4398 27720
rect 4986 27240 5042 27720
rect 5722 27240 5778 27720
rect 6366 27240 6422 27720
rect 7102 27240 7158 27720
rect 7746 27240 7802 27720
rect 8390 27240 8446 27720
rect 9126 27240 9182 27720
rect 9770 27240 9826 27720
rect 10506 27240 10562 27720
rect 11150 27240 11206 27720
rect 11886 27240 11942 27720
rect 12530 27240 12586 27720
rect 13174 27240 13230 27720
rect 13910 27240 13966 27720
rect 14554 27240 14610 27720
rect 15290 27240 15346 27720
rect 15934 27240 15990 27720
rect 16578 27240 16634 27720
rect 17314 27240 17370 27720
rect 17958 27240 18014 27720
rect 18694 27240 18750 27720
rect 19338 27240 19394 27720
rect 20074 27240 20130 27720
rect 20718 27240 20774 27720
rect 21362 27240 21418 27720
rect 22098 27240 22154 27720
rect 22742 27240 22798 27720
rect 23202 27424 23258 27433
rect 23202 27359 23258 27368
rect 308 27190 336 27240
rect 296 27184 348 27190
rect 296 27126 348 27132
rect 480 27184 532 27190
rect 480 27126 532 27132
rect 492 21886 520 27126
rect 480 21880 532 21886
rect 480 21822 532 21828
rect 480 21744 532 21750
rect 480 21686 532 21692
rect 492 10977 520 21686
rect 952 17369 980 27240
rect 938 17360 994 17369
rect 938 17295 994 17304
rect 1596 16825 1624 27240
rect 2332 17913 2360 27240
rect 2976 18457 3004 27240
rect 3422 22800 3478 22809
rect 3422 22735 3478 22744
rect 3436 20769 3464 22735
rect 3422 20760 3478 20769
rect 3422 20695 3478 20704
rect 3712 19137 3740 27240
rect 4356 23353 4384 27240
rect 4342 23344 4398 23353
rect 4342 23279 4398 23288
rect 5000 22265 5028 27240
rect 5736 24962 5764 27240
rect 5736 24934 6040 24962
rect 5622 24772 5918 24792
rect 5678 24770 5702 24772
rect 5758 24770 5782 24772
rect 5838 24770 5862 24772
rect 5700 24718 5702 24770
rect 5764 24718 5776 24770
rect 5838 24718 5840 24770
rect 5678 24716 5702 24718
rect 5758 24716 5782 24718
rect 5838 24716 5862 24718
rect 5622 24696 5918 24716
rect 5622 23684 5918 23704
rect 5678 23682 5702 23684
rect 5758 23682 5782 23684
rect 5838 23682 5862 23684
rect 5700 23630 5702 23682
rect 5764 23630 5776 23682
rect 5838 23630 5840 23682
rect 5678 23628 5702 23630
rect 5758 23628 5782 23630
rect 5838 23628 5862 23630
rect 5622 23608 5918 23628
rect 5622 22596 5918 22616
rect 5678 22594 5702 22596
rect 5758 22594 5782 22596
rect 5838 22594 5862 22596
rect 5700 22542 5702 22594
rect 5764 22542 5776 22594
rect 5838 22542 5840 22594
rect 5678 22540 5702 22542
rect 5758 22540 5782 22542
rect 5838 22540 5862 22542
rect 5622 22520 5918 22540
rect 4986 22256 5042 22265
rect 4986 22191 5042 22200
rect 5622 21508 5918 21528
rect 5678 21506 5702 21508
rect 5758 21506 5782 21508
rect 5838 21506 5862 21508
rect 5700 21454 5702 21506
rect 5764 21454 5776 21506
rect 5838 21454 5840 21506
rect 5678 21452 5702 21454
rect 5758 21452 5782 21454
rect 5838 21452 5862 21454
rect 5622 21432 5918 21452
rect 6012 20769 6040 24934
rect 6380 21585 6408 27240
rect 6366 21576 6422 21585
rect 6366 21511 6422 21520
rect 7116 21449 7144 27240
rect 7760 22401 7788 27240
rect 7746 22392 7802 22401
rect 7746 22327 7802 22336
rect 7102 21440 7158 21449
rect 7102 21375 7158 21384
rect 5998 20760 6054 20769
rect 5998 20695 6054 20704
rect 5622 20420 5918 20440
rect 5678 20418 5702 20420
rect 5758 20418 5782 20420
rect 5838 20418 5862 20420
rect 5700 20366 5702 20418
rect 5764 20366 5776 20418
rect 5838 20366 5840 20418
rect 5678 20364 5702 20366
rect 5758 20364 5782 20366
rect 5838 20364 5862 20366
rect 5622 20344 5918 20364
rect 5622 19332 5918 19352
rect 5678 19330 5702 19332
rect 5758 19330 5782 19332
rect 5838 19330 5862 19332
rect 5700 19278 5702 19330
rect 5764 19278 5776 19330
rect 5838 19278 5840 19330
rect 5678 19276 5702 19278
rect 5758 19276 5782 19278
rect 5838 19276 5862 19278
rect 5622 19256 5918 19276
rect 3698 19128 3754 19137
rect 3698 19063 3754 19072
rect 8404 19001 8432 27240
rect 9140 21177 9168 27240
rect 9784 24033 9812 27240
rect 10520 25506 10548 27240
rect 10520 25478 10732 25506
rect 10289 25316 10585 25336
rect 10345 25314 10369 25316
rect 10425 25314 10449 25316
rect 10505 25314 10529 25316
rect 10367 25262 10369 25314
rect 10431 25262 10443 25314
rect 10505 25262 10507 25314
rect 10345 25260 10369 25262
rect 10425 25260 10449 25262
rect 10505 25260 10529 25262
rect 10289 25240 10585 25260
rect 10289 24228 10585 24248
rect 10345 24226 10369 24228
rect 10425 24226 10449 24228
rect 10505 24226 10529 24228
rect 10367 24174 10369 24226
rect 10431 24174 10443 24226
rect 10505 24174 10507 24226
rect 10345 24172 10369 24174
rect 10425 24172 10449 24174
rect 10505 24172 10529 24174
rect 10289 24152 10585 24172
rect 10704 24169 10732 25478
rect 11060 24464 11112 24470
rect 11060 24406 11112 24412
rect 11072 24316 11100 24406
rect 10888 24288 11100 24316
rect 10690 24160 10746 24169
rect 10690 24095 10746 24104
rect 9770 24024 9826 24033
rect 9770 23959 9826 23968
rect 10289 23140 10585 23160
rect 10345 23138 10369 23140
rect 10425 23138 10449 23140
rect 10505 23138 10529 23140
rect 10367 23086 10369 23138
rect 10431 23086 10443 23138
rect 10505 23086 10507 23138
rect 10345 23084 10369 23086
rect 10425 23084 10449 23086
rect 10505 23084 10529 23086
rect 10289 23064 10585 23084
rect 10888 22770 10916 24288
rect 11060 23784 11112 23790
rect 10980 23732 11060 23738
rect 10980 23726 11112 23732
rect 10980 23710 11100 23726
rect 10980 23042 11008 23710
rect 11164 23625 11192 27240
rect 11428 24872 11480 24878
rect 11428 24814 11480 24820
rect 11244 24532 11296 24538
rect 11244 24474 11296 24480
rect 11256 24334 11284 24474
rect 11440 24470 11468 24814
rect 11428 24464 11480 24470
rect 11428 24406 11480 24412
rect 11244 24328 11296 24334
rect 11244 24270 11296 24276
rect 11796 24328 11848 24334
rect 11796 24270 11848 24276
rect 11150 23616 11206 23625
rect 11150 23551 11206 23560
rect 10968 23036 11020 23042
rect 10968 22978 11020 22984
rect 11060 23036 11112 23042
rect 11060 22978 11112 22984
rect 10876 22764 10928 22770
rect 10876 22706 10928 22712
rect 11072 22498 11100 22978
rect 11152 22900 11204 22906
rect 11152 22842 11204 22848
rect 11060 22492 11112 22498
rect 11060 22434 11112 22440
rect 11164 22294 11192 22842
rect 11256 22809 11284 24270
rect 11808 23790 11836 24270
rect 11796 23784 11848 23790
rect 11796 23726 11848 23732
rect 11336 23376 11388 23382
rect 11336 23318 11388 23324
rect 11242 22800 11298 22809
rect 11242 22735 11298 22744
rect 11348 22362 11376 23318
rect 11900 23042 11928 27240
rect 12544 24441 12572 27240
rect 13188 24577 13216 27240
rect 13174 24568 13230 24577
rect 13174 24503 13230 24512
rect 12530 24432 12586 24441
rect 12348 24396 12400 24402
rect 12530 24367 12586 24376
rect 12348 24338 12400 24344
rect 12164 23308 12216 23314
rect 12164 23250 12216 23256
rect 12176 23081 12204 23250
rect 12256 23240 12308 23246
rect 12256 23182 12308 23188
rect 12162 23072 12218 23081
rect 11888 23036 11940 23042
rect 12162 23007 12218 23016
rect 11888 22978 11940 22984
rect 12268 22838 12296 23182
rect 12360 23058 12388 24338
rect 13176 23988 13228 23994
rect 13176 23930 13228 23936
rect 13188 23586 13216 23930
rect 13820 23920 13872 23926
rect 13820 23862 13872 23868
rect 13450 23616 13506 23625
rect 13176 23580 13228 23586
rect 13450 23551 13452 23560
rect 13176 23522 13228 23528
rect 13504 23551 13506 23560
rect 13452 23522 13504 23528
rect 13832 23382 13860 23862
rect 13820 23376 13872 23382
rect 13820 23318 13872 23324
rect 13820 23240 13872 23246
rect 13820 23182 13872 23188
rect 12360 23030 12480 23058
rect 12452 22906 12480 23030
rect 12440 22900 12492 22906
rect 12440 22842 12492 22848
rect 12992 22900 13044 22906
rect 12992 22842 13044 22848
rect 11612 22832 11664 22838
rect 11612 22774 11664 22780
rect 12256 22832 12308 22838
rect 12256 22774 12308 22780
rect 12714 22800 12770 22809
rect 11336 22356 11388 22362
rect 11336 22298 11388 22304
rect 11624 22294 11652 22774
rect 12714 22735 12770 22744
rect 12728 22498 12756 22735
rect 13004 22498 13032 22842
rect 13728 22832 13780 22838
rect 13726 22800 13728 22809
rect 13780 22800 13782 22809
rect 13726 22735 13782 22744
rect 13728 22696 13780 22702
rect 13728 22638 13780 22644
rect 12716 22492 12768 22498
rect 12716 22434 12768 22440
rect 12992 22492 13044 22498
rect 12992 22434 13044 22440
rect 11152 22288 11204 22294
rect 11152 22230 11204 22236
rect 11612 22288 11664 22294
rect 11612 22230 11664 22236
rect 10289 22052 10585 22072
rect 10345 22050 10369 22052
rect 10425 22050 10449 22052
rect 10505 22050 10529 22052
rect 10367 21998 10369 22050
rect 10431 21998 10443 22050
rect 10505 21998 10507 22050
rect 10345 21996 10369 21998
rect 10425 21996 10449 21998
rect 10505 21996 10529 21998
rect 10289 21976 10585 21996
rect 11624 21954 11652 22230
rect 11796 22220 11848 22226
rect 11796 22162 11848 22168
rect 11612 21948 11664 21954
rect 11612 21890 11664 21896
rect 11518 21576 11574 21585
rect 11518 21511 11574 21520
rect 11532 21410 11560 21511
rect 11520 21404 11572 21410
rect 11520 21346 11572 21352
rect 9126 21168 9182 21177
rect 9126 21103 9182 21112
rect 11808 21070 11836 22162
rect 13740 22129 13768 22638
rect 13726 22120 13782 22129
rect 13726 22055 13782 22064
rect 13832 21818 13860 23182
rect 13820 21812 13872 21818
rect 13820 21754 13872 21760
rect 12624 21608 12676 21614
rect 12624 21550 12676 21556
rect 12636 21274 12664 21550
rect 12624 21268 12676 21274
rect 12624 21210 12676 21216
rect 11704 21064 11756 21070
rect 11704 21006 11756 21012
rect 11796 21064 11848 21070
rect 12440 21064 12492 21070
rect 11796 21006 11848 21012
rect 12268 21012 12440 21018
rect 12268 21006 12492 21012
rect 10289 20964 10585 20984
rect 10345 20962 10369 20964
rect 10425 20962 10449 20964
rect 10505 20962 10529 20964
rect 10367 20910 10369 20962
rect 10431 20910 10443 20962
rect 10505 20910 10507 20962
rect 10345 20908 10369 20910
rect 10425 20908 10449 20910
rect 10505 20908 10529 20910
rect 10289 20888 10585 20908
rect 10874 20080 10930 20089
rect 10874 20015 10876 20024
rect 10928 20015 10930 20024
rect 10876 19986 10928 19992
rect 10289 19876 10585 19896
rect 10345 19874 10369 19876
rect 10425 19874 10449 19876
rect 10505 19874 10529 19876
rect 10367 19822 10369 19874
rect 10431 19822 10443 19874
rect 10505 19822 10507 19874
rect 10345 19820 10369 19822
rect 10425 19820 10449 19822
rect 10505 19820 10529 19822
rect 10289 19800 10585 19820
rect 10888 19778 10916 19986
rect 11716 19778 11744 21006
rect 11808 20526 11836 21006
rect 12268 20990 12480 21006
rect 11796 20520 11848 20526
rect 11796 20462 11848 20468
rect 10876 19772 10928 19778
rect 10876 19714 10928 19720
rect 11704 19772 11756 19778
rect 11704 19714 11756 19720
rect 11716 19098 11744 19714
rect 11704 19092 11756 19098
rect 11704 19034 11756 19040
rect 8390 18992 8446 19001
rect 8390 18927 8446 18936
rect 10289 18788 10585 18808
rect 10345 18786 10369 18788
rect 10425 18786 10449 18788
rect 10505 18786 10529 18788
rect 10367 18734 10369 18786
rect 10431 18734 10443 18786
rect 10505 18734 10507 18786
rect 10345 18732 10369 18734
rect 10425 18732 10449 18734
rect 10505 18732 10529 18734
rect 10289 18712 10585 18732
rect 2962 18448 3018 18457
rect 2962 18383 3018 18392
rect 5622 18244 5918 18264
rect 5678 18242 5702 18244
rect 5758 18242 5782 18244
rect 5838 18242 5862 18244
rect 5700 18190 5702 18242
rect 5764 18190 5776 18242
rect 5838 18190 5840 18242
rect 5678 18188 5702 18190
rect 5758 18188 5782 18190
rect 5838 18188 5862 18190
rect 5622 18168 5918 18188
rect 2318 17904 2374 17913
rect 2318 17839 2374 17848
rect 10289 17700 10585 17720
rect 10345 17698 10369 17700
rect 10425 17698 10449 17700
rect 10505 17698 10529 17700
rect 10367 17646 10369 17698
rect 10431 17646 10443 17698
rect 10505 17646 10507 17698
rect 10345 17644 10369 17646
rect 10425 17644 10449 17646
rect 10505 17644 10529 17646
rect 10289 17624 10585 17644
rect 5622 17156 5918 17176
rect 5678 17154 5702 17156
rect 5758 17154 5782 17156
rect 5838 17154 5862 17156
rect 5700 17102 5702 17154
rect 5764 17102 5776 17154
rect 5838 17102 5840 17154
rect 5678 17100 5702 17102
rect 5758 17100 5782 17102
rect 5838 17100 5862 17102
rect 5622 17080 5918 17100
rect 11808 16961 11836 20462
rect 12268 18894 12296 20990
rect 12636 20798 12664 21210
rect 13542 21168 13598 21177
rect 13542 21103 13544 21112
rect 13596 21103 13598 21112
rect 13544 21074 13596 21080
rect 13832 20866 13860 21754
rect 13820 20860 13872 20866
rect 13820 20802 13872 20808
rect 12624 20792 12676 20798
rect 12624 20734 12676 20740
rect 12440 20656 12492 20662
rect 12440 20598 12492 20604
rect 12452 20322 12480 20598
rect 12440 20316 12492 20322
rect 12440 20258 12492 20264
rect 12452 20118 12480 20258
rect 12440 20112 12492 20118
rect 12440 20054 12492 20060
rect 12636 20050 12664 20734
rect 13820 20520 13872 20526
rect 13542 20488 13598 20497
rect 13820 20462 13872 20468
rect 13542 20423 13598 20432
rect 12716 20112 12768 20118
rect 12716 20054 12768 20060
rect 12992 20112 13044 20118
rect 12992 20054 13044 20060
rect 12624 20044 12676 20050
rect 12624 19986 12676 19992
rect 12728 19642 12756 20054
rect 13004 19778 13032 20054
rect 13268 20044 13320 20050
rect 13268 19986 13320 19992
rect 13280 19778 13308 19986
rect 12992 19772 13044 19778
rect 12992 19714 13044 19720
rect 13268 19772 13320 19778
rect 13268 19714 13320 19720
rect 12716 19636 12768 19642
rect 12716 19578 12768 19584
rect 12440 19568 12492 19574
rect 12440 19510 12492 19516
rect 12348 19160 12400 19166
rect 12348 19102 12400 19108
rect 12256 18888 12308 18894
rect 12256 18830 12308 18836
rect 12360 18690 12388 19102
rect 12452 19030 12480 19510
rect 13004 19098 13032 19714
rect 12992 19092 13044 19098
rect 12992 19034 13044 19040
rect 12440 19024 12492 19030
rect 12440 18966 12492 18972
rect 13450 18992 13506 19001
rect 13450 18927 13452 18936
rect 13504 18927 13506 18936
rect 13452 18898 13504 18904
rect 12348 18684 12400 18690
rect 12348 18626 12400 18632
rect 11794 16952 11850 16961
rect 11794 16887 11850 16896
rect 1582 16816 1638 16825
rect 1582 16751 1638 16760
rect 10289 16612 10585 16632
rect 10345 16610 10369 16612
rect 10425 16610 10449 16612
rect 10505 16610 10529 16612
rect 10367 16558 10369 16610
rect 10431 16558 10443 16610
rect 10505 16558 10507 16610
rect 10345 16556 10369 16558
rect 10425 16556 10449 16558
rect 10505 16556 10529 16558
rect 10289 16536 10585 16556
rect 5622 16068 5918 16088
rect 5678 16066 5702 16068
rect 5758 16066 5782 16068
rect 5838 16066 5862 16068
rect 5700 16014 5702 16066
rect 5764 16014 5776 16066
rect 5838 16014 5840 16066
rect 5678 16012 5702 16014
rect 5758 16012 5782 16014
rect 5838 16012 5862 16014
rect 5622 15992 5918 16012
rect 10289 15524 10585 15544
rect 10345 15522 10369 15524
rect 10425 15522 10449 15524
rect 10505 15522 10529 15524
rect 10367 15470 10369 15522
rect 10431 15470 10443 15522
rect 10505 15470 10507 15522
rect 10345 15468 10369 15470
rect 10425 15468 10449 15470
rect 10505 15468 10529 15470
rect 10289 15448 10585 15468
rect 5622 14980 5918 15000
rect 5678 14978 5702 14980
rect 5758 14978 5782 14980
rect 5838 14978 5862 14980
rect 5700 14926 5702 14978
rect 5764 14926 5776 14978
rect 5838 14926 5840 14978
rect 5678 14924 5702 14926
rect 5758 14924 5782 14926
rect 5838 14924 5862 14926
rect 5622 14904 5918 14924
rect 10289 14436 10585 14456
rect 10345 14434 10369 14436
rect 10425 14434 10449 14436
rect 10505 14434 10529 14436
rect 10367 14382 10369 14434
rect 10431 14382 10443 14434
rect 10505 14382 10507 14434
rect 10345 14380 10369 14382
rect 10425 14380 10449 14382
rect 10505 14380 10529 14382
rect 10289 14360 10585 14380
rect 13556 14338 13584 20423
rect 13832 20202 13860 20462
rect 13740 20174 13860 20202
rect 13740 20118 13768 20174
rect 13728 20112 13780 20118
rect 13728 20054 13780 20060
rect 13636 18888 13688 18894
rect 13634 18856 13636 18865
rect 13728 18888 13780 18894
rect 13688 18856 13690 18865
rect 13728 18830 13780 18836
rect 13634 18791 13690 18800
rect 13740 18690 13768 18830
rect 13728 18684 13780 18690
rect 13728 18626 13780 18632
rect 13636 15624 13688 15630
rect 13636 15566 13688 15572
rect 13648 15222 13676 15566
rect 13924 15465 13952 27240
rect 14280 23784 14332 23790
rect 14280 23726 14332 23732
rect 14292 23450 14320 23726
rect 14280 23444 14332 23450
rect 14280 23386 14332 23392
rect 14004 23240 14056 23246
rect 14004 23182 14056 23188
rect 14016 22129 14044 23182
rect 14292 22974 14320 23386
rect 14280 22968 14332 22974
rect 14280 22910 14332 22916
rect 14096 22696 14148 22702
rect 14096 22638 14148 22644
rect 14108 22362 14136 22638
rect 14292 22498 14320 22910
rect 14280 22492 14332 22498
rect 14280 22434 14332 22440
rect 14096 22356 14148 22362
rect 14096 22298 14148 22304
rect 14002 22120 14058 22129
rect 14002 22055 14058 22064
rect 14372 21948 14424 21954
rect 14372 21890 14424 21896
rect 14278 21712 14334 21721
rect 14278 21647 14280 21656
rect 14332 21647 14334 21656
rect 14280 21618 14332 21624
rect 14384 21410 14412 21890
rect 14372 21404 14424 21410
rect 14372 21346 14424 21352
rect 14568 20497 14596 27240
rect 14956 24772 15252 24792
rect 15012 24770 15036 24772
rect 15092 24770 15116 24772
rect 15172 24770 15196 24772
rect 15034 24718 15036 24770
rect 15098 24718 15110 24770
rect 15172 24718 15174 24770
rect 15012 24716 15036 24718
rect 15092 24716 15116 24718
rect 15172 24716 15196 24718
rect 14956 24696 15252 24716
rect 15304 24538 15332 27240
rect 15292 24532 15344 24538
rect 15292 24474 15344 24480
rect 15948 23994 15976 27240
rect 16212 24532 16264 24538
rect 16212 24474 16264 24480
rect 16118 24024 16174 24033
rect 15108 23988 15160 23994
rect 15108 23930 15160 23936
rect 15476 23988 15528 23994
rect 15476 23930 15528 23936
rect 15936 23988 15988 23994
rect 16118 23959 16174 23968
rect 15936 23930 15988 23936
rect 15120 23897 15148 23930
rect 15106 23888 15162 23897
rect 15106 23823 15162 23832
rect 14956 23684 15252 23704
rect 15012 23682 15036 23684
rect 15092 23682 15116 23684
rect 15172 23682 15196 23684
rect 15034 23630 15036 23682
rect 15098 23630 15110 23682
rect 15172 23630 15174 23682
rect 15012 23628 15036 23630
rect 15092 23628 15116 23630
rect 15172 23628 15196 23630
rect 14956 23608 15252 23628
rect 15292 23240 15344 23246
rect 15292 23182 15344 23188
rect 14830 23072 14886 23081
rect 14830 23007 14886 23016
rect 15198 23072 15254 23081
rect 15198 23007 15200 23016
rect 14844 21750 14872 23007
rect 15252 23007 15254 23016
rect 15200 22978 15252 22984
rect 14956 22596 15252 22616
rect 15012 22594 15036 22596
rect 15092 22594 15116 22596
rect 15172 22594 15196 22596
rect 15034 22542 15036 22594
rect 15098 22542 15110 22594
rect 15172 22542 15174 22594
rect 15012 22540 15036 22542
rect 15092 22540 15116 22542
rect 15172 22540 15196 22542
rect 14956 22520 15252 22540
rect 15304 21970 15332 23182
rect 15384 22356 15436 22362
rect 15384 22298 15436 22304
rect 15120 21954 15332 21970
rect 15108 21948 15332 21954
rect 15160 21942 15332 21948
rect 15108 21890 15160 21896
rect 14832 21744 14884 21750
rect 14832 21686 14884 21692
rect 14844 21410 14872 21686
rect 14956 21508 15252 21528
rect 15012 21506 15036 21508
rect 15092 21506 15116 21508
rect 15172 21506 15196 21508
rect 15034 21454 15036 21506
rect 15098 21454 15110 21506
rect 15172 21454 15174 21506
rect 15012 21452 15036 21454
rect 15092 21452 15116 21454
rect 15172 21452 15196 21454
rect 14956 21432 15252 21452
rect 14832 21404 14884 21410
rect 14832 21346 14884 21352
rect 14646 20896 14702 20905
rect 14646 20831 14648 20840
rect 14700 20831 14702 20840
rect 14648 20802 14700 20808
rect 15292 20724 15344 20730
rect 15292 20666 15344 20672
rect 14554 20488 14610 20497
rect 14554 20423 14610 20432
rect 14956 20420 15252 20440
rect 15012 20418 15036 20420
rect 15092 20418 15116 20420
rect 15172 20418 15196 20420
rect 15034 20366 15036 20418
rect 15098 20366 15110 20418
rect 15172 20366 15174 20418
rect 15012 20364 15036 20366
rect 15092 20364 15116 20366
rect 15172 20364 15196 20366
rect 14956 20344 15252 20364
rect 15304 20322 15332 20666
rect 15396 20662 15424 22298
rect 15384 20656 15436 20662
rect 15384 20598 15436 20604
rect 15384 20520 15436 20526
rect 15384 20462 15436 20468
rect 15292 20316 15344 20322
rect 15292 20258 15344 20264
rect 15396 20118 15424 20462
rect 15384 20112 15436 20118
rect 15384 20054 15436 20060
rect 14096 19976 14148 19982
rect 14096 19918 14148 19924
rect 15016 19976 15068 19982
rect 15016 19918 15068 19924
rect 14108 19710 14136 19918
rect 14096 19704 14148 19710
rect 14096 19646 14148 19652
rect 14108 19098 14136 19646
rect 15028 19642 15056 19918
rect 15396 19778 15424 20054
rect 15384 19772 15436 19778
rect 15384 19714 15436 19720
rect 14740 19636 14792 19642
rect 14740 19578 14792 19584
rect 15016 19636 15068 19642
rect 15016 19578 15068 19584
rect 14752 19234 14780 19578
rect 14956 19332 15252 19352
rect 15012 19330 15036 19332
rect 15092 19330 15116 19332
rect 15172 19330 15196 19332
rect 15034 19278 15036 19330
rect 15098 19278 15110 19330
rect 15172 19278 15174 19330
rect 15012 19276 15036 19278
rect 15092 19276 15116 19278
rect 15172 19276 15196 19278
rect 14956 19256 15252 19276
rect 14740 19228 14792 19234
rect 14740 19170 14792 19176
rect 14096 19092 14148 19098
rect 14096 19034 14148 19040
rect 14108 18690 14136 19034
rect 14648 18888 14700 18894
rect 14648 18830 14700 18836
rect 14096 18684 14148 18690
rect 14096 18626 14148 18632
rect 14660 17602 14688 18830
rect 14648 17596 14700 17602
rect 14648 17538 14700 17544
rect 14188 17460 14240 17466
rect 14188 17402 14240 17408
rect 14004 17256 14056 17262
rect 14004 17198 14056 17204
rect 14016 15970 14044 17198
rect 14200 16854 14228 17402
rect 14188 16848 14240 16854
rect 14186 16816 14188 16825
rect 14240 16816 14242 16825
rect 14186 16751 14242 16760
rect 14660 16718 14688 17538
rect 14752 17534 14780 19170
rect 15396 19098 15424 19714
rect 15384 19092 15436 19098
rect 15384 19034 15436 19040
rect 15396 18690 15424 19034
rect 15384 18684 15436 18690
rect 15384 18626 15436 18632
rect 14956 18244 15252 18264
rect 15012 18242 15036 18244
rect 15092 18242 15116 18244
rect 15172 18242 15196 18244
rect 15034 18190 15036 18242
rect 15098 18190 15110 18242
rect 15172 18190 15174 18242
rect 15012 18188 15036 18190
rect 15092 18188 15116 18190
rect 15172 18188 15196 18190
rect 14956 18168 15252 18188
rect 15382 18176 15438 18185
rect 15382 18111 15384 18120
rect 15436 18111 15438 18120
rect 15384 18082 15436 18088
rect 15292 17800 15344 17806
rect 15292 17742 15344 17748
rect 14740 17528 14792 17534
rect 14792 17476 14872 17482
rect 14740 17470 14872 17476
rect 14752 17454 14872 17470
rect 14740 17392 14792 17398
rect 14740 17334 14792 17340
rect 14752 16786 14780 17334
rect 14844 17058 14872 17454
rect 14956 17156 15252 17176
rect 15012 17154 15036 17156
rect 15092 17154 15116 17156
rect 15172 17154 15196 17156
rect 15034 17102 15036 17154
rect 15098 17102 15110 17154
rect 15172 17102 15174 17154
rect 15012 17100 15036 17102
rect 15092 17100 15116 17102
rect 15172 17100 15196 17102
rect 14956 17080 15252 17100
rect 14832 17052 14884 17058
rect 14832 16994 14884 17000
rect 14740 16780 14792 16786
rect 14740 16722 14792 16728
rect 14648 16712 14700 16718
rect 14648 16654 14700 16660
rect 14280 16304 14332 16310
rect 14280 16246 14332 16252
rect 14004 15964 14056 15970
rect 14004 15906 14056 15912
rect 14292 15630 14320 16246
rect 14280 15624 14332 15630
rect 14280 15566 14332 15572
rect 13910 15456 13966 15465
rect 13910 15391 13966 15400
rect 13910 15320 13966 15329
rect 13910 15255 13912 15264
rect 13964 15255 13966 15264
rect 13912 15226 13964 15232
rect 13636 15216 13688 15222
rect 13636 15158 13688 15164
rect 13648 14542 13676 15158
rect 13924 14882 13952 15226
rect 14660 14882 14688 16654
rect 14752 16446 14780 16722
rect 14740 16440 14792 16446
rect 14740 16382 14792 16388
rect 14752 15630 14780 16382
rect 14956 16068 15252 16088
rect 15012 16066 15036 16068
rect 15092 16066 15116 16068
rect 15172 16066 15196 16068
rect 15034 16014 15036 16066
rect 15098 16014 15110 16066
rect 15172 16014 15174 16066
rect 15012 16012 15036 16014
rect 15092 16012 15116 16014
rect 15172 16012 15196 16014
rect 14956 15992 15252 16012
rect 15304 15970 15332 17742
rect 15384 17256 15436 17262
rect 15384 17198 15436 17204
rect 15396 16854 15424 17198
rect 15384 16848 15436 16854
rect 15384 16790 15436 16796
rect 15396 16514 15424 16790
rect 15384 16508 15436 16514
rect 15384 16450 15436 16456
rect 15292 15964 15344 15970
rect 15292 15906 15344 15912
rect 14740 15624 14792 15630
rect 14740 15566 14792 15572
rect 14752 15426 14780 15566
rect 14740 15420 14792 15426
rect 14740 15362 14792 15368
rect 15292 15284 15344 15290
rect 15292 15226 15344 15232
rect 14956 14980 15252 15000
rect 15012 14978 15036 14980
rect 15092 14978 15116 14980
rect 15172 14978 15196 14980
rect 15034 14926 15036 14978
rect 15098 14926 15110 14978
rect 15172 14926 15174 14978
rect 15012 14924 15036 14926
rect 15092 14924 15116 14926
rect 15172 14924 15196 14926
rect 14956 14904 15252 14924
rect 15304 14882 15332 15226
rect 15488 14882 15516 23930
rect 16132 23926 16160 23959
rect 16120 23920 16172 23926
rect 16120 23862 16172 23868
rect 16132 23586 16160 23862
rect 16120 23580 16172 23586
rect 16120 23522 16172 23528
rect 15936 23308 15988 23314
rect 15936 23250 15988 23256
rect 15948 22362 15976 23250
rect 16028 22696 16080 22702
rect 16028 22638 16080 22644
rect 15936 22356 15988 22362
rect 15936 22298 15988 22304
rect 16040 22294 16068 22638
rect 16028 22288 16080 22294
rect 16028 22230 16080 22236
rect 15568 22220 15620 22226
rect 15568 22162 15620 22168
rect 15580 21410 15608 22162
rect 16028 21744 16080 21750
rect 16028 21686 16080 21692
rect 15752 21608 15804 21614
rect 15752 21550 15804 21556
rect 15568 21404 15620 21410
rect 15568 21346 15620 21352
rect 15764 20730 15792 21550
rect 16040 21410 16068 21686
rect 16028 21404 16080 21410
rect 16028 21346 16080 21352
rect 15844 21064 15896 21070
rect 15842 21032 15844 21041
rect 15896 21032 15898 21041
rect 15842 20967 15898 20976
rect 15752 20724 15804 20730
rect 15752 20666 15804 20672
rect 15660 20656 15712 20662
rect 15566 20624 15622 20633
rect 15660 20598 15712 20604
rect 15566 20559 15622 20568
rect 15580 18894 15608 20559
rect 15672 19982 15700 20598
rect 15660 19976 15712 19982
rect 15660 19918 15712 19924
rect 15672 19710 15700 19918
rect 15660 19704 15712 19710
rect 15660 19646 15712 19652
rect 15660 19568 15712 19574
rect 15660 19510 15712 19516
rect 15672 19030 15700 19510
rect 15660 19024 15712 19030
rect 15660 18966 15712 18972
rect 15568 18888 15620 18894
rect 15752 18888 15804 18894
rect 15568 18830 15620 18836
rect 15750 18856 15752 18865
rect 15804 18856 15806 18865
rect 15750 18791 15806 18800
rect 15764 18690 15792 18791
rect 15752 18684 15804 18690
rect 15752 18626 15804 18632
rect 16120 18344 16172 18350
rect 16120 18286 16172 18292
rect 15936 18004 15988 18010
rect 15936 17946 15988 17952
rect 15948 17534 15976 17946
rect 16132 17874 16160 18286
rect 16120 17868 16172 17874
rect 16120 17810 16172 17816
rect 15936 17528 15988 17534
rect 15936 17470 15988 17476
rect 15752 17460 15804 17466
rect 15752 17402 15804 17408
rect 15764 16378 15792 17402
rect 15948 17058 15976 17470
rect 15936 17052 15988 17058
rect 15936 16994 15988 17000
rect 15844 16508 15896 16514
rect 15844 16450 15896 16456
rect 15752 16372 15804 16378
rect 15752 16314 15804 16320
rect 15660 15624 15712 15630
rect 15658 15592 15660 15601
rect 15712 15592 15714 15601
rect 15658 15527 15714 15536
rect 13912 14876 13964 14882
rect 13912 14818 13964 14824
rect 14648 14876 14700 14882
rect 14648 14818 14700 14824
rect 15292 14876 15344 14882
rect 15292 14818 15344 14824
rect 15476 14876 15528 14882
rect 15476 14818 15528 14824
rect 15764 14814 15792 16314
rect 15856 15834 15884 16450
rect 16132 15902 16160 17810
rect 16120 15896 16172 15902
rect 16120 15838 16172 15844
rect 15844 15828 15896 15834
rect 15844 15770 15896 15776
rect 15856 15426 15884 15770
rect 15844 15420 15896 15426
rect 15844 15362 15896 15368
rect 15936 15080 15988 15086
rect 15936 15022 15988 15028
rect 15752 14808 15804 14814
rect 15948 14785 15976 15022
rect 15752 14750 15804 14756
rect 15934 14776 15990 14785
rect 15384 14672 15436 14678
rect 15384 14614 15436 14620
rect 13636 14536 13688 14542
rect 13636 14478 13688 14484
rect 13544 14332 13596 14338
rect 13544 14274 13596 14280
rect 13452 14196 13504 14202
rect 13452 14138 13504 14144
rect 5622 13892 5918 13912
rect 5678 13890 5702 13892
rect 5758 13890 5782 13892
rect 5838 13890 5862 13892
rect 5700 13838 5702 13890
rect 5764 13838 5776 13890
rect 5838 13838 5840 13890
rect 5678 13836 5702 13838
rect 5758 13836 5782 13838
rect 5838 13836 5862 13838
rect 5622 13816 5918 13836
rect 13464 13794 13492 14138
rect 13452 13788 13504 13794
rect 13452 13730 13504 13736
rect 13176 13448 13228 13454
rect 13176 13390 13228 13396
rect 10289 13348 10585 13368
rect 10345 13346 10369 13348
rect 10425 13346 10449 13348
rect 10505 13346 10529 13348
rect 10367 13294 10369 13346
rect 10431 13294 10443 13346
rect 10505 13294 10507 13346
rect 10345 13292 10369 13294
rect 10425 13292 10449 13294
rect 10505 13292 10529 13294
rect 10289 13272 10585 13292
rect 12992 13040 13044 13046
rect 12992 12982 13044 12988
rect 5622 12804 5918 12824
rect 5678 12802 5702 12804
rect 5758 12802 5782 12804
rect 5838 12802 5862 12804
rect 5700 12750 5702 12802
rect 5764 12750 5776 12802
rect 5838 12750 5840 12802
rect 5678 12748 5702 12750
rect 5758 12748 5782 12750
rect 5838 12748 5862 12750
rect 5622 12728 5918 12748
rect 13004 12706 13032 12982
rect 13188 12706 13216 13390
rect 13268 12904 13320 12910
rect 13268 12846 13320 12852
rect 12992 12700 13044 12706
rect 12992 12642 13044 12648
rect 13176 12700 13228 12706
rect 13176 12642 13228 12648
rect 13280 12570 13308 12846
rect 13268 12564 13320 12570
rect 13268 12506 13320 12512
rect 13084 12428 13136 12434
rect 13084 12370 13136 12376
rect 10289 12260 10585 12280
rect 10345 12258 10369 12260
rect 10425 12258 10449 12260
rect 10505 12258 10529 12260
rect 10367 12206 10369 12258
rect 10431 12206 10443 12258
rect 10505 12206 10507 12258
rect 10345 12204 10369 12206
rect 10425 12204 10449 12206
rect 10505 12204 10529 12206
rect 10289 12184 10585 12204
rect 12532 12020 12584 12026
rect 12532 11962 12584 11968
rect 5622 11716 5918 11736
rect 5678 11714 5702 11716
rect 5758 11714 5782 11716
rect 5838 11714 5862 11716
rect 5700 11662 5702 11714
rect 5764 11662 5776 11714
rect 5838 11662 5840 11714
rect 5678 11660 5702 11662
rect 5758 11660 5782 11662
rect 5838 11660 5862 11662
rect 5622 11640 5918 11660
rect 12544 11482 12572 11962
rect 12532 11476 12584 11482
rect 12532 11418 12584 11424
rect 10048 11408 10100 11414
rect 3422 11376 3478 11385
rect 10048 11350 10100 11356
rect 10138 11376 10194 11385
rect 3422 11311 3478 11320
rect 478 10968 534 10977
rect 478 10903 534 10912
rect 3436 6761 3464 11311
rect 10060 11074 10088 11350
rect 10138 11311 10140 11320
rect 10192 11311 10194 11320
rect 12808 11340 12860 11346
rect 10140 11282 10192 11288
rect 12808 11282 12860 11288
rect 10289 11172 10585 11192
rect 10345 11170 10369 11172
rect 10425 11170 10449 11172
rect 10505 11170 10529 11172
rect 10367 11118 10369 11170
rect 10431 11118 10443 11170
rect 10505 11118 10507 11170
rect 10345 11116 10369 11118
rect 10425 11116 10449 11118
rect 10505 11116 10529 11118
rect 10289 11096 10585 11116
rect 10048 11068 10100 11074
rect 10048 11010 10100 11016
rect 12820 10802 12848 11282
rect 13096 11074 13124 12370
rect 13280 12094 13308 12506
rect 13648 12094 13676 14478
rect 15396 13998 15424 14614
rect 15764 14270 15792 14750
rect 15934 14711 15990 14720
rect 15752 14264 15804 14270
rect 15752 14206 15804 14212
rect 15384 13992 15436 13998
rect 15384 13934 15436 13940
rect 14956 13892 15252 13912
rect 15012 13890 15036 13892
rect 15092 13890 15116 13892
rect 15172 13890 15196 13892
rect 15034 13838 15036 13890
rect 15098 13838 15110 13890
rect 15172 13838 15174 13890
rect 15012 13836 15036 13838
rect 15092 13836 15116 13838
rect 15172 13836 15196 13838
rect 14956 13816 15252 13836
rect 15396 13658 15424 13934
rect 15764 13794 15792 14206
rect 15752 13788 15804 13794
rect 15752 13730 15804 13736
rect 15936 13788 15988 13794
rect 15936 13730 15988 13736
rect 15384 13652 15436 13658
rect 15384 13594 15436 13600
rect 15292 13584 15344 13590
rect 15292 13526 15344 13532
rect 14956 12804 15252 12824
rect 15012 12802 15036 12804
rect 15092 12802 15116 12804
rect 15172 12802 15196 12804
rect 15034 12750 15036 12802
rect 15098 12750 15110 12802
rect 15172 12750 15174 12802
rect 15012 12748 15036 12750
rect 15092 12748 15116 12750
rect 15172 12748 15196 12750
rect 14956 12728 15252 12748
rect 15304 12706 15332 13526
rect 15844 12904 15896 12910
rect 15844 12846 15896 12852
rect 15292 12700 15344 12706
rect 15292 12642 15344 12648
rect 15856 12570 15884 12846
rect 15844 12564 15896 12570
rect 15844 12506 15896 12512
rect 15384 12428 15436 12434
rect 15384 12370 15436 12376
rect 13268 12088 13320 12094
rect 13268 12030 13320 12036
rect 13636 12088 13688 12094
rect 13636 12030 13688 12036
rect 13280 11618 13308 12030
rect 15292 12020 15344 12026
rect 15292 11962 15344 11968
rect 14372 11816 14424 11822
rect 14372 11758 14424 11764
rect 14384 11618 14412 11758
rect 14956 11716 15252 11736
rect 15012 11714 15036 11716
rect 15092 11714 15116 11716
rect 15172 11714 15196 11716
rect 15034 11662 15036 11714
rect 15098 11662 15110 11714
rect 15172 11662 15174 11714
rect 15012 11660 15036 11662
rect 15092 11660 15116 11662
rect 15172 11660 15196 11662
rect 14956 11640 15252 11660
rect 15304 11618 15332 11962
rect 13268 11612 13320 11618
rect 13268 11554 13320 11560
rect 14372 11612 14424 11618
rect 14372 11554 14424 11560
rect 15292 11612 15344 11618
rect 15292 11554 15344 11560
rect 13084 11068 13136 11074
rect 13084 11010 13136 11016
rect 13542 10968 13598 10977
rect 13176 10932 13228 10938
rect 13542 10903 13598 10912
rect 13176 10874 13228 10880
rect 12808 10796 12860 10802
rect 12808 10738 12860 10744
rect 5622 10628 5918 10648
rect 5678 10626 5702 10628
rect 5758 10626 5782 10628
rect 5838 10626 5862 10628
rect 5700 10574 5702 10626
rect 5764 10574 5776 10626
rect 5838 10574 5840 10626
rect 5678 10572 5702 10574
rect 5758 10572 5782 10574
rect 5838 10572 5862 10574
rect 5622 10552 5918 10572
rect 13188 10190 13216 10874
rect 13556 10870 13584 10903
rect 13544 10864 13596 10870
rect 13544 10806 13596 10812
rect 13728 10864 13780 10870
rect 13780 10812 13860 10818
rect 13728 10806 13860 10812
rect 13556 10462 13584 10806
rect 13740 10790 13860 10806
rect 15304 10802 15332 11554
rect 15396 11482 15424 12370
rect 15568 12360 15620 12366
rect 15568 12302 15620 12308
rect 15384 11476 15436 11482
rect 15384 11418 15436 11424
rect 15580 11074 15608 12302
rect 15948 12094 15976 13730
rect 15936 12088 15988 12094
rect 15936 12030 15988 12036
rect 15948 11618 15976 12030
rect 15936 11612 15988 11618
rect 15936 11554 15988 11560
rect 15568 11068 15620 11074
rect 15568 11010 15620 11016
rect 16028 11000 16080 11006
rect 16028 10942 16080 10948
rect 15660 10932 15712 10938
rect 15660 10874 15712 10880
rect 13832 10530 13860 10790
rect 15292 10796 15344 10802
rect 15292 10738 15344 10744
rect 14956 10628 15252 10648
rect 15012 10626 15036 10628
rect 15092 10626 15116 10628
rect 15172 10626 15196 10628
rect 15034 10574 15036 10626
rect 15098 10574 15110 10626
rect 15172 10574 15174 10626
rect 15012 10572 15036 10574
rect 15092 10572 15116 10574
rect 15172 10572 15196 10574
rect 14956 10552 15252 10572
rect 13820 10524 13872 10530
rect 13820 10466 13872 10472
rect 13544 10456 13596 10462
rect 13544 10398 13596 10404
rect 15672 10190 15700 10874
rect 16040 10530 16068 10942
rect 16028 10524 16080 10530
rect 16028 10466 16080 10472
rect 13176 10184 13228 10190
rect 13176 10126 13228 10132
rect 15660 10184 15712 10190
rect 15660 10126 15712 10132
rect 10289 10084 10585 10104
rect 10345 10082 10369 10084
rect 10425 10082 10449 10084
rect 10505 10082 10529 10084
rect 10367 10030 10369 10082
rect 10431 10030 10443 10082
rect 10505 10030 10507 10082
rect 10345 10028 10369 10030
rect 10425 10028 10449 10030
rect 10505 10028 10529 10030
rect 10289 10008 10585 10028
rect 5622 9540 5918 9560
rect 5678 9538 5702 9540
rect 5758 9538 5782 9540
rect 5838 9538 5862 9540
rect 5700 9486 5702 9538
rect 5764 9486 5776 9538
rect 5838 9486 5840 9538
rect 5678 9484 5702 9486
rect 5758 9484 5782 9486
rect 5838 9484 5862 9486
rect 5622 9464 5918 9484
rect 10289 8996 10585 9016
rect 10345 8994 10369 8996
rect 10425 8994 10449 8996
rect 10505 8994 10529 8996
rect 10367 8942 10369 8994
rect 10431 8942 10443 8994
rect 10505 8942 10507 8994
rect 10345 8940 10369 8942
rect 10425 8940 10449 8942
rect 10505 8940 10529 8942
rect 10289 8920 10585 8940
rect 5622 8452 5918 8472
rect 5678 8450 5702 8452
rect 5758 8450 5782 8452
rect 5838 8450 5862 8452
rect 5700 8398 5702 8450
rect 5764 8398 5776 8450
rect 5838 8398 5840 8450
rect 5678 8396 5702 8398
rect 5758 8396 5782 8398
rect 5838 8396 5862 8398
rect 5622 8376 5918 8396
rect 10289 7908 10585 7928
rect 10345 7906 10369 7908
rect 10425 7906 10449 7908
rect 10505 7906 10529 7908
rect 10367 7854 10369 7906
rect 10431 7854 10443 7906
rect 10505 7854 10507 7906
rect 10345 7852 10369 7854
rect 10425 7852 10449 7854
rect 10505 7852 10529 7854
rect 10289 7832 10585 7852
rect 5622 7364 5918 7384
rect 5678 7362 5702 7364
rect 5758 7362 5782 7364
rect 5838 7362 5862 7364
rect 5700 7310 5702 7362
rect 5764 7310 5776 7362
rect 5838 7310 5840 7362
rect 5678 7308 5702 7310
rect 5758 7308 5782 7310
rect 5838 7308 5862 7310
rect 5622 7288 5918 7308
rect 10289 6820 10585 6840
rect 10345 6818 10369 6820
rect 10425 6818 10449 6820
rect 10505 6818 10529 6820
rect 10367 6766 10369 6818
rect 10431 6766 10443 6818
rect 10505 6766 10507 6818
rect 10345 6764 10369 6766
rect 10425 6764 10449 6766
rect 10505 6764 10529 6766
rect 3422 6752 3478 6761
rect 10289 6744 10585 6764
rect 3422 6687 3478 6696
rect 5622 6276 5918 6296
rect 5678 6274 5702 6276
rect 5758 6274 5782 6276
rect 5838 6274 5862 6276
rect 5700 6222 5702 6274
rect 5764 6222 5776 6274
rect 5838 6222 5840 6274
rect 5678 6220 5702 6222
rect 5758 6220 5782 6222
rect 5838 6220 5862 6222
rect 5622 6200 5918 6220
rect 13188 6081 13216 10126
rect 14956 9540 15252 9560
rect 15012 9538 15036 9540
rect 15092 9538 15116 9540
rect 15172 9538 15196 9540
rect 15034 9486 15036 9538
rect 15098 9486 15110 9538
rect 15172 9486 15174 9538
rect 15012 9484 15036 9486
rect 15092 9484 15116 9486
rect 15172 9484 15196 9486
rect 14956 9464 15252 9484
rect 14956 8452 15252 8472
rect 15012 8450 15036 8452
rect 15092 8450 15116 8452
rect 15172 8450 15196 8452
rect 15034 8398 15036 8450
rect 15098 8398 15110 8450
rect 15172 8398 15174 8450
rect 15012 8396 15036 8398
rect 15092 8396 15116 8398
rect 15172 8396 15196 8398
rect 14956 8376 15252 8396
rect 15672 7713 15700 10126
rect 15658 7704 15714 7713
rect 15658 7639 15714 7648
rect 14956 7364 15252 7384
rect 15012 7362 15036 7364
rect 15092 7362 15116 7364
rect 15172 7362 15196 7364
rect 15034 7310 15036 7362
rect 15098 7310 15110 7362
rect 15172 7310 15174 7362
rect 15012 7308 15036 7310
rect 15092 7308 15116 7310
rect 15172 7308 15196 7310
rect 14956 7288 15252 7308
rect 14956 6276 15252 6296
rect 15012 6274 15036 6276
rect 15092 6274 15116 6276
rect 15172 6274 15196 6276
rect 15034 6222 15036 6274
rect 15098 6222 15110 6274
rect 15172 6222 15174 6274
rect 15012 6220 15036 6222
rect 15092 6220 15116 6222
rect 15172 6220 15196 6222
rect 14956 6200 15252 6220
rect 13174 6072 13230 6081
rect 13174 6007 13230 6016
rect 10289 5732 10585 5752
rect 10345 5730 10369 5732
rect 10425 5730 10449 5732
rect 10505 5730 10529 5732
rect 10367 5678 10369 5730
rect 10431 5678 10443 5730
rect 10505 5678 10507 5730
rect 10345 5676 10369 5678
rect 10425 5676 10449 5678
rect 10505 5676 10529 5678
rect 10289 5656 10585 5676
rect 5622 5188 5918 5208
rect 5678 5186 5702 5188
rect 5758 5186 5782 5188
rect 5838 5186 5862 5188
rect 5700 5134 5702 5186
rect 5764 5134 5776 5186
rect 5838 5134 5840 5186
rect 5678 5132 5702 5134
rect 5758 5132 5782 5134
rect 5838 5132 5862 5134
rect 5622 5112 5918 5132
rect 14956 5188 15252 5208
rect 15012 5186 15036 5188
rect 15092 5186 15116 5188
rect 15172 5186 15196 5188
rect 15034 5134 15036 5186
rect 15098 5134 15110 5186
rect 15172 5134 15174 5186
rect 15012 5132 15036 5134
rect 15092 5132 15116 5134
rect 15172 5132 15196 5134
rect 14956 5112 15252 5132
rect 16224 5090 16252 24474
rect 16304 23784 16356 23790
rect 16304 23726 16356 23732
rect 16316 22974 16344 23726
rect 16304 22968 16356 22974
rect 16304 22910 16356 22916
rect 16394 22800 16450 22809
rect 16394 22735 16396 22744
rect 16448 22735 16450 22744
rect 16396 22706 16448 22712
rect 16488 22288 16540 22294
rect 16488 22230 16540 22236
rect 16500 21614 16528 22230
rect 16396 21608 16448 21614
rect 16396 21550 16448 21556
rect 16488 21608 16540 21614
rect 16488 21550 16540 21556
rect 16408 21070 16436 21550
rect 16488 21268 16540 21274
rect 16488 21210 16540 21216
rect 16396 21064 16448 21070
rect 16396 21006 16448 21012
rect 16408 19273 16436 21006
rect 16500 20730 16528 21210
rect 16488 20724 16540 20730
rect 16488 20666 16540 20672
rect 16500 20322 16528 20666
rect 16488 20316 16540 20322
rect 16488 20258 16540 20264
rect 16394 19264 16450 19273
rect 16394 19199 16450 19208
rect 16396 18480 16448 18486
rect 16396 18422 16448 18428
rect 16408 17942 16436 18422
rect 16488 18344 16540 18350
rect 16488 18286 16540 18292
rect 16396 17936 16448 17942
rect 16394 17904 16396 17913
rect 16448 17904 16450 17913
rect 16394 17839 16450 17848
rect 16500 17641 16528 18286
rect 16486 17632 16542 17641
rect 16486 17567 16542 17576
rect 16304 17052 16356 17058
rect 16304 16994 16356 17000
rect 16316 16514 16344 16994
rect 16304 16508 16356 16514
rect 16304 16450 16356 16456
rect 16488 16304 16540 16310
rect 16488 16246 16540 16252
rect 16500 15970 16528 16246
rect 16488 15964 16540 15970
rect 16488 15906 16540 15912
rect 16500 15766 16528 15906
rect 16488 15760 16540 15766
rect 16488 15702 16540 15708
rect 16394 15456 16450 15465
rect 16394 15391 16396 15400
rect 16448 15391 16450 15400
rect 16396 15362 16448 15368
rect 16304 15284 16356 15290
rect 16304 15226 16356 15232
rect 16316 15057 16344 15226
rect 16302 15048 16358 15057
rect 16302 14983 16358 14992
rect 16408 14882 16436 15362
rect 16396 14876 16448 14882
rect 16396 14818 16448 14824
rect 16396 14196 16448 14202
rect 16396 14138 16448 14144
rect 16408 13833 16436 14138
rect 16394 13824 16450 13833
rect 16394 13759 16396 13768
rect 16448 13759 16450 13768
rect 16396 13730 16448 13736
rect 16408 13699 16436 13730
rect 16488 12564 16540 12570
rect 16488 12506 16540 12512
rect 16500 12162 16528 12506
rect 16488 12156 16540 12162
rect 16488 12098 16540 12104
rect 16304 10796 16356 10802
rect 16304 10738 16356 10744
rect 16316 10530 16344 10738
rect 16304 10524 16356 10530
rect 16304 10466 16356 10472
rect 16592 6194 16620 27240
rect 17328 24554 17356 27240
rect 16960 24526 17356 24554
rect 16856 24328 16908 24334
rect 16856 24270 16908 24276
rect 16868 23926 16896 24270
rect 16856 23920 16908 23926
rect 16856 23862 16908 23868
rect 16868 23314 16896 23862
rect 16856 23308 16908 23314
rect 16856 23250 16908 23256
rect 16856 21744 16908 21750
rect 16856 21686 16908 21692
rect 16868 21614 16896 21686
rect 16856 21608 16908 21614
rect 16856 21550 16908 21556
rect 16868 20866 16896 21550
rect 16856 20860 16908 20866
rect 16856 20802 16908 20808
rect 16854 19264 16910 19273
rect 16854 19199 16910 19208
rect 16868 18622 16896 19199
rect 16856 18616 16908 18622
rect 16856 18558 16908 18564
rect 16868 18146 16896 18558
rect 16856 18140 16908 18146
rect 16856 18082 16908 18088
rect 16856 15148 16908 15154
rect 16856 15090 16908 15096
rect 16868 14610 16896 15090
rect 16856 14604 16908 14610
rect 16856 14546 16908 14552
rect 16868 14338 16896 14546
rect 16856 14332 16908 14338
rect 16856 14274 16908 14280
rect 16960 13794 16988 24526
rect 17408 24328 17460 24334
rect 17408 24270 17460 24276
rect 17316 23308 17368 23314
rect 17316 23250 17368 23256
rect 17224 23240 17276 23246
rect 17224 23182 17276 23188
rect 17236 22838 17264 23182
rect 17224 22832 17276 22838
rect 17224 22774 17276 22780
rect 17236 21954 17264 22774
rect 17328 22498 17356 23250
rect 17420 23042 17448 24270
rect 17408 23036 17460 23042
rect 17408 22978 17460 22984
rect 17420 22498 17448 22978
rect 17316 22492 17368 22498
rect 17316 22434 17368 22440
rect 17408 22492 17460 22498
rect 17408 22434 17460 22440
rect 17224 21948 17276 21954
rect 17224 21890 17276 21896
rect 17040 21812 17092 21818
rect 17040 21754 17092 21760
rect 17052 21070 17080 21754
rect 17592 21268 17644 21274
rect 17592 21210 17644 21216
rect 17604 21070 17632 21210
rect 17972 21154 18000 27240
rect 18708 24538 18736 27240
rect 18696 24532 18748 24538
rect 18696 24474 18748 24480
rect 19156 24532 19208 24538
rect 19156 24474 19208 24480
rect 18418 24160 18474 24169
rect 18418 24095 18474 24104
rect 18144 23988 18196 23994
rect 18144 23930 18196 23936
rect 18156 23625 18184 23930
rect 18432 23926 18460 24095
rect 18420 23920 18472 23926
rect 18420 23862 18472 23868
rect 18328 23784 18380 23790
rect 18328 23726 18380 23732
rect 18142 23616 18198 23625
rect 18142 23551 18144 23560
rect 18196 23551 18198 23560
rect 18144 23522 18196 23528
rect 18144 23376 18196 23382
rect 18144 23318 18196 23324
rect 18052 22832 18104 22838
rect 18156 22820 18184 23318
rect 18340 23314 18368 23726
rect 18432 23586 18460 23862
rect 18696 23784 18748 23790
rect 18696 23726 18748 23732
rect 18420 23580 18472 23586
rect 18420 23522 18472 23528
rect 18708 23382 18736 23726
rect 18786 23616 18842 23625
rect 18786 23551 18842 23560
rect 18696 23376 18748 23382
rect 18696 23318 18748 23324
rect 18328 23308 18380 23314
rect 18328 23250 18380 23256
rect 18328 22900 18380 22906
rect 18328 22842 18380 22848
rect 18104 22792 18184 22820
rect 18052 22774 18104 22780
rect 18156 22537 18184 22792
rect 18142 22528 18198 22537
rect 18340 22498 18368 22842
rect 18142 22463 18144 22472
rect 18196 22463 18198 22472
rect 18328 22492 18380 22498
rect 18144 22434 18196 22440
rect 18328 22434 18380 22440
rect 18418 22120 18474 22129
rect 18418 22055 18474 22064
rect 18326 21848 18382 21857
rect 18326 21783 18328 21792
rect 18380 21783 18382 21792
rect 18328 21754 18380 21760
rect 18326 21712 18382 21721
rect 18326 21647 18382 21656
rect 18340 21313 18368 21647
rect 18326 21304 18382 21313
rect 18326 21239 18382 21248
rect 17972 21126 18276 21154
rect 17040 21064 17092 21070
rect 17040 21006 17092 21012
rect 17592 21064 17644 21070
rect 17592 21006 17644 21012
rect 18052 21064 18104 21070
rect 18052 21006 18104 21012
rect 18144 21064 18196 21070
rect 18144 21006 18196 21012
rect 17052 20905 17080 21006
rect 17038 20896 17094 20905
rect 17038 20831 17094 20840
rect 17604 20089 17632 21006
rect 17958 20760 18014 20769
rect 17958 20695 18014 20704
rect 17972 20662 18000 20695
rect 17960 20656 18012 20662
rect 17960 20598 18012 20604
rect 17972 20322 18000 20598
rect 17960 20316 18012 20322
rect 17960 20258 18012 20264
rect 17590 20080 17646 20089
rect 17590 20015 17646 20024
rect 17960 19772 18012 19778
rect 17960 19714 18012 19720
rect 17592 18548 17644 18554
rect 17592 18490 17644 18496
rect 17604 18146 17632 18490
rect 17132 18140 17184 18146
rect 17132 18082 17184 18088
rect 17592 18140 17644 18146
rect 17592 18082 17644 18088
rect 17144 17602 17172 18082
rect 17132 17596 17184 17602
rect 17132 17538 17184 17544
rect 17868 15760 17920 15766
rect 17972 15748 18000 19714
rect 18064 19030 18092 21006
rect 18156 19642 18184 21006
rect 18144 19636 18196 19642
rect 18144 19578 18196 19584
rect 18052 19024 18104 19030
rect 18052 18966 18104 18972
rect 18052 18480 18104 18486
rect 18052 18422 18104 18428
rect 18064 17890 18092 18422
rect 18064 17862 18184 17890
rect 18156 17806 18184 17862
rect 18144 17800 18196 17806
rect 18144 17742 18196 17748
rect 18052 17460 18104 17466
rect 18052 17402 18104 17408
rect 18064 16990 18092 17402
rect 18052 16984 18104 16990
rect 18052 16926 18104 16932
rect 17920 15720 18000 15748
rect 17868 15702 17920 15708
rect 16948 13788 17000 13794
rect 16948 13730 17000 13736
rect 17972 13726 18000 15720
rect 18156 14610 18184 17742
rect 18144 14604 18196 14610
rect 18144 14546 18196 14552
rect 18052 14536 18104 14542
rect 18052 14478 18104 14484
rect 18064 14202 18092 14478
rect 18052 14196 18104 14202
rect 18052 14138 18104 14144
rect 18064 13794 18092 14138
rect 18156 14134 18184 14546
rect 18144 14128 18196 14134
rect 18144 14070 18196 14076
rect 18248 14082 18276 21126
rect 18432 20798 18460 22055
rect 18604 21064 18656 21070
rect 18604 21006 18656 21012
rect 18616 20866 18644 21006
rect 18604 20860 18656 20866
rect 18604 20802 18656 20808
rect 18420 20792 18472 20798
rect 18420 20734 18472 20740
rect 18432 19778 18460 20734
rect 18420 19772 18472 19778
rect 18420 19714 18472 19720
rect 18696 19636 18748 19642
rect 18696 19578 18748 19584
rect 18708 19234 18736 19578
rect 18696 19228 18748 19234
rect 18696 19170 18748 19176
rect 18604 17868 18656 17874
rect 18604 17810 18656 17816
rect 18510 17632 18566 17641
rect 18510 17567 18512 17576
rect 18564 17567 18566 17576
rect 18512 17538 18564 17544
rect 18418 17496 18474 17505
rect 18418 17431 18420 17440
rect 18472 17431 18474 17440
rect 18420 17402 18472 17408
rect 18418 16952 18474 16961
rect 18418 16887 18420 16896
rect 18472 16887 18474 16896
rect 18420 16858 18472 16864
rect 18432 16786 18460 16858
rect 18420 16780 18472 16786
rect 18420 16722 18472 16728
rect 18524 16514 18552 17538
rect 18616 17398 18644 17810
rect 18604 17392 18656 17398
rect 18604 17334 18656 17340
rect 18616 17058 18644 17334
rect 18604 17052 18656 17058
rect 18604 16994 18656 17000
rect 18694 16816 18750 16825
rect 18694 16751 18750 16760
rect 18604 16712 18656 16718
rect 18604 16654 18656 16660
rect 18512 16508 18564 16514
rect 18512 16450 18564 16456
rect 18616 16378 18644 16654
rect 18708 16514 18736 16751
rect 18696 16508 18748 16514
rect 18696 16450 18748 16456
rect 18800 16394 18828 23551
rect 19064 20656 19116 20662
rect 19064 20598 19116 20604
rect 19076 20254 19104 20598
rect 19064 20248 19116 20254
rect 19064 20190 19116 20196
rect 18970 19672 19026 19681
rect 18970 19607 18972 19616
rect 19024 19607 19026 19616
rect 18972 19578 19024 19584
rect 18880 17256 18932 17262
rect 18880 17198 18932 17204
rect 19064 17256 19116 17262
rect 19064 17198 19116 17204
rect 18892 16514 18920 17198
rect 19076 16854 19104 17198
rect 19064 16848 19116 16854
rect 19064 16790 19116 16796
rect 19064 16712 19116 16718
rect 19064 16654 19116 16660
rect 18880 16508 18932 16514
rect 18880 16450 18932 16456
rect 19076 16417 19104 16654
rect 18604 16372 18656 16378
rect 18604 16314 18656 16320
rect 18708 16366 18828 16394
rect 19062 16408 19118 16417
rect 18418 15592 18474 15601
rect 18418 15527 18474 15536
rect 18432 14542 18460 15527
rect 18616 15426 18644 16314
rect 18708 15737 18736 16366
rect 19062 16343 19118 16352
rect 18788 16236 18840 16242
rect 18788 16178 18840 16184
rect 18694 15728 18750 15737
rect 18694 15663 18750 15672
rect 18696 15624 18748 15630
rect 18696 15566 18748 15572
rect 18604 15420 18656 15426
rect 18604 15362 18656 15368
rect 18420 14536 18472 14542
rect 18420 14478 18472 14484
rect 18708 14241 18736 15566
rect 18800 15426 18828 16178
rect 18880 15692 18932 15698
rect 18880 15634 18932 15640
rect 18788 15420 18840 15426
rect 18788 15362 18840 15368
rect 18788 15216 18840 15222
rect 18788 15158 18840 15164
rect 18800 14610 18828 15158
rect 18892 14882 18920 15634
rect 18972 15624 19024 15630
rect 18972 15566 19024 15572
rect 18880 14876 18932 14882
rect 18880 14818 18932 14824
rect 18788 14604 18840 14610
rect 18788 14546 18840 14552
rect 18694 14232 18750 14241
rect 18694 14167 18750 14176
rect 18052 13788 18104 13794
rect 18052 13730 18104 13736
rect 17960 13720 18012 13726
rect 17960 13662 18012 13668
rect 16948 13584 17000 13590
rect 16948 13526 17000 13532
rect 16960 13182 16988 13526
rect 16948 13176 17000 13182
rect 16948 13118 17000 13124
rect 16672 13108 16724 13114
rect 16672 13050 16724 13056
rect 16684 12638 16712 13050
rect 16672 12632 16724 12638
rect 16672 12574 16724 12580
rect 16764 12156 16816 12162
rect 16764 12098 16816 12104
rect 16776 11414 16804 12098
rect 16764 11408 16816 11414
rect 16764 11350 16816 11356
rect 16776 11074 16804 11350
rect 16764 11068 16816 11074
rect 16764 11010 16816 11016
rect 17774 7296 17830 7305
rect 17774 7231 17776 7240
rect 17828 7231 17830 7240
rect 17776 7202 17828 7208
rect 16500 6178 16620 6194
rect 16488 6172 16620 6178
rect 16540 6166 16620 6172
rect 16488 6114 16540 6120
rect 16854 5936 16910 5945
rect 16854 5871 16856 5880
rect 16908 5871 16910 5880
rect 16856 5842 16908 5848
rect 16212 5084 16264 5090
rect 16212 5026 16264 5032
rect 15934 4848 15990 4857
rect 15934 4783 15936 4792
rect 15988 4783 15990 4792
rect 15936 4754 15988 4760
rect 10289 4644 10585 4664
rect 10345 4642 10369 4644
rect 10425 4642 10449 4644
rect 10505 4642 10529 4644
rect 10367 4590 10369 4642
rect 10431 4590 10443 4642
rect 10505 4590 10507 4642
rect 10345 4588 10369 4590
rect 10425 4588 10449 4590
rect 10505 4588 10529 4590
rect 10289 4568 10585 4588
rect 17972 4313 18000 13662
rect 18156 13590 18184 14070
rect 18248 14054 18736 14082
rect 18144 13584 18196 13590
rect 18144 13526 18196 13532
rect 18052 13040 18104 13046
rect 18052 12982 18104 12988
rect 18064 12706 18092 12982
rect 18052 12700 18104 12706
rect 18052 12642 18104 12648
rect 18064 12502 18092 12642
rect 18052 12496 18104 12502
rect 18052 12438 18104 12444
rect 18052 12020 18104 12026
rect 18052 11962 18104 11968
rect 18064 11278 18092 11962
rect 18156 11958 18184 13526
rect 18604 12564 18656 12570
rect 18604 12506 18656 12512
rect 18144 11952 18196 11958
rect 18144 11894 18196 11900
rect 18156 11618 18184 11894
rect 18616 11618 18644 12506
rect 18144 11612 18196 11618
rect 18144 11554 18196 11560
rect 18604 11612 18656 11618
rect 18604 11554 18656 11560
rect 18052 11272 18104 11278
rect 18052 11214 18104 11220
rect 18064 11074 18092 11214
rect 18052 11068 18104 11074
rect 18052 11010 18104 11016
rect 18708 7305 18736 14054
rect 18984 13794 19012 15566
rect 19062 14776 19118 14785
rect 19062 14711 19064 14720
rect 19116 14711 19118 14720
rect 19064 14682 19116 14688
rect 18972 13788 19024 13794
rect 18972 13730 19024 13736
rect 18878 13688 18934 13697
rect 18878 13623 18934 13632
rect 18892 13522 18920 13623
rect 18880 13516 18932 13522
rect 18880 13458 18932 13464
rect 18892 13250 18920 13458
rect 18880 13244 18932 13250
rect 18880 13186 18932 13192
rect 18972 11408 19024 11414
rect 18972 11350 19024 11356
rect 18984 11006 19012 11350
rect 18972 11000 19024 11006
rect 18972 10942 19024 10948
rect 19168 7577 19196 24474
rect 19248 23988 19300 23994
rect 19248 23930 19300 23936
rect 19260 23058 19288 23930
rect 19352 23314 19380 27240
rect 20088 27138 20116 27240
rect 20088 27110 20300 27138
rect 19622 25316 19918 25336
rect 19678 25314 19702 25316
rect 19758 25314 19782 25316
rect 19838 25314 19862 25316
rect 19700 25262 19702 25314
rect 19764 25262 19776 25314
rect 19838 25262 19840 25314
rect 19678 25260 19702 25262
rect 19758 25260 19782 25262
rect 19838 25260 19862 25262
rect 19622 25240 19918 25260
rect 19622 24228 19918 24248
rect 19678 24226 19702 24228
rect 19758 24226 19782 24228
rect 19838 24226 19862 24228
rect 19700 24174 19702 24226
rect 19764 24174 19776 24226
rect 19838 24174 19840 24226
rect 19678 24172 19702 24174
rect 19758 24172 19782 24174
rect 19838 24172 19862 24174
rect 19622 24152 19918 24172
rect 19982 23888 20038 23897
rect 19432 23852 19484 23858
rect 19982 23823 19984 23832
rect 19432 23794 19484 23800
rect 20036 23823 20038 23832
rect 19984 23794 20036 23800
rect 19444 23382 19472 23794
rect 19996 23586 20024 23794
rect 19984 23580 20036 23586
rect 19984 23522 20036 23528
rect 19432 23376 19484 23382
rect 19432 23318 19484 23324
rect 19340 23308 19392 23314
rect 19340 23250 19392 23256
rect 19260 23030 19380 23058
rect 19444 23042 19472 23318
rect 19622 23140 19918 23160
rect 19678 23138 19702 23140
rect 19758 23138 19782 23140
rect 19838 23138 19862 23140
rect 19700 23086 19702 23138
rect 19764 23086 19776 23138
rect 19838 23086 19840 23138
rect 19678 23084 19702 23086
rect 19758 23084 19782 23086
rect 19838 23084 19862 23086
rect 19622 23064 19918 23084
rect 19352 22974 19380 23030
rect 19432 23036 19484 23042
rect 19432 22978 19484 22984
rect 19340 22968 19392 22974
rect 19340 22910 19392 22916
rect 19622 22052 19918 22072
rect 19678 22050 19702 22052
rect 19758 22050 19782 22052
rect 19838 22050 19862 22052
rect 19700 21998 19702 22050
rect 19764 21998 19776 22050
rect 19838 21998 19840 22050
rect 19678 21996 19702 21998
rect 19758 21996 19782 21998
rect 19838 21996 19862 21998
rect 19622 21976 19918 21996
rect 19984 21880 20036 21886
rect 19984 21822 20036 21828
rect 19996 21410 20024 21822
rect 20168 21744 20220 21750
rect 20168 21686 20220 21692
rect 19984 21404 20036 21410
rect 19984 21346 20036 21352
rect 19248 21268 19300 21274
rect 19248 21210 19300 21216
rect 19260 20338 19288 21210
rect 20180 21070 20208 21686
rect 20168 21064 20220 21070
rect 20168 21006 20220 21012
rect 19622 20964 19918 20984
rect 19678 20962 19702 20964
rect 19758 20962 19782 20964
rect 19838 20962 19862 20964
rect 19700 20910 19702 20962
rect 19764 20910 19776 20962
rect 19838 20910 19840 20962
rect 19678 20908 19702 20910
rect 19758 20908 19782 20910
rect 19838 20908 19862 20910
rect 19622 20888 19918 20908
rect 20180 20662 20208 21006
rect 20168 20656 20220 20662
rect 20168 20598 20220 20604
rect 19260 20322 19380 20338
rect 19260 20316 19392 20322
rect 19260 20310 19340 20316
rect 19340 20258 19392 20264
rect 20180 20050 20208 20598
rect 19248 20044 19300 20050
rect 19248 19986 19300 19992
rect 20168 20044 20220 20050
rect 20168 19986 20220 19992
rect 19260 17618 19288 19986
rect 19622 19876 19918 19896
rect 19678 19874 19702 19876
rect 19758 19874 19782 19876
rect 19838 19874 19862 19876
rect 19700 19822 19702 19874
rect 19764 19822 19776 19874
rect 19838 19822 19840 19874
rect 19678 19820 19702 19822
rect 19758 19820 19782 19822
rect 19838 19820 19862 19822
rect 19622 19800 19918 19820
rect 19622 18788 19918 18808
rect 19678 18786 19702 18788
rect 19758 18786 19782 18788
rect 19838 18786 19862 18788
rect 19700 18734 19702 18786
rect 19764 18734 19776 18786
rect 19838 18734 19840 18786
rect 19678 18732 19702 18734
rect 19758 18732 19782 18734
rect 19838 18732 19862 18734
rect 19622 18712 19918 18732
rect 19432 18344 19484 18350
rect 19432 18286 19484 18292
rect 19444 17874 19472 18286
rect 19432 17868 19484 17874
rect 19432 17810 19484 17816
rect 19260 17590 19380 17618
rect 19352 17466 19380 17590
rect 19340 17460 19392 17466
rect 19340 17402 19392 17408
rect 19352 17058 19380 17402
rect 19444 17398 19472 17810
rect 19984 17800 20036 17806
rect 19984 17742 20036 17748
rect 19622 17700 19918 17720
rect 19678 17698 19702 17700
rect 19758 17698 19782 17700
rect 19838 17698 19862 17700
rect 19700 17646 19702 17698
rect 19764 17646 19776 17698
rect 19838 17646 19840 17698
rect 19678 17644 19702 17646
rect 19758 17644 19782 17646
rect 19838 17644 19862 17646
rect 19622 17624 19918 17644
rect 19892 17460 19944 17466
rect 19996 17448 20024 17742
rect 19944 17420 20024 17448
rect 19892 17402 19944 17408
rect 19432 17392 19484 17398
rect 19432 17334 19484 17340
rect 19340 17052 19392 17058
rect 19340 16994 19392 17000
rect 19904 16786 19932 17402
rect 20272 16972 20300 27110
rect 20732 24470 20760 27240
rect 21376 24538 21404 27240
rect 21364 24532 21416 24538
rect 21364 24474 21416 24480
rect 22008 24532 22060 24538
rect 22008 24474 22060 24480
rect 20720 24464 20772 24470
rect 20720 24406 20772 24412
rect 21640 24464 21692 24470
rect 21640 24406 21692 24412
rect 21088 23988 21140 23994
rect 21088 23930 21140 23936
rect 20536 23784 20588 23790
rect 20536 23726 20588 23732
rect 20548 23450 20576 23726
rect 20536 23444 20588 23450
rect 20536 23386 20588 23392
rect 20536 23308 20588 23314
rect 20536 23250 20588 23256
rect 20352 22900 20404 22906
rect 20352 22842 20404 22848
rect 20364 22498 20392 22842
rect 20444 22696 20496 22702
rect 20444 22638 20496 22644
rect 20352 22492 20404 22498
rect 20352 22434 20404 22440
rect 20456 22294 20484 22638
rect 20444 22288 20496 22294
rect 20444 22230 20496 22236
rect 20456 21886 20484 22230
rect 20444 21880 20496 21886
rect 20444 21822 20496 21828
rect 20548 21426 20576 23250
rect 20720 23240 20772 23246
rect 20640 23200 20720 23228
rect 20640 22362 20668 23200
rect 20720 23182 20772 23188
rect 20996 22832 21048 22838
rect 20996 22774 21048 22780
rect 21008 22537 21036 22774
rect 20994 22528 21050 22537
rect 20994 22463 20996 22472
rect 21048 22463 21050 22472
rect 20996 22434 21048 22440
rect 21008 22403 21036 22434
rect 20628 22356 20680 22362
rect 20628 22298 20680 22304
rect 20718 22256 20774 22265
rect 20718 22191 20720 22200
rect 20772 22191 20774 22200
rect 20720 22162 20772 22168
rect 20904 22152 20956 22158
rect 20904 22094 20956 22100
rect 20548 21398 20668 21426
rect 20536 21268 20588 21274
rect 20536 21210 20588 21216
rect 20548 20798 20576 21210
rect 20536 20792 20588 20798
rect 20536 20734 20588 20740
rect 20548 20322 20576 20734
rect 20536 20316 20588 20322
rect 20536 20258 20588 20264
rect 20536 18480 20588 18486
rect 20536 18422 20588 18428
rect 20548 17058 20576 18422
rect 20536 17052 20588 17058
rect 20536 16994 20588 17000
rect 20272 16944 20484 16972
rect 19340 16780 19392 16786
rect 19340 16722 19392 16728
rect 19892 16780 19944 16786
rect 19892 16722 19944 16728
rect 19352 16310 19380 16722
rect 19622 16612 19918 16632
rect 19678 16610 19702 16612
rect 19758 16610 19782 16612
rect 19838 16610 19862 16612
rect 19700 16558 19702 16610
rect 19764 16558 19776 16610
rect 19838 16558 19840 16610
rect 19678 16556 19702 16558
rect 19758 16556 19782 16558
rect 19838 16556 19862 16558
rect 19622 16536 19918 16556
rect 19432 16508 19484 16514
rect 19432 16450 19484 16456
rect 19340 16304 19392 16310
rect 19340 16246 19392 16252
rect 19444 15970 19472 16450
rect 19432 15964 19484 15970
rect 19432 15906 19484 15912
rect 19248 15828 19300 15834
rect 19248 15770 19300 15776
rect 19260 15358 19288 15770
rect 20352 15692 20404 15698
rect 20352 15634 20404 15640
rect 19622 15524 19918 15544
rect 19678 15522 19702 15524
rect 19758 15522 19782 15524
rect 19838 15522 19862 15524
rect 19700 15470 19702 15522
rect 19764 15470 19776 15522
rect 19838 15470 19840 15522
rect 19678 15468 19702 15470
rect 19758 15468 19782 15470
rect 19838 15468 19862 15470
rect 19622 15448 19918 15468
rect 20364 15426 20392 15634
rect 20352 15420 20404 15426
rect 20352 15362 20404 15368
rect 19248 15352 19300 15358
rect 19248 15294 19300 15300
rect 19260 15034 19288 15294
rect 19260 15006 19380 15034
rect 19352 14882 19380 15006
rect 19340 14876 19392 14882
rect 19340 14818 19392 14824
rect 19248 14536 19300 14542
rect 19248 14478 19300 14484
rect 19260 13153 19288 14478
rect 19352 14338 19380 14818
rect 19524 14740 19576 14746
rect 19524 14682 19576 14688
rect 19340 14332 19392 14338
rect 19340 14274 19392 14280
rect 19536 14202 19564 14682
rect 19622 14436 19918 14456
rect 19678 14434 19702 14436
rect 19758 14434 19782 14436
rect 19838 14434 19862 14436
rect 19700 14382 19702 14434
rect 19764 14382 19776 14434
rect 19838 14382 19840 14434
rect 19678 14380 19702 14382
rect 19758 14380 19782 14382
rect 19838 14380 19862 14382
rect 19622 14360 19918 14380
rect 19524 14196 19576 14202
rect 19524 14138 19576 14144
rect 19536 13794 19564 14138
rect 20258 13824 20314 13833
rect 19524 13788 19576 13794
rect 20258 13759 20260 13768
rect 19524 13730 19576 13736
rect 20312 13759 20314 13768
rect 20260 13730 20312 13736
rect 19622 13348 19918 13368
rect 19678 13346 19702 13348
rect 19758 13346 19782 13348
rect 19838 13346 19862 13348
rect 19700 13294 19702 13346
rect 19764 13294 19776 13346
rect 19838 13294 19840 13346
rect 19678 13292 19702 13294
rect 19758 13292 19782 13294
rect 19838 13292 19862 13294
rect 19622 13272 19918 13292
rect 19246 13144 19302 13153
rect 19246 13079 19302 13088
rect 19616 13108 19668 13114
rect 19616 13050 19668 13056
rect 19892 13108 19944 13114
rect 19892 13050 19944 13056
rect 19628 12706 19656 13050
rect 19616 12700 19668 12706
rect 19616 12642 19668 12648
rect 19904 12502 19932 13050
rect 19524 12496 19576 12502
rect 19524 12438 19576 12444
rect 19892 12496 19944 12502
rect 19892 12438 19944 12444
rect 19536 12162 19564 12438
rect 19622 12260 19918 12280
rect 19678 12258 19702 12260
rect 19758 12258 19782 12260
rect 19838 12258 19862 12260
rect 19700 12206 19702 12258
rect 19764 12206 19776 12258
rect 19838 12206 19840 12258
rect 19678 12204 19702 12206
rect 19758 12204 19782 12206
rect 19838 12204 19862 12206
rect 19622 12184 19918 12204
rect 19524 12156 19576 12162
rect 19524 12098 19576 12104
rect 19246 11512 19302 11521
rect 19246 11447 19302 11456
rect 19432 11476 19484 11482
rect 19260 11414 19288 11447
rect 19432 11418 19484 11424
rect 19248 11408 19300 11414
rect 19248 11350 19300 11356
rect 19248 11272 19300 11278
rect 19248 11214 19300 11220
rect 19154 7568 19210 7577
rect 19154 7503 19210 7512
rect 18694 7296 18750 7305
rect 18694 7231 18750 7240
rect 18234 7160 18290 7169
rect 18234 7095 18236 7104
rect 18288 7095 18290 7104
rect 18236 7066 18288 7072
rect 19260 5401 19288 11214
rect 19444 11074 19472 11418
rect 19622 11172 19918 11192
rect 19678 11170 19702 11172
rect 19758 11170 19782 11172
rect 19838 11170 19862 11172
rect 19700 11118 19702 11170
rect 19764 11118 19776 11170
rect 19838 11118 19840 11170
rect 19678 11116 19702 11118
rect 19758 11116 19782 11118
rect 19838 11116 19862 11118
rect 19622 11096 19918 11116
rect 19432 11068 19484 11074
rect 19432 11010 19484 11016
rect 19622 10084 19918 10104
rect 19678 10082 19702 10084
rect 19758 10082 19782 10084
rect 19838 10082 19862 10084
rect 19700 10030 19702 10082
rect 19764 10030 19776 10082
rect 19838 10030 19840 10082
rect 19678 10028 19702 10030
rect 19758 10028 19782 10030
rect 19838 10028 19862 10030
rect 19622 10008 19918 10028
rect 20456 9345 20484 16944
rect 20442 9336 20498 9345
rect 20442 9271 20498 9280
rect 20640 9073 20668 21398
rect 20916 21206 20944 22094
rect 20904 21200 20956 21206
rect 20904 21142 20956 21148
rect 20996 21132 21048 21138
rect 20996 21074 21048 21080
rect 20904 21064 20956 21070
rect 20904 21006 20956 21012
rect 20916 20769 20944 21006
rect 20902 20760 20958 20769
rect 20902 20695 20958 20704
rect 20812 20520 20864 20526
rect 20812 20462 20864 20468
rect 20824 20254 20852 20462
rect 20812 20248 20864 20254
rect 20812 20190 20864 20196
rect 21008 20186 21036 21074
rect 20996 20180 21048 20186
rect 20996 20122 21048 20128
rect 20996 19432 21048 19438
rect 20996 19374 21048 19380
rect 21008 19098 21036 19374
rect 20996 19092 21048 19098
rect 20996 19034 21048 19040
rect 20720 18888 20772 18894
rect 20720 18830 20772 18836
rect 20732 18457 20760 18830
rect 21008 18690 21036 19034
rect 20996 18684 21048 18690
rect 20996 18626 21048 18632
rect 20904 18480 20956 18486
rect 20718 18448 20774 18457
rect 20904 18422 20956 18428
rect 20718 18383 20774 18392
rect 20916 17942 20944 18422
rect 21008 17942 21036 18626
rect 20904 17936 20956 17942
rect 20904 17878 20956 17884
rect 20996 17936 21048 17942
rect 20996 17878 21048 17884
rect 20720 17800 20772 17806
rect 20720 17742 20772 17748
rect 20732 17534 20760 17742
rect 21008 17602 21036 17878
rect 20996 17596 21048 17602
rect 20996 17538 21048 17544
rect 20720 17528 20772 17534
rect 20720 17470 20772 17476
rect 20732 15834 20760 17470
rect 20720 15828 20772 15834
rect 20720 15770 20772 15776
rect 20732 15290 20760 15770
rect 20720 15284 20772 15290
rect 20720 15226 20772 15232
rect 20718 14776 20774 14785
rect 20718 14711 20720 14720
rect 20772 14711 20774 14720
rect 20720 14682 20772 14688
rect 20904 14536 20956 14542
rect 20904 14478 20956 14484
rect 20812 14196 20864 14202
rect 20812 14138 20864 14144
rect 20824 13726 20852 14138
rect 20812 13720 20864 13726
rect 20916 13697 20944 14478
rect 21100 14270 21128 23930
rect 21456 23852 21508 23858
rect 21456 23794 21508 23800
rect 21468 23450 21496 23794
rect 21456 23444 21508 23450
rect 21456 23386 21508 23392
rect 21180 22968 21232 22974
rect 21180 22910 21232 22916
rect 21192 22158 21220 22910
rect 21364 22900 21416 22906
rect 21364 22842 21416 22848
rect 21376 22537 21404 22842
rect 21362 22528 21418 22537
rect 21362 22463 21418 22472
rect 21180 22152 21232 22158
rect 21180 22094 21232 22100
rect 21548 21608 21600 21614
rect 21548 21550 21600 21556
rect 21560 21274 21588 21550
rect 21548 21268 21600 21274
rect 21548 21210 21600 21216
rect 21548 19432 21600 19438
rect 21548 19374 21600 19380
rect 21560 19273 21588 19374
rect 21546 19264 21602 19273
rect 21546 19199 21602 19208
rect 21272 18888 21324 18894
rect 21456 18888 21508 18894
rect 21324 18848 21404 18876
rect 21272 18830 21324 18836
rect 21376 18350 21404 18848
rect 21456 18830 21508 18836
rect 21468 18554 21496 18830
rect 21456 18548 21508 18554
rect 21456 18490 21508 18496
rect 21364 18344 21416 18350
rect 21364 18286 21416 18292
rect 21178 17360 21234 17369
rect 21178 17295 21234 17304
rect 21192 16446 21220 17295
rect 21180 16440 21232 16446
rect 21180 16382 21232 16388
rect 21192 15970 21220 16382
rect 21272 16304 21324 16310
rect 21272 16246 21324 16252
rect 21180 15964 21232 15970
rect 21180 15906 21232 15912
rect 21284 15698 21312 16246
rect 21272 15692 21324 15698
rect 21272 15634 21324 15640
rect 21272 15284 21324 15290
rect 21272 15226 21324 15232
rect 21284 14882 21312 15226
rect 21376 15057 21404 18286
rect 21560 16378 21588 19199
rect 21652 18978 21680 24406
rect 21732 22152 21784 22158
rect 21732 22094 21784 22100
rect 21643 18950 21680 18978
rect 21643 18865 21671 18950
rect 21638 18856 21694 18865
rect 21638 18791 21694 18800
rect 21744 17505 21772 22094
rect 21822 17768 21878 17777
rect 21822 17703 21878 17712
rect 21836 17602 21864 17703
rect 21824 17596 21876 17602
rect 21824 17538 21876 17544
rect 21730 17496 21786 17505
rect 21730 17431 21786 17440
rect 21744 16786 21772 17431
rect 21732 16780 21784 16786
rect 21732 16722 21784 16728
rect 21916 16712 21968 16718
rect 21916 16654 21968 16660
rect 21928 16553 21956 16654
rect 21914 16544 21970 16553
rect 21914 16479 21970 16488
rect 21548 16372 21600 16378
rect 21548 16314 21600 16320
rect 21560 15630 21588 16314
rect 21732 15692 21784 15698
rect 21732 15634 21784 15640
rect 21548 15624 21600 15630
rect 21548 15566 21600 15572
rect 21362 15048 21418 15057
rect 21362 14983 21418 14992
rect 21272 14876 21324 14882
rect 21272 14818 21324 14824
rect 21088 14264 21140 14270
rect 21088 14206 21140 14212
rect 20812 13662 20864 13668
rect 20902 13688 20958 13697
rect 20902 13623 20958 13632
rect 20812 13584 20864 13590
rect 20812 13526 20864 13532
rect 20824 12162 20852 13526
rect 21284 13182 21312 14818
rect 21272 13176 21324 13182
rect 21272 13118 21324 13124
rect 21364 12904 21416 12910
rect 21364 12846 21416 12852
rect 21376 12434 21404 12846
rect 21364 12428 21416 12434
rect 21364 12370 21416 12376
rect 20812 12156 20864 12162
rect 20812 12098 20864 12104
rect 21180 12020 21232 12026
rect 21180 11962 21232 11968
rect 21192 11414 21220 11962
rect 21376 11958 21404 12370
rect 21456 12020 21508 12026
rect 21456 11962 21508 11968
rect 21364 11952 21416 11958
rect 21364 11894 21416 11900
rect 21376 11618 21404 11894
rect 21468 11618 21496 11962
rect 21364 11612 21416 11618
rect 21364 11554 21416 11560
rect 21456 11612 21508 11618
rect 21456 11554 21508 11560
rect 21468 11521 21496 11554
rect 21454 11512 21510 11521
rect 21454 11447 21510 11456
rect 21180 11408 21232 11414
rect 21178 11376 21180 11385
rect 21232 11376 21234 11385
rect 21178 11311 21234 11320
rect 20626 9064 20682 9073
rect 19622 8996 19918 9016
rect 20626 8999 20682 9008
rect 19678 8994 19702 8996
rect 19758 8994 19782 8996
rect 19838 8994 19862 8996
rect 19700 8942 19702 8994
rect 19764 8942 19776 8994
rect 19838 8942 19840 8994
rect 19678 8940 19702 8942
rect 19758 8940 19782 8942
rect 19838 8940 19862 8942
rect 19622 8920 19918 8940
rect 19622 7908 19918 7928
rect 19678 7906 19702 7908
rect 19758 7906 19782 7908
rect 19838 7906 19862 7908
rect 19700 7854 19702 7906
rect 19764 7854 19776 7906
rect 19838 7854 19840 7906
rect 19678 7852 19702 7854
rect 19758 7852 19782 7854
rect 19838 7852 19862 7854
rect 19622 7832 19918 7852
rect 19622 6820 19918 6840
rect 19678 6818 19702 6820
rect 19758 6818 19782 6820
rect 19838 6818 19862 6820
rect 19700 6766 19702 6818
rect 19764 6766 19776 6818
rect 19838 6766 19840 6818
rect 19678 6764 19702 6766
rect 19758 6764 19782 6766
rect 19838 6764 19862 6766
rect 19622 6744 19918 6764
rect 19622 5732 19918 5752
rect 19678 5730 19702 5732
rect 19758 5730 19782 5732
rect 19838 5730 19862 5732
rect 19700 5678 19702 5730
rect 19764 5678 19776 5730
rect 19838 5678 19840 5730
rect 19678 5676 19702 5678
rect 19758 5676 19782 5678
rect 19838 5676 19862 5678
rect 19622 5656 19918 5676
rect 19246 5392 19302 5401
rect 19246 5327 19302 5336
rect 21560 4993 21588 15566
rect 21744 15290 21772 15634
rect 21732 15284 21784 15290
rect 21732 15226 21784 15232
rect 21744 14882 21772 15226
rect 21732 14876 21784 14882
rect 21732 14818 21784 14824
rect 21824 13516 21876 13522
rect 21824 13458 21876 13464
rect 21836 13250 21864 13458
rect 21824 13244 21876 13250
rect 21824 13186 21876 13192
rect 22020 10569 22048 24474
rect 22112 23738 22140 27240
rect 22560 24464 22612 24470
rect 22558 24432 22560 24441
rect 22612 24432 22614 24441
rect 22558 24367 22614 24376
rect 22756 24130 22784 27240
rect 22836 25076 22888 25082
rect 22836 25018 22888 25024
rect 22848 24606 22876 25018
rect 22836 24600 22888 24606
rect 22834 24568 22836 24577
rect 22888 24568 22890 24577
rect 22834 24503 22890 24512
rect 22848 24477 22876 24503
rect 22744 24124 22796 24130
rect 22744 24066 22796 24072
rect 22284 23988 22336 23994
rect 22284 23930 22336 23936
rect 22112 23710 22232 23738
rect 22098 23616 22154 23625
rect 22098 23551 22154 23560
rect 22112 23518 22140 23551
rect 22100 23512 22152 23518
rect 22100 23454 22152 23460
rect 22204 20866 22232 23710
rect 22296 22673 22324 23930
rect 22836 23444 22888 23450
rect 22836 23386 22888 23392
rect 22374 23344 22430 23353
rect 22374 23279 22376 23288
rect 22428 23279 22430 23288
rect 22376 23250 22428 23256
rect 22848 22702 22876 23386
rect 22468 22696 22520 22702
rect 22282 22664 22338 22673
rect 22468 22638 22520 22644
rect 22836 22696 22888 22702
rect 22836 22638 22888 22644
rect 22282 22599 22338 22608
rect 22480 22362 22508 22638
rect 22468 22356 22520 22362
rect 22468 22298 22520 22304
rect 22848 22226 22876 22638
rect 23216 22498 23244 27359
rect 23478 27240 23534 27720
rect 24122 27240 24178 27720
rect 24766 27240 24822 27720
rect 25502 27240 25558 27720
rect 26146 27240 26202 27720
rect 26882 27240 26938 27720
rect 27526 27240 27582 27720
rect 23386 26200 23442 26209
rect 23386 26135 23442 26144
rect 23294 25656 23350 25665
rect 23294 25591 23350 25600
rect 23308 23858 23336 25591
rect 23400 24334 23428 26135
rect 23388 24328 23440 24334
rect 23388 24270 23440 24276
rect 23296 23852 23348 23858
rect 23296 23794 23348 23800
rect 23204 22492 23256 22498
rect 23204 22434 23256 22440
rect 22836 22220 22888 22226
rect 22836 22162 22888 22168
rect 23388 22220 23440 22226
rect 23388 22162 23440 22168
rect 22926 21712 22982 21721
rect 22926 21647 22982 21656
rect 22940 21410 22968 21647
rect 23400 21614 23428 22162
rect 23388 21608 23440 21614
rect 23492 21596 23520 27240
rect 23570 26880 23626 26889
rect 23570 26815 23626 26824
rect 23584 25218 23612 26815
rect 23572 25212 23624 25218
rect 23572 25154 23624 25160
rect 23756 24532 23808 24538
rect 24136 24520 24164 27240
rect 24780 25370 24808 27240
rect 24688 25342 24808 25370
rect 24289 24772 24585 24792
rect 24345 24770 24369 24772
rect 24425 24770 24449 24772
rect 24505 24770 24529 24772
rect 24367 24718 24369 24770
rect 24431 24718 24443 24770
rect 24505 24718 24507 24770
rect 24345 24716 24369 24718
rect 24425 24716 24449 24718
rect 24505 24716 24529 24718
rect 24289 24696 24585 24716
rect 24688 24538 24716 25342
rect 24768 25212 24820 25218
rect 24768 25154 24820 25160
rect 24780 25121 24808 25154
rect 24766 25112 24822 25121
rect 24766 25047 24822 25056
rect 24768 25008 24820 25014
rect 24768 24950 24820 24956
rect 23756 24474 23808 24480
rect 24044 24492 24164 24520
rect 24676 24532 24728 24538
rect 23664 23988 23716 23994
rect 23664 23930 23716 23936
rect 23676 23586 23704 23930
rect 23664 23580 23716 23586
rect 23664 23522 23716 23528
rect 23664 23376 23716 23382
rect 23664 23318 23716 23324
rect 23572 23240 23624 23246
rect 23572 23182 23624 23188
rect 23584 23042 23612 23182
rect 23572 23036 23624 23042
rect 23572 22978 23624 22984
rect 23492 21568 23612 21596
rect 23388 21550 23440 21556
rect 23400 21426 23428 21550
rect 22928 21404 22980 21410
rect 23400 21398 23520 21426
rect 22928 21346 22980 21352
rect 22192 20860 22244 20866
rect 22192 20802 22244 20808
rect 22836 20520 22888 20526
rect 22836 20462 22888 20468
rect 22848 20118 22876 20462
rect 23492 20322 23520 21398
rect 23480 20316 23532 20322
rect 23480 20258 23532 20264
rect 22560 20112 22612 20118
rect 22560 20054 22612 20060
rect 22836 20112 22888 20118
rect 22836 20054 22888 20060
rect 23480 20112 23532 20118
rect 23480 20054 23532 20060
rect 22572 19574 22600 20054
rect 22652 19976 22704 19982
rect 22652 19918 22704 19924
rect 22100 19568 22152 19574
rect 22100 19510 22152 19516
rect 22560 19568 22612 19574
rect 22560 19510 22612 19516
rect 22112 19166 22140 19510
rect 22100 19160 22152 19166
rect 22098 19128 22100 19137
rect 22152 19128 22154 19137
rect 22098 19063 22154 19072
rect 22572 19030 22600 19510
rect 22664 19098 22692 19918
rect 22848 19574 22876 20054
rect 22836 19568 22888 19574
rect 22836 19510 22888 19516
rect 22652 19092 22704 19098
rect 22652 19034 22704 19040
rect 22100 19024 22152 19030
rect 22100 18966 22152 18972
rect 22560 19024 22612 19030
rect 22560 18966 22612 18972
rect 22112 17602 22140 18966
rect 22572 18690 22600 18966
rect 23294 18856 23350 18865
rect 23294 18791 23350 18800
rect 22560 18684 22612 18690
rect 22560 18626 22612 18632
rect 22192 18548 22244 18554
rect 22192 18490 22244 18496
rect 22204 18146 22232 18490
rect 22192 18140 22244 18146
rect 22192 18082 22244 18088
rect 22376 18140 22428 18146
rect 22376 18082 22428 18088
rect 22100 17596 22152 17602
rect 22100 17538 22152 17544
rect 22112 16990 22140 17538
rect 22192 17460 22244 17466
rect 22192 17402 22244 17408
rect 22204 17058 22232 17402
rect 22388 17398 22416 18082
rect 22376 17392 22428 17398
rect 22376 17334 22428 17340
rect 22192 17052 22244 17058
rect 22192 16994 22244 17000
rect 22100 16984 22152 16990
rect 22100 16926 22152 16932
rect 22284 16916 22336 16922
rect 22284 16858 22336 16864
rect 22190 16408 22246 16417
rect 22190 16343 22246 16352
rect 22204 14542 22232 16343
rect 22296 16310 22324 16858
rect 22388 16802 22416 17334
rect 22388 16774 22508 16802
rect 22376 16712 22428 16718
rect 22376 16654 22428 16660
rect 22388 16514 22416 16654
rect 22376 16508 22428 16514
rect 22376 16450 22428 16456
rect 22480 16446 22508 16774
rect 22468 16440 22520 16446
rect 22468 16382 22520 16388
rect 22560 16372 22612 16378
rect 22560 16314 22612 16320
rect 22284 16304 22336 16310
rect 22284 16246 22336 16252
rect 22296 15766 22324 16246
rect 22284 15760 22336 15766
rect 22284 15702 22336 15708
rect 22296 15426 22324 15702
rect 22284 15420 22336 15426
rect 22284 15362 22336 15368
rect 22572 14678 22600 16314
rect 23020 15420 23072 15426
rect 23020 15362 23072 15368
rect 23032 14746 23060 15362
rect 23020 14740 23072 14746
rect 23020 14682 23072 14688
rect 22560 14672 22612 14678
rect 22560 14614 22612 14620
rect 22192 14536 22244 14542
rect 22192 14478 22244 14484
rect 22572 14338 22600 14614
rect 22928 14536 22980 14542
rect 22928 14478 22980 14484
rect 22560 14332 22612 14338
rect 22560 14274 22612 14280
rect 22100 13652 22152 13658
rect 22100 13594 22152 13600
rect 22112 12706 22140 13594
rect 22100 12700 22152 12706
rect 22100 12642 22152 12648
rect 22940 10705 22968 14478
rect 23032 14338 23060 14682
rect 23020 14332 23072 14338
rect 23020 14274 23072 14280
rect 22926 10696 22982 10705
rect 22926 10631 22982 10640
rect 22006 10560 22062 10569
rect 22006 10495 22062 10504
rect 23308 9986 23336 18791
rect 23492 16242 23520 20054
rect 23584 16310 23612 21568
rect 23676 21449 23704 23318
rect 23662 21440 23718 21449
rect 23662 21375 23718 21384
rect 23664 21064 23716 21070
rect 23664 21006 23716 21012
rect 23676 20633 23704 21006
rect 23662 20624 23718 20633
rect 23662 20559 23718 20568
rect 23768 20202 23796 24474
rect 23848 24464 23900 24470
rect 23848 24406 23900 24412
rect 23860 24334 23888 24406
rect 23848 24328 23900 24334
rect 23848 24270 23900 24276
rect 23860 22809 23888 24270
rect 23940 22832 23992 22838
rect 23846 22800 23902 22809
rect 23940 22774 23992 22780
rect 23846 22735 23902 22744
rect 23846 22664 23902 22673
rect 23846 22599 23902 22608
rect 23860 20882 23888 22599
rect 23952 22537 23980 22774
rect 23938 22528 23994 22537
rect 23938 22463 23940 22472
rect 23992 22463 23994 22472
rect 23940 22434 23992 22440
rect 23952 21886 23980 22434
rect 23940 21880 23992 21886
rect 23940 21822 23992 21828
rect 24044 21120 24072 24492
rect 24676 24474 24728 24480
rect 24216 24464 24268 24470
rect 24216 24406 24268 24412
rect 24228 24062 24256 24406
rect 24676 24396 24728 24402
rect 24676 24338 24728 24344
rect 24216 24056 24268 24062
rect 24216 23998 24268 24004
rect 24688 23994 24716 24338
rect 24780 24334 24808 24950
rect 25134 24432 25190 24441
rect 25134 24367 25190 24376
rect 25148 24334 25176 24367
rect 24768 24328 24820 24334
rect 24768 24270 24820 24276
rect 25136 24328 25188 24334
rect 25136 24270 25188 24276
rect 24676 23988 24728 23994
rect 24676 23930 24728 23936
rect 24216 23784 24268 23790
rect 24216 23726 24268 23732
rect 24228 23382 24256 23726
rect 24289 23684 24585 23704
rect 24345 23682 24369 23684
rect 24425 23682 24449 23684
rect 24505 23682 24529 23684
rect 24367 23630 24369 23682
rect 24431 23630 24443 23682
rect 24505 23630 24507 23682
rect 24345 23628 24369 23630
rect 24425 23628 24449 23630
rect 24505 23628 24529 23630
rect 24289 23608 24585 23628
rect 24688 23586 24716 23930
rect 24676 23580 24728 23586
rect 24676 23522 24728 23528
rect 24780 23450 24808 24270
rect 25134 23888 25190 23897
rect 25134 23823 25136 23832
rect 25188 23823 25190 23832
rect 25228 23852 25280 23858
rect 25136 23794 25188 23800
rect 25228 23794 25280 23800
rect 24768 23444 24820 23450
rect 24768 23386 24820 23392
rect 24216 23376 24268 23382
rect 24216 23318 24268 23324
rect 24124 23036 24176 23042
rect 24124 22978 24176 22984
rect 24136 22498 24164 22978
rect 24216 22968 24268 22974
rect 24216 22910 24268 22916
rect 24124 22492 24176 22498
rect 24124 22434 24176 22440
rect 24228 22158 24256 22910
rect 24860 22696 24912 22702
rect 24674 22664 24730 22673
rect 24289 22596 24585 22616
rect 24860 22638 24912 22644
rect 24674 22599 24730 22608
rect 24345 22594 24369 22596
rect 24425 22594 24449 22596
rect 24505 22594 24529 22596
rect 24367 22542 24369 22594
rect 24431 22542 24443 22594
rect 24505 22542 24507 22594
rect 24345 22540 24369 22542
rect 24425 22540 24449 22542
rect 24505 22540 24529 22542
rect 24289 22520 24585 22540
rect 24216 22152 24268 22158
rect 24216 22094 24268 22100
rect 24228 21954 24256 22094
rect 24216 21948 24268 21954
rect 24216 21890 24268 21896
rect 24124 21812 24176 21818
rect 24124 21754 24176 21760
rect 24136 21585 24164 21754
rect 24688 21721 24716 22599
rect 24766 22392 24822 22401
rect 24766 22327 24822 22336
rect 24780 22294 24808 22327
rect 24768 22288 24820 22294
rect 24768 22230 24820 22236
rect 24674 21712 24730 21721
rect 24674 21647 24730 21656
rect 24768 21608 24820 21614
rect 24122 21576 24178 21585
rect 24768 21550 24820 21556
rect 24122 21511 24178 21520
rect 24136 21410 24164 21511
rect 24289 21508 24585 21528
rect 24345 21506 24369 21508
rect 24425 21506 24449 21508
rect 24505 21506 24529 21508
rect 24367 21454 24369 21506
rect 24431 21454 24443 21506
rect 24505 21454 24507 21506
rect 24345 21452 24369 21454
rect 24425 21452 24449 21454
rect 24505 21452 24529 21454
rect 24289 21432 24585 21452
rect 24780 21449 24808 21550
rect 24766 21440 24822 21449
rect 24124 21404 24176 21410
rect 24766 21375 24822 21384
rect 24124 21346 24176 21352
rect 24044 21092 24256 21120
rect 23860 20854 23980 20882
rect 23846 20760 23902 20769
rect 23846 20695 23848 20704
rect 23900 20695 23902 20704
rect 23848 20666 23900 20672
rect 23860 20322 23888 20666
rect 23848 20316 23900 20322
rect 23848 20258 23900 20264
rect 23768 20174 23888 20202
rect 23664 19432 23716 19438
rect 23664 19374 23716 19380
rect 23676 18554 23704 19374
rect 23664 18548 23716 18554
rect 23664 18490 23716 18496
rect 23676 18146 23704 18490
rect 23754 18176 23810 18185
rect 23664 18140 23716 18146
rect 23754 18111 23810 18120
rect 23664 18082 23716 18088
rect 23664 17800 23716 17806
rect 23662 17768 23664 17777
rect 23716 17768 23718 17777
rect 23662 17703 23718 17712
rect 23664 16780 23716 16786
rect 23664 16722 23716 16728
rect 23572 16304 23624 16310
rect 23572 16246 23624 16252
rect 23480 16236 23532 16242
rect 23480 16178 23532 16184
rect 23676 15850 23704 16722
rect 23768 16378 23796 18111
rect 23756 16372 23808 16378
rect 23756 16314 23808 16320
rect 23768 15970 23796 16314
rect 23756 15964 23808 15970
rect 23756 15906 23808 15912
rect 23676 15822 23796 15850
rect 23664 15624 23716 15630
rect 23664 15566 23716 15572
rect 23676 15329 23704 15566
rect 23662 15320 23718 15329
rect 23480 15284 23532 15290
rect 23662 15255 23718 15264
rect 23480 15226 23532 15232
rect 23386 15048 23442 15057
rect 23386 14983 23442 14992
rect 23400 14218 23428 14983
rect 23492 14814 23520 15226
rect 23676 15222 23704 15255
rect 23664 15216 23716 15222
rect 23664 15158 23716 15164
rect 23664 15080 23716 15086
rect 23664 15022 23716 15028
rect 23480 14808 23532 14814
rect 23480 14750 23532 14756
rect 23492 14338 23520 14750
rect 23676 14678 23704 15022
rect 23664 14672 23716 14678
rect 23664 14614 23716 14620
rect 23480 14332 23532 14338
rect 23480 14274 23532 14280
rect 23662 14232 23718 14241
rect 23400 14190 23520 14218
rect 23492 12042 23520 14190
rect 23662 14167 23664 14176
rect 23716 14167 23718 14176
rect 23664 14138 23716 14144
rect 23676 13794 23704 14138
rect 23664 13788 23716 13794
rect 23664 13730 23716 13736
rect 23492 12014 23612 12042
rect 23296 9980 23348 9986
rect 23296 9922 23348 9928
rect 23478 6616 23534 6625
rect 23478 6551 23534 6560
rect 23492 5401 23520 6551
rect 23478 5392 23534 5401
rect 23478 5327 23534 5336
rect 21546 4984 21602 4993
rect 21546 4919 21602 4928
rect 23478 4712 23534 4721
rect 19622 4644 19918 4664
rect 23478 4647 23534 4656
rect 19678 4642 19702 4644
rect 19758 4642 19782 4644
rect 19838 4642 19862 4644
rect 19700 4590 19702 4642
rect 19764 4590 19776 4642
rect 19838 4590 19840 4642
rect 19678 4588 19702 4590
rect 19758 4588 19782 4590
rect 19838 4588 19862 4590
rect 19622 4568 19918 4588
rect 17958 4304 18014 4313
rect 17958 4239 18014 4248
rect 5622 4100 5918 4120
rect 5678 4098 5702 4100
rect 5758 4098 5782 4100
rect 5838 4098 5862 4100
rect 5700 4046 5702 4098
rect 5764 4046 5776 4098
rect 5838 4046 5840 4098
rect 5678 4044 5702 4046
rect 5758 4044 5782 4046
rect 5838 4044 5862 4046
rect 5622 4024 5918 4044
rect 14956 4100 15252 4120
rect 15012 4098 15036 4100
rect 15092 4098 15116 4100
rect 15172 4098 15196 4100
rect 15034 4046 15036 4098
rect 15098 4046 15110 4098
rect 15172 4046 15174 4098
rect 15012 4044 15036 4046
rect 15092 4044 15116 4046
rect 15172 4044 15196 4046
rect 14956 4024 15252 4044
rect 10289 3556 10585 3576
rect 10345 3554 10369 3556
rect 10425 3554 10449 3556
rect 10505 3554 10529 3556
rect 10367 3502 10369 3554
rect 10431 3502 10443 3554
rect 10505 3502 10507 3554
rect 10345 3500 10369 3502
rect 10425 3500 10449 3502
rect 10505 3500 10529 3502
rect 10289 3480 10585 3500
rect 19622 3556 19918 3576
rect 19678 3554 19702 3556
rect 19758 3554 19782 3556
rect 19838 3554 19862 3556
rect 19700 3502 19702 3554
rect 19764 3502 19776 3554
rect 19838 3502 19840 3554
rect 19678 3500 19702 3502
rect 19758 3500 19782 3502
rect 19838 3500 19862 3502
rect 19622 3480 19918 3500
rect 5622 3012 5918 3032
rect 5678 3010 5702 3012
rect 5758 3010 5782 3012
rect 5838 3010 5862 3012
rect 5700 2958 5702 3010
rect 5764 2958 5776 3010
rect 5838 2958 5840 3010
rect 5678 2956 5702 2958
rect 5758 2956 5782 2958
rect 5838 2956 5862 2958
rect 5622 2936 5918 2956
rect 14956 3012 15252 3032
rect 15012 3010 15036 3012
rect 15092 3010 15116 3012
rect 15172 3010 15196 3012
rect 15034 2958 15036 3010
rect 15098 2958 15110 3010
rect 15172 2958 15174 3010
rect 15012 2956 15036 2958
rect 15092 2956 15116 2958
rect 15172 2956 15196 2958
rect 14956 2936 15252 2956
rect 10289 2468 10585 2488
rect 10345 2466 10369 2468
rect 10425 2466 10449 2468
rect 10505 2466 10529 2468
rect 10367 2414 10369 2466
rect 10431 2414 10443 2466
rect 10505 2414 10507 2466
rect 10345 2412 10369 2414
rect 10425 2412 10449 2414
rect 10505 2412 10529 2414
rect 10289 2392 10585 2412
rect 19622 2468 19918 2488
rect 19678 2466 19702 2468
rect 19758 2466 19782 2468
rect 19838 2466 19862 2468
rect 19700 2414 19702 2466
rect 19764 2414 19776 2466
rect 19838 2414 19840 2466
rect 19678 2412 19702 2414
rect 19758 2412 19782 2414
rect 19838 2412 19862 2414
rect 19622 2392 19918 2412
rect 23492 2409 23520 4647
rect 23478 2400 23534 2409
rect 23478 2335 23534 2344
rect 5622 1924 5918 1944
rect 5678 1922 5702 1924
rect 5758 1922 5782 1924
rect 5838 1922 5862 1924
rect 5700 1870 5702 1922
rect 5764 1870 5776 1922
rect 5838 1870 5840 1922
rect 5678 1868 5702 1870
rect 5758 1868 5782 1870
rect 5838 1868 5862 1870
rect 5622 1848 5918 1868
rect 14956 1924 15252 1944
rect 15012 1922 15036 1924
rect 15092 1922 15116 1924
rect 15172 1922 15196 1924
rect 15034 1870 15036 1922
rect 15098 1870 15110 1922
rect 15172 1870 15174 1922
rect 15012 1868 15036 1870
rect 15092 1868 15116 1870
rect 15172 1868 15196 1870
rect 14956 1848 15252 1868
rect 23584 97 23612 12014
rect 23662 7704 23718 7713
rect 23662 7639 23718 7648
rect 23676 5401 23704 7639
rect 23662 5392 23718 5401
rect 23662 5327 23718 5336
rect 23662 4984 23718 4993
rect 23662 4919 23718 4928
rect 23676 641 23704 4919
rect 23768 2137 23796 15822
rect 23860 13250 23888 20174
rect 23952 20118 23980 20854
rect 23940 20112 23992 20118
rect 23940 20054 23992 20060
rect 24032 19636 24084 19642
rect 24032 19578 24084 19584
rect 24044 19234 24072 19578
rect 24124 19568 24176 19574
rect 24124 19510 24176 19516
rect 24032 19228 24084 19234
rect 24032 19170 24084 19176
rect 24044 18690 24072 19170
rect 24136 19166 24164 19510
rect 24124 19160 24176 19166
rect 24124 19102 24176 19108
rect 24032 18684 24084 18690
rect 24032 18626 24084 18632
rect 24136 18622 24164 19102
rect 24124 18616 24176 18622
rect 24124 18558 24176 18564
rect 24124 17868 24176 17874
rect 24124 17810 24176 17816
rect 24136 17466 24164 17810
rect 24124 17460 24176 17466
rect 24124 17402 24176 17408
rect 23940 16848 23992 16854
rect 23938 16816 23940 16825
rect 23992 16816 23994 16825
rect 23938 16751 23994 16760
rect 24030 16544 24086 16553
rect 24030 16479 24086 16488
rect 23940 16236 23992 16242
rect 23940 16178 23992 16184
rect 23952 13794 23980 16178
rect 24044 15426 24072 16479
rect 24124 16304 24176 16310
rect 24124 16246 24176 16252
rect 24032 15420 24084 15426
rect 24032 15362 24084 15368
rect 24136 15306 24164 16246
rect 24044 15278 24164 15306
rect 23940 13788 23992 13794
rect 23940 13730 23992 13736
rect 23848 13244 23900 13250
rect 23848 13186 23900 13192
rect 23938 13144 23994 13153
rect 23938 13079 23994 13088
rect 23952 10326 23980 13079
rect 24044 12162 24072 15278
rect 24124 15216 24176 15222
rect 24124 15158 24176 15164
rect 24136 14882 24164 15158
rect 24124 14876 24176 14882
rect 24124 14818 24176 14824
rect 24228 12706 24256 21092
rect 24676 20860 24728 20866
rect 24676 20802 24728 20808
rect 24289 20420 24585 20440
rect 24345 20418 24369 20420
rect 24425 20418 24449 20420
rect 24505 20418 24529 20420
rect 24367 20366 24369 20418
rect 24431 20366 24443 20418
rect 24505 20366 24507 20418
rect 24345 20364 24369 20366
rect 24425 20364 24449 20366
rect 24505 20364 24529 20366
rect 24289 20344 24585 20364
rect 24289 19332 24585 19352
rect 24345 19330 24369 19332
rect 24425 19330 24449 19332
rect 24505 19330 24529 19332
rect 24367 19278 24369 19330
rect 24431 19278 24443 19330
rect 24505 19278 24507 19330
rect 24345 19276 24369 19278
rect 24425 19276 24449 19278
rect 24505 19276 24529 19278
rect 24289 19256 24585 19276
rect 24289 18244 24585 18264
rect 24345 18242 24369 18244
rect 24425 18242 24449 18244
rect 24505 18242 24529 18244
rect 24367 18190 24369 18242
rect 24431 18190 24443 18242
rect 24505 18190 24507 18242
rect 24345 18188 24369 18190
rect 24425 18188 24449 18190
rect 24505 18188 24529 18190
rect 24289 18168 24585 18188
rect 24289 17156 24585 17176
rect 24345 17154 24369 17156
rect 24425 17154 24449 17156
rect 24505 17154 24529 17156
rect 24367 17102 24369 17154
rect 24431 17102 24443 17154
rect 24505 17102 24507 17154
rect 24345 17100 24369 17102
rect 24425 17100 24449 17102
rect 24505 17100 24529 17102
rect 24289 17080 24585 17100
rect 24289 16068 24585 16088
rect 24345 16066 24369 16068
rect 24425 16066 24449 16068
rect 24505 16066 24529 16068
rect 24367 16014 24369 16066
rect 24431 16014 24443 16066
rect 24505 16014 24507 16066
rect 24345 16012 24369 16014
rect 24425 16012 24449 16014
rect 24505 16012 24529 16014
rect 24289 15992 24585 16012
rect 24688 15850 24716 20802
rect 24872 20798 24900 22638
rect 24952 22152 25004 22158
rect 24950 22120 24952 22129
rect 25004 22120 25006 22129
rect 24950 22055 25006 22064
rect 25136 21200 25188 21206
rect 25134 21168 25136 21177
rect 25188 21168 25190 21177
rect 25134 21103 25190 21112
rect 24860 20792 24912 20798
rect 24860 20734 24912 20740
rect 24860 20656 24912 20662
rect 24860 20598 24912 20604
rect 24768 19772 24820 19778
rect 24768 19714 24820 19720
rect 24780 19234 24808 19714
rect 24872 19642 24900 20598
rect 25134 20352 25190 20361
rect 25134 20287 25136 20296
rect 25188 20287 25190 20296
rect 25136 20258 25188 20264
rect 24952 19976 25004 19982
rect 24952 19918 25004 19924
rect 24964 19681 24992 19918
rect 24950 19672 25006 19681
rect 24860 19636 24912 19642
rect 24950 19607 25006 19616
rect 24860 19578 24912 19584
rect 24768 19228 24820 19234
rect 24768 19170 24820 19176
rect 25134 19128 25190 19137
rect 25134 19063 25190 19072
rect 25148 18894 25176 19063
rect 25136 18888 25188 18894
rect 25136 18830 25188 18836
rect 25136 18480 25188 18486
rect 25136 18422 25188 18428
rect 25148 17942 25176 18422
rect 25136 17936 25188 17942
rect 24766 17904 24822 17913
rect 25136 17878 25188 17884
rect 24766 17839 24822 17848
rect 24780 17602 24808 17839
rect 25240 17754 25268 23794
rect 25516 23353 25544 27240
rect 26160 23858 26188 27240
rect 26148 23852 26200 23858
rect 26148 23794 26200 23800
rect 25502 23344 25558 23353
rect 25502 23279 25558 23288
rect 25410 23072 25466 23081
rect 25410 23007 25412 23016
rect 25464 23007 25466 23016
rect 25412 22978 25464 22984
rect 25688 22900 25740 22906
rect 25688 22842 25740 22848
rect 25700 22158 25728 22842
rect 25688 22152 25740 22158
rect 25688 22094 25740 22100
rect 25700 21857 25728 22094
rect 25686 21848 25742 21857
rect 25686 21783 25742 21792
rect 26240 21132 26292 21138
rect 26240 21074 26292 21080
rect 25320 21064 25372 21070
rect 25320 21006 25372 21012
rect 25332 20905 25360 21006
rect 25318 20896 25374 20905
rect 25318 20831 25374 20840
rect 25320 20724 25372 20730
rect 25320 20666 25372 20672
rect 25332 20322 25360 20666
rect 25504 20656 25556 20662
rect 25504 20598 25556 20604
rect 25320 20316 25372 20322
rect 25320 20258 25372 20264
rect 25412 19772 25464 19778
rect 25412 19714 25464 19720
rect 25424 19681 25452 19714
rect 25410 19672 25466 19681
rect 25410 19607 25466 19616
rect 25516 19030 25544 20598
rect 25594 20216 25650 20225
rect 25594 20151 25650 20160
rect 25504 19024 25556 19030
rect 25504 18966 25556 18972
rect 25318 18448 25374 18457
rect 25318 18383 25374 18392
rect 25332 18146 25360 18383
rect 25320 18140 25372 18146
rect 25320 18082 25372 18088
rect 25148 17726 25268 17754
rect 24768 17596 24820 17602
rect 24768 17538 24820 17544
rect 25044 17460 25096 17466
rect 25044 17402 25096 17408
rect 25056 17058 25084 17402
rect 25044 17052 25096 17058
rect 25044 16994 25096 17000
rect 24766 16136 24822 16145
rect 24766 16071 24822 16080
rect 24780 15970 24808 16071
rect 24768 15964 24820 15970
rect 24768 15906 24820 15912
rect 24688 15822 24808 15850
rect 24676 15760 24728 15766
rect 24676 15702 24728 15708
rect 24289 14980 24585 15000
rect 24345 14978 24369 14980
rect 24425 14978 24449 14980
rect 24505 14978 24529 14980
rect 24367 14926 24369 14978
rect 24431 14926 24443 14978
rect 24505 14926 24507 14978
rect 24345 14924 24369 14926
rect 24425 14924 24449 14926
rect 24505 14924 24529 14926
rect 24289 14904 24585 14924
rect 24688 14746 24716 15702
rect 24676 14740 24728 14746
rect 24676 14682 24728 14688
rect 24584 14672 24636 14678
rect 24584 14614 24636 14620
rect 24596 14338 24624 14614
rect 24584 14332 24636 14338
rect 24584 14274 24636 14280
rect 24289 13892 24585 13912
rect 24345 13890 24369 13892
rect 24425 13890 24449 13892
rect 24505 13890 24529 13892
rect 24367 13838 24369 13890
rect 24431 13838 24443 13890
rect 24505 13838 24507 13890
rect 24345 13836 24369 13838
rect 24425 13836 24449 13838
rect 24505 13836 24529 13838
rect 24289 13816 24585 13836
rect 24289 12804 24585 12824
rect 24345 12802 24369 12804
rect 24425 12802 24449 12804
rect 24505 12802 24529 12804
rect 24367 12750 24369 12802
rect 24431 12750 24443 12802
rect 24505 12750 24507 12802
rect 24345 12748 24369 12750
rect 24425 12748 24449 12750
rect 24505 12748 24529 12750
rect 24289 12728 24585 12748
rect 24216 12700 24268 12706
rect 24216 12642 24268 12648
rect 24674 12600 24730 12609
rect 24674 12535 24676 12544
rect 24728 12535 24730 12544
rect 24676 12506 24728 12512
rect 24032 12156 24084 12162
rect 24032 12098 24084 12104
rect 24584 12020 24636 12026
rect 24584 11962 24636 11968
rect 24596 11929 24624 11962
rect 24582 11920 24638 11929
rect 24638 11878 24716 11906
rect 24582 11855 24638 11864
rect 24289 11716 24585 11736
rect 24345 11714 24369 11716
rect 24425 11714 24449 11716
rect 24505 11714 24529 11716
rect 24367 11662 24369 11714
rect 24431 11662 24443 11714
rect 24505 11662 24507 11714
rect 24345 11660 24369 11662
rect 24425 11660 24449 11662
rect 24505 11660 24529 11662
rect 24289 11640 24585 11660
rect 24688 11618 24716 11878
rect 24676 11612 24728 11618
rect 24676 11554 24728 11560
rect 24780 11074 24808 15822
rect 24860 15420 24912 15426
rect 24860 15362 24912 15368
rect 24872 14882 24900 15362
rect 24860 14876 24912 14882
rect 24860 14818 24912 14824
rect 25044 14536 25096 14542
rect 25044 14478 25096 14484
rect 25056 14270 25084 14478
rect 25148 14338 25176 17726
rect 25410 17360 25466 17369
rect 25410 17295 25466 17304
rect 25424 17058 25452 17295
rect 25412 17052 25464 17058
rect 25412 16994 25464 17000
rect 25410 16680 25466 16689
rect 25410 16615 25466 16624
rect 25424 16514 25452 16615
rect 25412 16508 25464 16514
rect 25412 16450 25464 16456
rect 25228 16372 25280 16378
rect 25228 16314 25280 16320
rect 25240 15970 25268 16314
rect 25228 15964 25280 15970
rect 25228 15906 25280 15912
rect 25502 15456 25558 15465
rect 25608 15426 25636 20151
rect 25872 19636 25924 19642
rect 25872 19578 25924 19584
rect 25884 19234 25912 19578
rect 25872 19228 25924 19234
rect 25872 19170 25924 19176
rect 25502 15391 25558 15400
rect 25596 15420 25648 15426
rect 25516 14882 25544 15391
rect 25596 15362 25648 15368
rect 25872 15284 25924 15290
rect 25872 15226 25924 15232
rect 25884 14921 25912 15226
rect 25870 14912 25926 14921
rect 25504 14876 25556 14882
rect 25870 14847 25872 14856
rect 25504 14818 25556 14824
rect 25924 14847 25926 14856
rect 25872 14818 25924 14824
rect 25884 14787 25912 14818
rect 25594 14368 25650 14377
rect 25136 14332 25188 14338
rect 25594 14303 25650 14312
rect 25136 14274 25188 14280
rect 25044 14264 25096 14270
rect 25044 14206 25096 14212
rect 25608 14202 25636 14303
rect 25596 14196 25648 14202
rect 25596 14138 25648 14144
rect 25608 13794 25636 14138
rect 25596 13788 25648 13794
rect 25596 13730 25648 13736
rect 25226 13688 25282 13697
rect 25226 13623 25228 13632
rect 25280 13623 25282 13632
rect 25228 13594 25280 13600
rect 25042 13144 25098 13153
rect 25042 13079 25044 13088
rect 25096 13079 25098 13088
rect 25044 13050 25096 13056
rect 25056 12706 25084 13050
rect 25044 12700 25096 12706
rect 25044 12642 25096 12648
rect 24768 11068 24820 11074
rect 24768 11010 24820 11016
rect 24676 10932 24728 10938
rect 24676 10874 24728 10880
rect 24688 10705 24716 10874
rect 24030 10696 24086 10705
rect 24674 10696 24730 10705
rect 24030 10631 24086 10640
rect 23940 10320 23992 10326
rect 23940 10262 23992 10268
rect 24044 3225 24072 10631
rect 24289 10628 24585 10648
rect 24674 10631 24730 10640
rect 24345 10626 24369 10628
rect 24425 10626 24449 10628
rect 24505 10626 24529 10628
rect 24367 10574 24369 10626
rect 24431 10574 24443 10626
rect 24505 10574 24507 10626
rect 24345 10572 24369 10574
rect 24425 10572 24449 10574
rect 24505 10572 24529 10574
rect 24122 10560 24178 10569
rect 24289 10552 24585 10572
rect 24688 10530 24716 10631
rect 24122 10495 24178 10504
rect 24676 10524 24728 10530
rect 24136 10462 24164 10495
rect 24676 10466 24728 10472
rect 24124 10456 24176 10462
rect 24124 10398 24176 10404
rect 24124 10320 24176 10326
rect 24124 10262 24176 10268
rect 24030 3216 24086 3225
rect 24030 3151 24086 3160
rect 23754 2128 23810 2137
rect 23754 2063 23810 2072
rect 24136 1185 24164 10262
rect 25228 10184 25280 10190
rect 25226 10152 25228 10161
rect 25280 10152 25282 10161
rect 25226 10087 25282 10096
rect 24676 9844 24728 9850
rect 24676 9786 24728 9792
rect 24688 9617 24716 9786
rect 24674 9608 24730 9617
rect 24289 9540 24585 9560
rect 24674 9543 24730 9552
rect 25226 9608 25282 9617
rect 25226 9543 25282 9552
rect 24345 9538 24369 9540
rect 24425 9538 24449 9540
rect 24505 9538 24529 9540
rect 24367 9486 24369 9538
rect 24431 9486 24443 9538
rect 24505 9486 24507 9538
rect 24345 9484 24369 9486
rect 24425 9484 24449 9486
rect 24505 9484 24529 9486
rect 24289 9464 24585 9484
rect 25240 9374 25268 9543
rect 24768 9368 24820 9374
rect 24766 9336 24768 9345
rect 25228 9368 25280 9374
rect 24820 9336 24822 9345
rect 25228 9310 25280 9316
rect 24766 9271 24822 9280
rect 24492 9096 24544 9102
rect 24492 9038 24544 9044
rect 24766 9064 24822 9073
rect 24504 8937 24532 9038
rect 24766 8999 24822 9008
rect 24490 8928 24546 8937
rect 24780 8898 24808 8999
rect 24490 8863 24546 8872
rect 24768 8892 24820 8898
rect 24768 8834 24820 8840
rect 24676 8756 24728 8762
rect 24676 8698 24728 8704
rect 24289 8452 24585 8472
rect 24345 8450 24369 8452
rect 24425 8450 24449 8452
rect 24505 8450 24529 8452
rect 24367 8398 24369 8450
rect 24431 8398 24443 8450
rect 24505 8398 24507 8450
rect 24345 8396 24369 8398
rect 24425 8396 24449 8398
rect 24505 8396 24529 8398
rect 24289 8376 24585 8396
rect 24688 8393 24716 8698
rect 24674 8384 24730 8393
rect 24674 8319 24676 8328
rect 24728 8319 24730 8328
rect 24676 8290 24728 8296
rect 24582 7704 24638 7713
rect 24582 7639 24584 7648
rect 24636 7639 24638 7648
rect 24584 7610 24636 7616
rect 24596 7554 24624 7610
rect 24766 7568 24822 7577
rect 24596 7526 24716 7554
rect 24289 7364 24585 7384
rect 24345 7362 24369 7364
rect 24425 7362 24449 7364
rect 24505 7362 24529 7364
rect 24367 7310 24369 7362
rect 24431 7310 24443 7362
rect 24505 7310 24507 7362
rect 24345 7308 24369 7310
rect 24425 7308 24449 7310
rect 24505 7308 24529 7310
rect 24289 7288 24585 7308
rect 24688 7266 24716 7526
rect 24766 7503 24768 7512
rect 24820 7503 24822 7512
rect 24768 7474 24820 7480
rect 24676 7260 24728 7266
rect 24676 7202 24728 7208
rect 24289 6276 24585 6296
rect 24345 6274 24369 6276
rect 24425 6274 24449 6276
rect 24505 6274 24529 6276
rect 24367 6222 24369 6274
rect 24431 6222 24443 6274
rect 24505 6222 24507 6274
rect 24345 6220 24369 6222
rect 24425 6220 24449 6222
rect 24505 6220 24529 6222
rect 24289 6200 24585 6220
rect 24674 6072 24730 6081
rect 24674 6007 24730 6016
rect 24289 5188 24585 5208
rect 24345 5186 24369 5188
rect 24425 5186 24449 5188
rect 24505 5186 24529 5188
rect 24367 5134 24369 5186
rect 24431 5134 24443 5186
rect 24505 5134 24507 5186
rect 24345 5132 24369 5134
rect 24425 5132 24449 5134
rect 24505 5132 24529 5134
rect 24289 5112 24585 5132
rect 24688 4177 24716 6007
rect 24674 4168 24730 4177
rect 24289 4100 24585 4120
rect 24674 4103 24730 4112
rect 24345 4098 24369 4100
rect 24425 4098 24449 4100
rect 24505 4098 24529 4100
rect 24367 4046 24369 4098
rect 24431 4046 24443 4098
rect 24505 4046 24507 4098
rect 24345 4044 24369 4046
rect 24425 4044 24449 4046
rect 24505 4044 24529 4046
rect 24289 4024 24585 4044
rect 26252 3769 26280 21074
rect 26896 20225 26924 27240
rect 27540 21138 27568 27240
rect 27528 21132 27580 21138
rect 27528 21074 27580 21080
rect 26882 20216 26938 20225
rect 26882 20151 26938 20160
rect 24766 3760 24822 3769
rect 24766 3695 24822 3704
rect 26238 3760 26294 3769
rect 26238 3695 26294 3704
rect 24780 3662 24808 3695
rect 24768 3656 24820 3662
rect 25228 3656 25280 3662
rect 24768 3598 24820 3604
rect 25226 3624 25228 3633
rect 25280 3624 25282 3633
rect 25226 3559 25282 3568
rect 24289 3012 24585 3032
rect 24345 3010 24369 3012
rect 24425 3010 24449 3012
rect 24505 3010 24529 3012
rect 24367 2958 24369 3010
rect 24431 2958 24443 3010
rect 24505 2958 24507 3010
rect 24345 2956 24369 2958
rect 24425 2956 24449 2958
rect 24505 2956 24529 2958
rect 24289 2936 24585 2956
rect 24289 1924 24585 1944
rect 24345 1922 24369 1924
rect 24425 1922 24449 1924
rect 24505 1922 24529 1924
rect 24367 1870 24369 1922
rect 24431 1870 24443 1922
rect 24505 1870 24507 1922
rect 24345 1868 24369 1870
rect 24425 1868 24449 1870
rect 24505 1868 24529 1870
rect 24289 1848 24585 1868
rect 24122 1176 24178 1185
rect 24122 1111 24178 1120
rect 23662 632 23718 641
rect 23662 567 23718 576
rect 23570 88 23626 97
rect 23570 23 23626 32
<< via2 >>
rect 23202 27368 23258 27424
rect 938 17304 994 17360
rect 3422 22744 3478 22800
rect 3422 20704 3478 20760
rect 4342 23288 4398 23344
rect 5622 24770 5678 24772
rect 5702 24770 5758 24772
rect 5782 24770 5838 24772
rect 5862 24770 5918 24772
rect 5622 24718 5648 24770
rect 5648 24718 5678 24770
rect 5702 24718 5712 24770
rect 5712 24718 5758 24770
rect 5782 24718 5828 24770
rect 5828 24718 5838 24770
rect 5862 24718 5892 24770
rect 5892 24718 5918 24770
rect 5622 24716 5678 24718
rect 5702 24716 5758 24718
rect 5782 24716 5838 24718
rect 5862 24716 5918 24718
rect 5622 23682 5678 23684
rect 5702 23682 5758 23684
rect 5782 23682 5838 23684
rect 5862 23682 5918 23684
rect 5622 23630 5648 23682
rect 5648 23630 5678 23682
rect 5702 23630 5712 23682
rect 5712 23630 5758 23682
rect 5782 23630 5828 23682
rect 5828 23630 5838 23682
rect 5862 23630 5892 23682
rect 5892 23630 5918 23682
rect 5622 23628 5678 23630
rect 5702 23628 5758 23630
rect 5782 23628 5838 23630
rect 5862 23628 5918 23630
rect 5622 22594 5678 22596
rect 5702 22594 5758 22596
rect 5782 22594 5838 22596
rect 5862 22594 5918 22596
rect 5622 22542 5648 22594
rect 5648 22542 5678 22594
rect 5702 22542 5712 22594
rect 5712 22542 5758 22594
rect 5782 22542 5828 22594
rect 5828 22542 5838 22594
rect 5862 22542 5892 22594
rect 5892 22542 5918 22594
rect 5622 22540 5678 22542
rect 5702 22540 5758 22542
rect 5782 22540 5838 22542
rect 5862 22540 5918 22542
rect 4986 22200 5042 22256
rect 5622 21506 5678 21508
rect 5702 21506 5758 21508
rect 5782 21506 5838 21508
rect 5862 21506 5918 21508
rect 5622 21454 5648 21506
rect 5648 21454 5678 21506
rect 5702 21454 5712 21506
rect 5712 21454 5758 21506
rect 5782 21454 5828 21506
rect 5828 21454 5838 21506
rect 5862 21454 5892 21506
rect 5892 21454 5918 21506
rect 5622 21452 5678 21454
rect 5702 21452 5758 21454
rect 5782 21452 5838 21454
rect 5862 21452 5918 21454
rect 6366 21520 6422 21576
rect 7746 22336 7802 22392
rect 7102 21384 7158 21440
rect 5998 20704 6054 20760
rect 5622 20418 5678 20420
rect 5702 20418 5758 20420
rect 5782 20418 5838 20420
rect 5862 20418 5918 20420
rect 5622 20366 5648 20418
rect 5648 20366 5678 20418
rect 5702 20366 5712 20418
rect 5712 20366 5758 20418
rect 5782 20366 5828 20418
rect 5828 20366 5838 20418
rect 5862 20366 5892 20418
rect 5892 20366 5918 20418
rect 5622 20364 5678 20366
rect 5702 20364 5758 20366
rect 5782 20364 5838 20366
rect 5862 20364 5918 20366
rect 5622 19330 5678 19332
rect 5702 19330 5758 19332
rect 5782 19330 5838 19332
rect 5862 19330 5918 19332
rect 5622 19278 5648 19330
rect 5648 19278 5678 19330
rect 5702 19278 5712 19330
rect 5712 19278 5758 19330
rect 5782 19278 5828 19330
rect 5828 19278 5838 19330
rect 5862 19278 5892 19330
rect 5892 19278 5918 19330
rect 5622 19276 5678 19278
rect 5702 19276 5758 19278
rect 5782 19276 5838 19278
rect 5862 19276 5918 19278
rect 3698 19072 3754 19128
rect 10289 25314 10345 25316
rect 10369 25314 10425 25316
rect 10449 25314 10505 25316
rect 10529 25314 10585 25316
rect 10289 25262 10315 25314
rect 10315 25262 10345 25314
rect 10369 25262 10379 25314
rect 10379 25262 10425 25314
rect 10449 25262 10495 25314
rect 10495 25262 10505 25314
rect 10529 25262 10559 25314
rect 10559 25262 10585 25314
rect 10289 25260 10345 25262
rect 10369 25260 10425 25262
rect 10449 25260 10505 25262
rect 10529 25260 10585 25262
rect 10289 24226 10345 24228
rect 10369 24226 10425 24228
rect 10449 24226 10505 24228
rect 10529 24226 10585 24228
rect 10289 24174 10315 24226
rect 10315 24174 10345 24226
rect 10369 24174 10379 24226
rect 10379 24174 10425 24226
rect 10449 24174 10495 24226
rect 10495 24174 10505 24226
rect 10529 24174 10559 24226
rect 10559 24174 10585 24226
rect 10289 24172 10345 24174
rect 10369 24172 10425 24174
rect 10449 24172 10505 24174
rect 10529 24172 10585 24174
rect 10690 24104 10746 24160
rect 9770 23968 9826 24024
rect 10289 23138 10345 23140
rect 10369 23138 10425 23140
rect 10449 23138 10505 23140
rect 10529 23138 10585 23140
rect 10289 23086 10315 23138
rect 10315 23086 10345 23138
rect 10369 23086 10379 23138
rect 10379 23086 10425 23138
rect 10449 23086 10495 23138
rect 10495 23086 10505 23138
rect 10529 23086 10559 23138
rect 10559 23086 10585 23138
rect 10289 23084 10345 23086
rect 10369 23084 10425 23086
rect 10449 23084 10505 23086
rect 10529 23084 10585 23086
rect 11150 23560 11206 23616
rect 11242 22744 11298 22800
rect 13174 24512 13230 24568
rect 12530 24376 12586 24432
rect 12162 23016 12218 23072
rect 13450 23580 13506 23616
rect 13450 23560 13452 23580
rect 13452 23560 13504 23580
rect 13504 23560 13506 23580
rect 12714 22744 12770 22800
rect 13726 22780 13728 22800
rect 13728 22780 13780 22800
rect 13780 22780 13782 22800
rect 13726 22744 13782 22780
rect 10289 22050 10345 22052
rect 10369 22050 10425 22052
rect 10449 22050 10505 22052
rect 10529 22050 10585 22052
rect 10289 21998 10315 22050
rect 10315 21998 10345 22050
rect 10369 21998 10379 22050
rect 10379 21998 10425 22050
rect 10449 21998 10495 22050
rect 10495 21998 10505 22050
rect 10529 21998 10559 22050
rect 10559 21998 10585 22050
rect 10289 21996 10345 21998
rect 10369 21996 10425 21998
rect 10449 21996 10505 21998
rect 10529 21996 10585 21998
rect 11518 21520 11574 21576
rect 9126 21112 9182 21168
rect 13726 22064 13782 22120
rect 10289 20962 10345 20964
rect 10369 20962 10425 20964
rect 10449 20962 10505 20964
rect 10529 20962 10585 20964
rect 10289 20910 10315 20962
rect 10315 20910 10345 20962
rect 10369 20910 10379 20962
rect 10379 20910 10425 20962
rect 10449 20910 10495 20962
rect 10495 20910 10505 20962
rect 10529 20910 10559 20962
rect 10559 20910 10585 20962
rect 10289 20908 10345 20910
rect 10369 20908 10425 20910
rect 10449 20908 10505 20910
rect 10529 20908 10585 20910
rect 10874 20044 10930 20080
rect 10874 20024 10876 20044
rect 10876 20024 10928 20044
rect 10928 20024 10930 20044
rect 10289 19874 10345 19876
rect 10369 19874 10425 19876
rect 10449 19874 10505 19876
rect 10529 19874 10585 19876
rect 10289 19822 10315 19874
rect 10315 19822 10345 19874
rect 10369 19822 10379 19874
rect 10379 19822 10425 19874
rect 10449 19822 10495 19874
rect 10495 19822 10505 19874
rect 10529 19822 10559 19874
rect 10559 19822 10585 19874
rect 10289 19820 10345 19822
rect 10369 19820 10425 19822
rect 10449 19820 10505 19822
rect 10529 19820 10585 19822
rect 8390 18936 8446 18992
rect 10289 18786 10345 18788
rect 10369 18786 10425 18788
rect 10449 18786 10505 18788
rect 10529 18786 10585 18788
rect 10289 18734 10315 18786
rect 10315 18734 10345 18786
rect 10369 18734 10379 18786
rect 10379 18734 10425 18786
rect 10449 18734 10495 18786
rect 10495 18734 10505 18786
rect 10529 18734 10559 18786
rect 10559 18734 10585 18786
rect 10289 18732 10345 18734
rect 10369 18732 10425 18734
rect 10449 18732 10505 18734
rect 10529 18732 10585 18734
rect 2962 18392 3018 18448
rect 5622 18242 5678 18244
rect 5702 18242 5758 18244
rect 5782 18242 5838 18244
rect 5862 18242 5918 18244
rect 5622 18190 5648 18242
rect 5648 18190 5678 18242
rect 5702 18190 5712 18242
rect 5712 18190 5758 18242
rect 5782 18190 5828 18242
rect 5828 18190 5838 18242
rect 5862 18190 5892 18242
rect 5892 18190 5918 18242
rect 5622 18188 5678 18190
rect 5702 18188 5758 18190
rect 5782 18188 5838 18190
rect 5862 18188 5918 18190
rect 2318 17848 2374 17904
rect 10289 17698 10345 17700
rect 10369 17698 10425 17700
rect 10449 17698 10505 17700
rect 10529 17698 10585 17700
rect 10289 17646 10315 17698
rect 10315 17646 10345 17698
rect 10369 17646 10379 17698
rect 10379 17646 10425 17698
rect 10449 17646 10495 17698
rect 10495 17646 10505 17698
rect 10529 17646 10559 17698
rect 10559 17646 10585 17698
rect 10289 17644 10345 17646
rect 10369 17644 10425 17646
rect 10449 17644 10505 17646
rect 10529 17644 10585 17646
rect 5622 17154 5678 17156
rect 5702 17154 5758 17156
rect 5782 17154 5838 17156
rect 5862 17154 5918 17156
rect 5622 17102 5648 17154
rect 5648 17102 5678 17154
rect 5702 17102 5712 17154
rect 5712 17102 5758 17154
rect 5782 17102 5828 17154
rect 5828 17102 5838 17154
rect 5862 17102 5892 17154
rect 5892 17102 5918 17154
rect 5622 17100 5678 17102
rect 5702 17100 5758 17102
rect 5782 17100 5838 17102
rect 5862 17100 5918 17102
rect 13542 21132 13598 21168
rect 13542 21112 13544 21132
rect 13544 21112 13596 21132
rect 13596 21112 13598 21132
rect 13542 20432 13598 20488
rect 13450 18956 13506 18992
rect 13450 18936 13452 18956
rect 13452 18936 13504 18956
rect 13504 18936 13506 18956
rect 11794 16896 11850 16952
rect 1582 16760 1638 16816
rect 10289 16610 10345 16612
rect 10369 16610 10425 16612
rect 10449 16610 10505 16612
rect 10529 16610 10585 16612
rect 10289 16558 10315 16610
rect 10315 16558 10345 16610
rect 10369 16558 10379 16610
rect 10379 16558 10425 16610
rect 10449 16558 10495 16610
rect 10495 16558 10505 16610
rect 10529 16558 10559 16610
rect 10559 16558 10585 16610
rect 10289 16556 10345 16558
rect 10369 16556 10425 16558
rect 10449 16556 10505 16558
rect 10529 16556 10585 16558
rect 5622 16066 5678 16068
rect 5702 16066 5758 16068
rect 5782 16066 5838 16068
rect 5862 16066 5918 16068
rect 5622 16014 5648 16066
rect 5648 16014 5678 16066
rect 5702 16014 5712 16066
rect 5712 16014 5758 16066
rect 5782 16014 5828 16066
rect 5828 16014 5838 16066
rect 5862 16014 5892 16066
rect 5892 16014 5918 16066
rect 5622 16012 5678 16014
rect 5702 16012 5758 16014
rect 5782 16012 5838 16014
rect 5862 16012 5918 16014
rect 10289 15522 10345 15524
rect 10369 15522 10425 15524
rect 10449 15522 10505 15524
rect 10529 15522 10585 15524
rect 10289 15470 10315 15522
rect 10315 15470 10345 15522
rect 10369 15470 10379 15522
rect 10379 15470 10425 15522
rect 10449 15470 10495 15522
rect 10495 15470 10505 15522
rect 10529 15470 10559 15522
rect 10559 15470 10585 15522
rect 10289 15468 10345 15470
rect 10369 15468 10425 15470
rect 10449 15468 10505 15470
rect 10529 15468 10585 15470
rect 5622 14978 5678 14980
rect 5702 14978 5758 14980
rect 5782 14978 5838 14980
rect 5862 14978 5918 14980
rect 5622 14926 5648 14978
rect 5648 14926 5678 14978
rect 5702 14926 5712 14978
rect 5712 14926 5758 14978
rect 5782 14926 5828 14978
rect 5828 14926 5838 14978
rect 5862 14926 5892 14978
rect 5892 14926 5918 14978
rect 5622 14924 5678 14926
rect 5702 14924 5758 14926
rect 5782 14924 5838 14926
rect 5862 14924 5918 14926
rect 10289 14434 10345 14436
rect 10369 14434 10425 14436
rect 10449 14434 10505 14436
rect 10529 14434 10585 14436
rect 10289 14382 10315 14434
rect 10315 14382 10345 14434
rect 10369 14382 10379 14434
rect 10379 14382 10425 14434
rect 10449 14382 10495 14434
rect 10495 14382 10505 14434
rect 10529 14382 10559 14434
rect 10559 14382 10585 14434
rect 10289 14380 10345 14382
rect 10369 14380 10425 14382
rect 10449 14380 10505 14382
rect 10529 14380 10585 14382
rect 13634 18836 13636 18856
rect 13636 18836 13688 18856
rect 13688 18836 13690 18856
rect 13634 18800 13690 18836
rect 14002 22064 14058 22120
rect 14278 21676 14334 21712
rect 14278 21656 14280 21676
rect 14280 21656 14332 21676
rect 14332 21656 14334 21676
rect 14956 24770 15012 24772
rect 15036 24770 15092 24772
rect 15116 24770 15172 24772
rect 15196 24770 15252 24772
rect 14956 24718 14982 24770
rect 14982 24718 15012 24770
rect 15036 24718 15046 24770
rect 15046 24718 15092 24770
rect 15116 24718 15162 24770
rect 15162 24718 15172 24770
rect 15196 24718 15226 24770
rect 15226 24718 15252 24770
rect 14956 24716 15012 24718
rect 15036 24716 15092 24718
rect 15116 24716 15172 24718
rect 15196 24716 15252 24718
rect 16118 23968 16174 24024
rect 15106 23832 15162 23888
rect 14956 23682 15012 23684
rect 15036 23682 15092 23684
rect 15116 23682 15172 23684
rect 15196 23682 15252 23684
rect 14956 23630 14982 23682
rect 14982 23630 15012 23682
rect 15036 23630 15046 23682
rect 15046 23630 15092 23682
rect 15116 23630 15162 23682
rect 15162 23630 15172 23682
rect 15196 23630 15226 23682
rect 15226 23630 15252 23682
rect 14956 23628 15012 23630
rect 15036 23628 15092 23630
rect 15116 23628 15172 23630
rect 15196 23628 15252 23630
rect 14830 23016 14886 23072
rect 15198 23036 15254 23072
rect 15198 23016 15200 23036
rect 15200 23016 15252 23036
rect 15252 23016 15254 23036
rect 14956 22594 15012 22596
rect 15036 22594 15092 22596
rect 15116 22594 15172 22596
rect 15196 22594 15252 22596
rect 14956 22542 14982 22594
rect 14982 22542 15012 22594
rect 15036 22542 15046 22594
rect 15046 22542 15092 22594
rect 15116 22542 15162 22594
rect 15162 22542 15172 22594
rect 15196 22542 15226 22594
rect 15226 22542 15252 22594
rect 14956 22540 15012 22542
rect 15036 22540 15092 22542
rect 15116 22540 15172 22542
rect 15196 22540 15252 22542
rect 14956 21506 15012 21508
rect 15036 21506 15092 21508
rect 15116 21506 15172 21508
rect 15196 21506 15252 21508
rect 14956 21454 14982 21506
rect 14982 21454 15012 21506
rect 15036 21454 15046 21506
rect 15046 21454 15092 21506
rect 15116 21454 15162 21506
rect 15162 21454 15172 21506
rect 15196 21454 15226 21506
rect 15226 21454 15252 21506
rect 14956 21452 15012 21454
rect 15036 21452 15092 21454
rect 15116 21452 15172 21454
rect 15196 21452 15252 21454
rect 14646 20860 14702 20896
rect 14646 20840 14648 20860
rect 14648 20840 14700 20860
rect 14700 20840 14702 20860
rect 14554 20432 14610 20488
rect 14956 20418 15012 20420
rect 15036 20418 15092 20420
rect 15116 20418 15172 20420
rect 15196 20418 15252 20420
rect 14956 20366 14982 20418
rect 14982 20366 15012 20418
rect 15036 20366 15046 20418
rect 15046 20366 15092 20418
rect 15116 20366 15162 20418
rect 15162 20366 15172 20418
rect 15196 20366 15226 20418
rect 15226 20366 15252 20418
rect 14956 20364 15012 20366
rect 15036 20364 15092 20366
rect 15116 20364 15172 20366
rect 15196 20364 15252 20366
rect 14956 19330 15012 19332
rect 15036 19330 15092 19332
rect 15116 19330 15172 19332
rect 15196 19330 15252 19332
rect 14956 19278 14982 19330
rect 14982 19278 15012 19330
rect 15036 19278 15046 19330
rect 15046 19278 15092 19330
rect 15116 19278 15162 19330
rect 15162 19278 15172 19330
rect 15196 19278 15226 19330
rect 15226 19278 15252 19330
rect 14956 19276 15012 19278
rect 15036 19276 15092 19278
rect 15116 19276 15172 19278
rect 15196 19276 15252 19278
rect 14186 16796 14188 16816
rect 14188 16796 14240 16816
rect 14240 16796 14242 16816
rect 14186 16760 14242 16796
rect 14956 18242 15012 18244
rect 15036 18242 15092 18244
rect 15116 18242 15172 18244
rect 15196 18242 15252 18244
rect 14956 18190 14982 18242
rect 14982 18190 15012 18242
rect 15036 18190 15046 18242
rect 15046 18190 15092 18242
rect 15116 18190 15162 18242
rect 15162 18190 15172 18242
rect 15196 18190 15226 18242
rect 15226 18190 15252 18242
rect 14956 18188 15012 18190
rect 15036 18188 15092 18190
rect 15116 18188 15172 18190
rect 15196 18188 15252 18190
rect 15382 18140 15438 18176
rect 15382 18120 15384 18140
rect 15384 18120 15436 18140
rect 15436 18120 15438 18140
rect 14956 17154 15012 17156
rect 15036 17154 15092 17156
rect 15116 17154 15172 17156
rect 15196 17154 15252 17156
rect 14956 17102 14982 17154
rect 14982 17102 15012 17154
rect 15036 17102 15046 17154
rect 15046 17102 15092 17154
rect 15116 17102 15162 17154
rect 15162 17102 15172 17154
rect 15196 17102 15226 17154
rect 15226 17102 15252 17154
rect 14956 17100 15012 17102
rect 15036 17100 15092 17102
rect 15116 17100 15172 17102
rect 15196 17100 15252 17102
rect 13910 15400 13966 15456
rect 13910 15284 13966 15320
rect 13910 15264 13912 15284
rect 13912 15264 13964 15284
rect 13964 15264 13966 15284
rect 14956 16066 15012 16068
rect 15036 16066 15092 16068
rect 15116 16066 15172 16068
rect 15196 16066 15252 16068
rect 14956 16014 14982 16066
rect 14982 16014 15012 16066
rect 15036 16014 15046 16066
rect 15046 16014 15092 16066
rect 15116 16014 15162 16066
rect 15162 16014 15172 16066
rect 15196 16014 15226 16066
rect 15226 16014 15252 16066
rect 14956 16012 15012 16014
rect 15036 16012 15092 16014
rect 15116 16012 15172 16014
rect 15196 16012 15252 16014
rect 14956 14978 15012 14980
rect 15036 14978 15092 14980
rect 15116 14978 15172 14980
rect 15196 14978 15252 14980
rect 14956 14926 14982 14978
rect 14982 14926 15012 14978
rect 15036 14926 15046 14978
rect 15046 14926 15092 14978
rect 15116 14926 15162 14978
rect 15162 14926 15172 14978
rect 15196 14926 15226 14978
rect 15226 14926 15252 14978
rect 14956 14924 15012 14926
rect 15036 14924 15092 14926
rect 15116 14924 15172 14926
rect 15196 14924 15252 14926
rect 15842 21012 15844 21032
rect 15844 21012 15896 21032
rect 15896 21012 15898 21032
rect 15842 20976 15898 21012
rect 15566 20568 15622 20624
rect 15750 18836 15752 18856
rect 15752 18836 15804 18856
rect 15804 18836 15806 18856
rect 15750 18800 15806 18836
rect 15658 15572 15660 15592
rect 15660 15572 15712 15592
rect 15712 15572 15714 15592
rect 15658 15536 15714 15572
rect 5622 13890 5678 13892
rect 5702 13890 5758 13892
rect 5782 13890 5838 13892
rect 5862 13890 5918 13892
rect 5622 13838 5648 13890
rect 5648 13838 5678 13890
rect 5702 13838 5712 13890
rect 5712 13838 5758 13890
rect 5782 13838 5828 13890
rect 5828 13838 5838 13890
rect 5862 13838 5892 13890
rect 5892 13838 5918 13890
rect 5622 13836 5678 13838
rect 5702 13836 5758 13838
rect 5782 13836 5838 13838
rect 5862 13836 5918 13838
rect 10289 13346 10345 13348
rect 10369 13346 10425 13348
rect 10449 13346 10505 13348
rect 10529 13346 10585 13348
rect 10289 13294 10315 13346
rect 10315 13294 10345 13346
rect 10369 13294 10379 13346
rect 10379 13294 10425 13346
rect 10449 13294 10495 13346
rect 10495 13294 10505 13346
rect 10529 13294 10559 13346
rect 10559 13294 10585 13346
rect 10289 13292 10345 13294
rect 10369 13292 10425 13294
rect 10449 13292 10505 13294
rect 10529 13292 10585 13294
rect 5622 12802 5678 12804
rect 5702 12802 5758 12804
rect 5782 12802 5838 12804
rect 5862 12802 5918 12804
rect 5622 12750 5648 12802
rect 5648 12750 5678 12802
rect 5702 12750 5712 12802
rect 5712 12750 5758 12802
rect 5782 12750 5828 12802
rect 5828 12750 5838 12802
rect 5862 12750 5892 12802
rect 5892 12750 5918 12802
rect 5622 12748 5678 12750
rect 5702 12748 5758 12750
rect 5782 12748 5838 12750
rect 5862 12748 5918 12750
rect 10289 12258 10345 12260
rect 10369 12258 10425 12260
rect 10449 12258 10505 12260
rect 10529 12258 10585 12260
rect 10289 12206 10315 12258
rect 10315 12206 10345 12258
rect 10369 12206 10379 12258
rect 10379 12206 10425 12258
rect 10449 12206 10495 12258
rect 10495 12206 10505 12258
rect 10529 12206 10559 12258
rect 10559 12206 10585 12258
rect 10289 12204 10345 12206
rect 10369 12204 10425 12206
rect 10449 12204 10505 12206
rect 10529 12204 10585 12206
rect 5622 11714 5678 11716
rect 5702 11714 5758 11716
rect 5782 11714 5838 11716
rect 5862 11714 5918 11716
rect 5622 11662 5648 11714
rect 5648 11662 5678 11714
rect 5702 11662 5712 11714
rect 5712 11662 5758 11714
rect 5782 11662 5828 11714
rect 5828 11662 5838 11714
rect 5862 11662 5892 11714
rect 5892 11662 5918 11714
rect 5622 11660 5678 11662
rect 5702 11660 5758 11662
rect 5782 11660 5838 11662
rect 5862 11660 5918 11662
rect 3422 11320 3478 11376
rect 478 10912 534 10968
rect 10138 11340 10194 11376
rect 10138 11320 10140 11340
rect 10140 11320 10192 11340
rect 10192 11320 10194 11340
rect 10289 11170 10345 11172
rect 10369 11170 10425 11172
rect 10449 11170 10505 11172
rect 10529 11170 10585 11172
rect 10289 11118 10315 11170
rect 10315 11118 10345 11170
rect 10369 11118 10379 11170
rect 10379 11118 10425 11170
rect 10449 11118 10495 11170
rect 10495 11118 10505 11170
rect 10529 11118 10559 11170
rect 10559 11118 10585 11170
rect 10289 11116 10345 11118
rect 10369 11116 10425 11118
rect 10449 11116 10505 11118
rect 10529 11116 10585 11118
rect 15934 14720 15990 14776
rect 14956 13890 15012 13892
rect 15036 13890 15092 13892
rect 15116 13890 15172 13892
rect 15196 13890 15252 13892
rect 14956 13838 14982 13890
rect 14982 13838 15012 13890
rect 15036 13838 15046 13890
rect 15046 13838 15092 13890
rect 15116 13838 15162 13890
rect 15162 13838 15172 13890
rect 15196 13838 15226 13890
rect 15226 13838 15252 13890
rect 14956 13836 15012 13838
rect 15036 13836 15092 13838
rect 15116 13836 15172 13838
rect 15196 13836 15252 13838
rect 14956 12802 15012 12804
rect 15036 12802 15092 12804
rect 15116 12802 15172 12804
rect 15196 12802 15252 12804
rect 14956 12750 14982 12802
rect 14982 12750 15012 12802
rect 15036 12750 15046 12802
rect 15046 12750 15092 12802
rect 15116 12750 15162 12802
rect 15162 12750 15172 12802
rect 15196 12750 15226 12802
rect 15226 12750 15252 12802
rect 14956 12748 15012 12750
rect 15036 12748 15092 12750
rect 15116 12748 15172 12750
rect 15196 12748 15252 12750
rect 14956 11714 15012 11716
rect 15036 11714 15092 11716
rect 15116 11714 15172 11716
rect 15196 11714 15252 11716
rect 14956 11662 14982 11714
rect 14982 11662 15012 11714
rect 15036 11662 15046 11714
rect 15046 11662 15092 11714
rect 15116 11662 15162 11714
rect 15162 11662 15172 11714
rect 15196 11662 15226 11714
rect 15226 11662 15252 11714
rect 14956 11660 15012 11662
rect 15036 11660 15092 11662
rect 15116 11660 15172 11662
rect 15196 11660 15252 11662
rect 13542 10912 13598 10968
rect 5622 10626 5678 10628
rect 5702 10626 5758 10628
rect 5782 10626 5838 10628
rect 5862 10626 5918 10628
rect 5622 10574 5648 10626
rect 5648 10574 5678 10626
rect 5702 10574 5712 10626
rect 5712 10574 5758 10626
rect 5782 10574 5828 10626
rect 5828 10574 5838 10626
rect 5862 10574 5892 10626
rect 5892 10574 5918 10626
rect 5622 10572 5678 10574
rect 5702 10572 5758 10574
rect 5782 10572 5838 10574
rect 5862 10572 5918 10574
rect 14956 10626 15012 10628
rect 15036 10626 15092 10628
rect 15116 10626 15172 10628
rect 15196 10626 15252 10628
rect 14956 10574 14982 10626
rect 14982 10574 15012 10626
rect 15036 10574 15046 10626
rect 15046 10574 15092 10626
rect 15116 10574 15162 10626
rect 15162 10574 15172 10626
rect 15196 10574 15226 10626
rect 15226 10574 15252 10626
rect 14956 10572 15012 10574
rect 15036 10572 15092 10574
rect 15116 10572 15172 10574
rect 15196 10572 15252 10574
rect 10289 10082 10345 10084
rect 10369 10082 10425 10084
rect 10449 10082 10505 10084
rect 10529 10082 10585 10084
rect 10289 10030 10315 10082
rect 10315 10030 10345 10082
rect 10369 10030 10379 10082
rect 10379 10030 10425 10082
rect 10449 10030 10495 10082
rect 10495 10030 10505 10082
rect 10529 10030 10559 10082
rect 10559 10030 10585 10082
rect 10289 10028 10345 10030
rect 10369 10028 10425 10030
rect 10449 10028 10505 10030
rect 10529 10028 10585 10030
rect 5622 9538 5678 9540
rect 5702 9538 5758 9540
rect 5782 9538 5838 9540
rect 5862 9538 5918 9540
rect 5622 9486 5648 9538
rect 5648 9486 5678 9538
rect 5702 9486 5712 9538
rect 5712 9486 5758 9538
rect 5782 9486 5828 9538
rect 5828 9486 5838 9538
rect 5862 9486 5892 9538
rect 5892 9486 5918 9538
rect 5622 9484 5678 9486
rect 5702 9484 5758 9486
rect 5782 9484 5838 9486
rect 5862 9484 5918 9486
rect 10289 8994 10345 8996
rect 10369 8994 10425 8996
rect 10449 8994 10505 8996
rect 10529 8994 10585 8996
rect 10289 8942 10315 8994
rect 10315 8942 10345 8994
rect 10369 8942 10379 8994
rect 10379 8942 10425 8994
rect 10449 8942 10495 8994
rect 10495 8942 10505 8994
rect 10529 8942 10559 8994
rect 10559 8942 10585 8994
rect 10289 8940 10345 8942
rect 10369 8940 10425 8942
rect 10449 8940 10505 8942
rect 10529 8940 10585 8942
rect 5622 8450 5678 8452
rect 5702 8450 5758 8452
rect 5782 8450 5838 8452
rect 5862 8450 5918 8452
rect 5622 8398 5648 8450
rect 5648 8398 5678 8450
rect 5702 8398 5712 8450
rect 5712 8398 5758 8450
rect 5782 8398 5828 8450
rect 5828 8398 5838 8450
rect 5862 8398 5892 8450
rect 5892 8398 5918 8450
rect 5622 8396 5678 8398
rect 5702 8396 5758 8398
rect 5782 8396 5838 8398
rect 5862 8396 5918 8398
rect 10289 7906 10345 7908
rect 10369 7906 10425 7908
rect 10449 7906 10505 7908
rect 10529 7906 10585 7908
rect 10289 7854 10315 7906
rect 10315 7854 10345 7906
rect 10369 7854 10379 7906
rect 10379 7854 10425 7906
rect 10449 7854 10495 7906
rect 10495 7854 10505 7906
rect 10529 7854 10559 7906
rect 10559 7854 10585 7906
rect 10289 7852 10345 7854
rect 10369 7852 10425 7854
rect 10449 7852 10505 7854
rect 10529 7852 10585 7854
rect 5622 7362 5678 7364
rect 5702 7362 5758 7364
rect 5782 7362 5838 7364
rect 5862 7362 5918 7364
rect 5622 7310 5648 7362
rect 5648 7310 5678 7362
rect 5702 7310 5712 7362
rect 5712 7310 5758 7362
rect 5782 7310 5828 7362
rect 5828 7310 5838 7362
rect 5862 7310 5892 7362
rect 5892 7310 5918 7362
rect 5622 7308 5678 7310
rect 5702 7308 5758 7310
rect 5782 7308 5838 7310
rect 5862 7308 5918 7310
rect 10289 6818 10345 6820
rect 10369 6818 10425 6820
rect 10449 6818 10505 6820
rect 10529 6818 10585 6820
rect 10289 6766 10315 6818
rect 10315 6766 10345 6818
rect 10369 6766 10379 6818
rect 10379 6766 10425 6818
rect 10449 6766 10495 6818
rect 10495 6766 10505 6818
rect 10529 6766 10559 6818
rect 10559 6766 10585 6818
rect 10289 6764 10345 6766
rect 10369 6764 10425 6766
rect 10449 6764 10505 6766
rect 10529 6764 10585 6766
rect 3422 6696 3478 6752
rect 5622 6274 5678 6276
rect 5702 6274 5758 6276
rect 5782 6274 5838 6276
rect 5862 6274 5918 6276
rect 5622 6222 5648 6274
rect 5648 6222 5678 6274
rect 5702 6222 5712 6274
rect 5712 6222 5758 6274
rect 5782 6222 5828 6274
rect 5828 6222 5838 6274
rect 5862 6222 5892 6274
rect 5892 6222 5918 6274
rect 5622 6220 5678 6222
rect 5702 6220 5758 6222
rect 5782 6220 5838 6222
rect 5862 6220 5918 6222
rect 14956 9538 15012 9540
rect 15036 9538 15092 9540
rect 15116 9538 15172 9540
rect 15196 9538 15252 9540
rect 14956 9486 14982 9538
rect 14982 9486 15012 9538
rect 15036 9486 15046 9538
rect 15046 9486 15092 9538
rect 15116 9486 15162 9538
rect 15162 9486 15172 9538
rect 15196 9486 15226 9538
rect 15226 9486 15252 9538
rect 14956 9484 15012 9486
rect 15036 9484 15092 9486
rect 15116 9484 15172 9486
rect 15196 9484 15252 9486
rect 14956 8450 15012 8452
rect 15036 8450 15092 8452
rect 15116 8450 15172 8452
rect 15196 8450 15252 8452
rect 14956 8398 14982 8450
rect 14982 8398 15012 8450
rect 15036 8398 15046 8450
rect 15046 8398 15092 8450
rect 15116 8398 15162 8450
rect 15162 8398 15172 8450
rect 15196 8398 15226 8450
rect 15226 8398 15252 8450
rect 14956 8396 15012 8398
rect 15036 8396 15092 8398
rect 15116 8396 15172 8398
rect 15196 8396 15252 8398
rect 15658 7648 15714 7704
rect 14956 7362 15012 7364
rect 15036 7362 15092 7364
rect 15116 7362 15172 7364
rect 15196 7362 15252 7364
rect 14956 7310 14982 7362
rect 14982 7310 15012 7362
rect 15036 7310 15046 7362
rect 15046 7310 15092 7362
rect 15116 7310 15162 7362
rect 15162 7310 15172 7362
rect 15196 7310 15226 7362
rect 15226 7310 15252 7362
rect 14956 7308 15012 7310
rect 15036 7308 15092 7310
rect 15116 7308 15172 7310
rect 15196 7308 15252 7310
rect 14956 6274 15012 6276
rect 15036 6274 15092 6276
rect 15116 6274 15172 6276
rect 15196 6274 15252 6276
rect 14956 6222 14982 6274
rect 14982 6222 15012 6274
rect 15036 6222 15046 6274
rect 15046 6222 15092 6274
rect 15116 6222 15162 6274
rect 15162 6222 15172 6274
rect 15196 6222 15226 6274
rect 15226 6222 15252 6274
rect 14956 6220 15012 6222
rect 15036 6220 15092 6222
rect 15116 6220 15172 6222
rect 15196 6220 15252 6222
rect 13174 6016 13230 6072
rect 10289 5730 10345 5732
rect 10369 5730 10425 5732
rect 10449 5730 10505 5732
rect 10529 5730 10585 5732
rect 10289 5678 10315 5730
rect 10315 5678 10345 5730
rect 10369 5678 10379 5730
rect 10379 5678 10425 5730
rect 10449 5678 10495 5730
rect 10495 5678 10505 5730
rect 10529 5678 10559 5730
rect 10559 5678 10585 5730
rect 10289 5676 10345 5678
rect 10369 5676 10425 5678
rect 10449 5676 10505 5678
rect 10529 5676 10585 5678
rect 5622 5186 5678 5188
rect 5702 5186 5758 5188
rect 5782 5186 5838 5188
rect 5862 5186 5918 5188
rect 5622 5134 5648 5186
rect 5648 5134 5678 5186
rect 5702 5134 5712 5186
rect 5712 5134 5758 5186
rect 5782 5134 5828 5186
rect 5828 5134 5838 5186
rect 5862 5134 5892 5186
rect 5892 5134 5918 5186
rect 5622 5132 5678 5134
rect 5702 5132 5758 5134
rect 5782 5132 5838 5134
rect 5862 5132 5918 5134
rect 14956 5186 15012 5188
rect 15036 5186 15092 5188
rect 15116 5186 15172 5188
rect 15196 5186 15252 5188
rect 14956 5134 14982 5186
rect 14982 5134 15012 5186
rect 15036 5134 15046 5186
rect 15046 5134 15092 5186
rect 15116 5134 15162 5186
rect 15162 5134 15172 5186
rect 15196 5134 15226 5186
rect 15226 5134 15252 5186
rect 14956 5132 15012 5134
rect 15036 5132 15092 5134
rect 15116 5132 15172 5134
rect 15196 5132 15252 5134
rect 16394 22764 16450 22800
rect 16394 22744 16396 22764
rect 16396 22744 16448 22764
rect 16448 22744 16450 22764
rect 16394 19208 16450 19264
rect 16394 17884 16396 17904
rect 16396 17884 16448 17904
rect 16448 17884 16450 17904
rect 16394 17848 16450 17884
rect 16486 17576 16542 17632
rect 16394 15420 16450 15456
rect 16394 15400 16396 15420
rect 16396 15400 16448 15420
rect 16448 15400 16450 15420
rect 16302 14992 16358 15048
rect 16394 13788 16450 13824
rect 16394 13768 16396 13788
rect 16396 13768 16448 13788
rect 16448 13768 16450 13788
rect 16854 19208 16910 19264
rect 18418 24104 18474 24160
rect 18142 23580 18198 23616
rect 18142 23560 18144 23580
rect 18144 23560 18196 23580
rect 18196 23560 18198 23580
rect 18786 23560 18842 23616
rect 18142 22492 18198 22528
rect 18142 22472 18144 22492
rect 18144 22472 18196 22492
rect 18196 22472 18198 22492
rect 18418 22064 18474 22120
rect 18326 21812 18382 21848
rect 18326 21792 18328 21812
rect 18328 21792 18380 21812
rect 18380 21792 18382 21812
rect 18326 21656 18382 21712
rect 18326 21248 18382 21304
rect 17038 20840 17094 20896
rect 17958 20704 18014 20760
rect 17590 20024 17646 20080
rect 18510 17596 18566 17632
rect 18510 17576 18512 17596
rect 18512 17576 18564 17596
rect 18564 17576 18566 17596
rect 18418 17460 18474 17496
rect 18418 17440 18420 17460
rect 18420 17440 18472 17460
rect 18472 17440 18474 17460
rect 18418 16916 18474 16952
rect 18418 16896 18420 16916
rect 18420 16896 18472 16916
rect 18472 16896 18474 16916
rect 18694 16760 18750 16816
rect 18970 19636 19026 19672
rect 18970 19616 18972 19636
rect 18972 19616 19024 19636
rect 19024 19616 19026 19636
rect 18418 15536 18474 15592
rect 19062 16352 19118 16408
rect 18694 15672 18750 15728
rect 18694 14176 18750 14232
rect 17774 7260 17830 7296
rect 17774 7240 17776 7260
rect 17776 7240 17828 7260
rect 17828 7240 17830 7260
rect 16854 5900 16910 5936
rect 16854 5880 16856 5900
rect 16856 5880 16908 5900
rect 16908 5880 16910 5900
rect 15934 4812 15990 4848
rect 15934 4792 15936 4812
rect 15936 4792 15988 4812
rect 15988 4792 15990 4812
rect 10289 4642 10345 4644
rect 10369 4642 10425 4644
rect 10449 4642 10505 4644
rect 10529 4642 10585 4644
rect 10289 4590 10315 4642
rect 10315 4590 10345 4642
rect 10369 4590 10379 4642
rect 10379 4590 10425 4642
rect 10449 4590 10495 4642
rect 10495 4590 10505 4642
rect 10529 4590 10559 4642
rect 10559 4590 10585 4642
rect 10289 4588 10345 4590
rect 10369 4588 10425 4590
rect 10449 4588 10505 4590
rect 10529 4588 10585 4590
rect 19062 14740 19118 14776
rect 19062 14720 19064 14740
rect 19064 14720 19116 14740
rect 19116 14720 19118 14740
rect 18878 13632 18934 13688
rect 19622 25314 19678 25316
rect 19702 25314 19758 25316
rect 19782 25314 19838 25316
rect 19862 25314 19918 25316
rect 19622 25262 19648 25314
rect 19648 25262 19678 25314
rect 19702 25262 19712 25314
rect 19712 25262 19758 25314
rect 19782 25262 19828 25314
rect 19828 25262 19838 25314
rect 19862 25262 19892 25314
rect 19892 25262 19918 25314
rect 19622 25260 19678 25262
rect 19702 25260 19758 25262
rect 19782 25260 19838 25262
rect 19862 25260 19918 25262
rect 19622 24226 19678 24228
rect 19702 24226 19758 24228
rect 19782 24226 19838 24228
rect 19862 24226 19918 24228
rect 19622 24174 19648 24226
rect 19648 24174 19678 24226
rect 19702 24174 19712 24226
rect 19712 24174 19758 24226
rect 19782 24174 19828 24226
rect 19828 24174 19838 24226
rect 19862 24174 19892 24226
rect 19892 24174 19918 24226
rect 19622 24172 19678 24174
rect 19702 24172 19758 24174
rect 19782 24172 19838 24174
rect 19862 24172 19918 24174
rect 19982 23852 20038 23888
rect 19982 23832 19984 23852
rect 19984 23832 20036 23852
rect 20036 23832 20038 23852
rect 19622 23138 19678 23140
rect 19702 23138 19758 23140
rect 19782 23138 19838 23140
rect 19862 23138 19918 23140
rect 19622 23086 19648 23138
rect 19648 23086 19678 23138
rect 19702 23086 19712 23138
rect 19712 23086 19758 23138
rect 19782 23086 19828 23138
rect 19828 23086 19838 23138
rect 19862 23086 19892 23138
rect 19892 23086 19918 23138
rect 19622 23084 19678 23086
rect 19702 23084 19758 23086
rect 19782 23084 19838 23086
rect 19862 23084 19918 23086
rect 19622 22050 19678 22052
rect 19702 22050 19758 22052
rect 19782 22050 19838 22052
rect 19862 22050 19918 22052
rect 19622 21998 19648 22050
rect 19648 21998 19678 22050
rect 19702 21998 19712 22050
rect 19712 21998 19758 22050
rect 19782 21998 19828 22050
rect 19828 21998 19838 22050
rect 19862 21998 19892 22050
rect 19892 21998 19918 22050
rect 19622 21996 19678 21998
rect 19702 21996 19758 21998
rect 19782 21996 19838 21998
rect 19862 21996 19918 21998
rect 19622 20962 19678 20964
rect 19702 20962 19758 20964
rect 19782 20962 19838 20964
rect 19862 20962 19918 20964
rect 19622 20910 19648 20962
rect 19648 20910 19678 20962
rect 19702 20910 19712 20962
rect 19712 20910 19758 20962
rect 19782 20910 19828 20962
rect 19828 20910 19838 20962
rect 19862 20910 19892 20962
rect 19892 20910 19918 20962
rect 19622 20908 19678 20910
rect 19702 20908 19758 20910
rect 19782 20908 19838 20910
rect 19862 20908 19918 20910
rect 19622 19874 19678 19876
rect 19702 19874 19758 19876
rect 19782 19874 19838 19876
rect 19862 19874 19918 19876
rect 19622 19822 19648 19874
rect 19648 19822 19678 19874
rect 19702 19822 19712 19874
rect 19712 19822 19758 19874
rect 19782 19822 19828 19874
rect 19828 19822 19838 19874
rect 19862 19822 19892 19874
rect 19892 19822 19918 19874
rect 19622 19820 19678 19822
rect 19702 19820 19758 19822
rect 19782 19820 19838 19822
rect 19862 19820 19918 19822
rect 19622 18786 19678 18788
rect 19702 18786 19758 18788
rect 19782 18786 19838 18788
rect 19862 18786 19918 18788
rect 19622 18734 19648 18786
rect 19648 18734 19678 18786
rect 19702 18734 19712 18786
rect 19712 18734 19758 18786
rect 19782 18734 19828 18786
rect 19828 18734 19838 18786
rect 19862 18734 19892 18786
rect 19892 18734 19918 18786
rect 19622 18732 19678 18734
rect 19702 18732 19758 18734
rect 19782 18732 19838 18734
rect 19862 18732 19918 18734
rect 19622 17698 19678 17700
rect 19702 17698 19758 17700
rect 19782 17698 19838 17700
rect 19862 17698 19918 17700
rect 19622 17646 19648 17698
rect 19648 17646 19678 17698
rect 19702 17646 19712 17698
rect 19712 17646 19758 17698
rect 19782 17646 19828 17698
rect 19828 17646 19838 17698
rect 19862 17646 19892 17698
rect 19892 17646 19918 17698
rect 19622 17644 19678 17646
rect 19702 17644 19758 17646
rect 19782 17644 19838 17646
rect 19862 17644 19918 17646
rect 20994 22492 21050 22528
rect 20994 22472 20996 22492
rect 20996 22472 21048 22492
rect 21048 22472 21050 22492
rect 20718 22220 20774 22256
rect 20718 22200 20720 22220
rect 20720 22200 20772 22220
rect 20772 22200 20774 22220
rect 19622 16610 19678 16612
rect 19702 16610 19758 16612
rect 19782 16610 19838 16612
rect 19862 16610 19918 16612
rect 19622 16558 19648 16610
rect 19648 16558 19678 16610
rect 19702 16558 19712 16610
rect 19712 16558 19758 16610
rect 19782 16558 19828 16610
rect 19828 16558 19838 16610
rect 19862 16558 19892 16610
rect 19892 16558 19918 16610
rect 19622 16556 19678 16558
rect 19702 16556 19758 16558
rect 19782 16556 19838 16558
rect 19862 16556 19918 16558
rect 19622 15522 19678 15524
rect 19702 15522 19758 15524
rect 19782 15522 19838 15524
rect 19862 15522 19918 15524
rect 19622 15470 19648 15522
rect 19648 15470 19678 15522
rect 19702 15470 19712 15522
rect 19712 15470 19758 15522
rect 19782 15470 19828 15522
rect 19828 15470 19838 15522
rect 19862 15470 19892 15522
rect 19892 15470 19918 15522
rect 19622 15468 19678 15470
rect 19702 15468 19758 15470
rect 19782 15468 19838 15470
rect 19862 15468 19918 15470
rect 19622 14434 19678 14436
rect 19702 14434 19758 14436
rect 19782 14434 19838 14436
rect 19862 14434 19918 14436
rect 19622 14382 19648 14434
rect 19648 14382 19678 14434
rect 19702 14382 19712 14434
rect 19712 14382 19758 14434
rect 19782 14382 19828 14434
rect 19828 14382 19838 14434
rect 19862 14382 19892 14434
rect 19892 14382 19918 14434
rect 19622 14380 19678 14382
rect 19702 14380 19758 14382
rect 19782 14380 19838 14382
rect 19862 14380 19918 14382
rect 20258 13788 20314 13824
rect 20258 13768 20260 13788
rect 20260 13768 20312 13788
rect 20312 13768 20314 13788
rect 19622 13346 19678 13348
rect 19702 13346 19758 13348
rect 19782 13346 19838 13348
rect 19862 13346 19918 13348
rect 19622 13294 19648 13346
rect 19648 13294 19678 13346
rect 19702 13294 19712 13346
rect 19712 13294 19758 13346
rect 19782 13294 19828 13346
rect 19828 13294 19838 13346
rect 19862 13294 19892 13346
rect 19892 13294 19918 13346
rect 19622 13292 19678 13294
rect 19702 13292 19758 13294
rect 19782 13292 19838 13294
rect 19862 13292 19918 13294
rect 19246 13088 19302 13144
rect 19622 12258 19678 12260
rect 19702 12258 19758 12260
rect 19782 12258 19838 12260
rect 19862 12258 19918 12260
rect 19622 12206 19648 12258
rect 19648 12206 19678 12258
rect 19702 12206 19712 12258
rect 19712 12206 19758 12258
rect 19782 12206 19828 12258
rect 19828 12206 19838 12258
rect 19862 12206 19892 12258
rect 19892 12206 19918 12258
rect 19622 12204 19678 12206
rect 19702 12204 19758 12206
rect 19782 12204 19838 12206
rect 19862 12204 19918 12206
rect 19246 11456 19302 11512
rect 19154 7512 19210 7568
rect 18694 7240 18750 7296
rect 18234 7124 18290 7160
rect 18234 7104 18236 7124
rect 18236 7104 18288 7124
rect 18288 7104 18290 7124
rect 19622 11170 19678 11172
rect 19702 11170 19758 11172
rect 19782 11170 19838 11172
rect 19862 11170 19918 11172
rect 19622 11118 19648 11170
rect 19648 11118 19678 11170
rect 19702 11118 19712 11170
rect 19712 11118 19758 11170
rect 19782 11118 19828 11170
rect 19828 11118 19838 11170
rect 19862 11118 19892 11170
rect 19892 11118 19918 11170
rect 19622 11116 19678 11118
rect 19702 11116 19758 11118
rect 19782 11116 19838 11118
rect 19862 11116 19918 11118
rect 19622 10082 19678 10084
rect 19702 10082 19758 10084
rect 19782 10082 19838 10084
rect 19862 10082 19918 10084
rect 19622 10030 19648 10082
rect 19648 10030 19678 10082
rect 19702 10030 19712 10082
rect 19712 10030 19758 10082
rect 19782 10030 19828 10082
rect 19828 10030 19838 10082
rect 19862 10030 19892 10082
rect 19892 10030 19918 10082
rect 19622 10028 19678 10030
rect 19702 10028 19758 10030
rect 19782 10028 19838 10030
rect 19862 10028 19918 10030
rect 20442 9280 20498 9336
rect 20902 20704 20958 20760
rect 20718 18392 20774 18448
rect 20718 14740 20774 14776
rect 20718 14720 20720 14740
rect 20720 14720 20772 14740
rect 20772 14720 20774 14740
rect 21362 22472 21418 22528
rect 21546 19208 21602 19264
rect 21178 17304 21234 17360
rect 21638 18800 21694 18856
rect 21822 17712 21878 17768
rect 21730 17440 21786 17496
rect 21914 16488 21970 16544
rect 21362 14992 21418 15048
rect 20902 13632 20958 13688
rect 21454 11456 21510 11512
rect 21178 11356 21180 11376
rect 21180 11356 21232 11376
rect 21232 11356 21234 11376
rect 21178 11320 21234 11356
rect 20626 9008 20682 9064
rect 19622 8994 19678 8996
rect 19702 8994 19758 8996
rect 19782 8994 19838 8996
rect 19862 8994 19918 8996
rect 19622 8942 19648 8994
rect 19648 8942 19678 8994
rect 19702 8942 19712 8994
rect 19712 8942 19758 8994
rect 19782 8942 19828 8994
rect 19828 8942 19838 8994
rect 19862 8942 19892 8994
rect 19892 8942 19918 8994
rect 19622 8940 19678 8942
rect 19702 8940 19758 8942
rect 19782 8940 19838 8942
rect 19862 8940 19918 8942
rect 19622 7906 19678 7908
rect 19702 7906 19758 7908
rect 19782 7906 19838 7908
rect 19862 7906 19918 7908
rect 19622 7854 19648 7906
rect 19648 7854 19678 7906
rect 19702 7854 19712 7906
rect 19712 7854 19758 7906
rect 19782 7854 19828 7906
rect 19828 7854 19838 7906
rect 19862 7854 19892 7906
rect 19892 7854 19918 7906
rect 19622 7852 19678 7854
rect 19702 7852 19758 7854
rect 19782 7852 19838 7854
rect 19862 7852 19918 7854
rect 19622 6818 19678 6820
rect 19702 6818 19758 6820
rect 19782 6818 19838 6820
rect 19862 6818 19918 6820
rect 19622 6766 19648 6818
rect 19648 6766 19678 6818
rect 19702 6766 19712 6818
rect 19712 6766 19758 6818
rect 19782 6766 19828 6818
rect 19828 6766 19838 6818
rect 19862 6766 19892 6818
rect 19892 6766 19918 6818
rect 19622 6764 19678 6766
rect 19702 6764 19758 6766
rect 19782 6764 19838 6766
rect 19862 6764 19918 6766
rect 19622 5730 19678 5732
rect 19702 5730 19758 5732
rect 19782 5730 19838 5732
rect 19862 5730 19918 5732
rect 19622 5678 19648 5730
rect 19648 5678 19678 5730
rect 19702 5678 19712 5730
rect 19712 5678 19758 5730
rect 19782 5678 19828 5730
rect 19828 5678 19838 5730
rect 19862 5678 19892 5730
rect 19892 5678 19918 5730
rect 19622 5676 19678 5678
rect 19702 5676 19758 5678
rect 19782 5676 19838 5678
rect 19862 5676 19918 5678
rect 19246 5336 19302 5392
rect 22558 24412 22560 24432
rect 22560 24412 22612 24432
rect 22612 24412 22614 24432
rect 22558 24376 22614 24412
rect 22834 24548 22836 24568
rect 22836 24548 22888 24568
rect 22888 24548 22890 24568
rect 22834 24512 22890 24548
rect 22098 23560 22154 23616
rect 22374 23308 22430 23344
rect 22374 23288 22376 23308
rect 22376 23288 22428 23308
rect 22428 23288 22430 23308
rect 22282 22608 22338 22664
rect 23386 26144 23442 26200
rect 23294 25600 23350 25656
rect 22926 21656 22982 21712
rect 23570 26824 23626 26880
rect 24289 24770 24345 24772
rect 24369 24770 24425 24772
rect 24449 24770 24505 24772
rect 24529 24770 24585 24772
rect 24289 24718 24315 24770
rect 24315 24718 24345 24770
rect 24369 24718 24379 24770
rect 24379 24718 24425 24770
rect 24449 24718 24495 24770
rect 24495 24718 24505 24770
rect 24529 24718 24559 24770
rect 24559 24718 24585 24770
rect 24289 24716 24345 24718
rect 24369 24716 24425 24718
rect 24449 24716 24505 24718
rect 24529 24716 24585 24718
rect 24766 25056 24822 25112
rect 22098 19108 22100 19128
rect 22100 19108 22152 19128
rect 22152 19108 22154 19128
rect 22098 19072 22154 19108
rect 23294 18800 23350 18856
rect 22190 16352 22246 16408
rect 22926 10640 22982 10696
rect 22006 10504 22062 10560
rect 23662 21384 23718 21440
rect 23662 20568 23718 20624
rect 23846 22744 23902 22800
rect 23846 22608 23902 22664
rect 23938 22492 23994 22528
rect 23938 22472 23940 22492
rect 23940 22472 23992 22492
rect 23992 22472 23994 22492
rect 25134 24376 25190 24432
rect 24289 23682 24345 23684
rect 24369 23682 24425 23684
rect 24449 23682 24505 23684
rect 24529 23682 24585 23684
rect 24289 23630 24315 23682
rect 24315 23630 24345 23682
rect 24369 23630 24379 23682
rect 24379 23630 24425 23682
rect 24449 23630 24495 23682
rect 24495 23630 24505 23682
rect 24529 23630 24559 23682
rect 24559 23630 24585 23682
rect 24289 23628 24345 23630
rect 24369 23628 24425 23630
rect 24449 23628 24505 23630
rect 24529 23628 24585 23630
rect 25134 23852 25190 23888
rect 25134 23832 25136 23852
rect 25136 23832 25188 23852
rect 25188 23832 25190 23852
rect 24674 22608 24730 22664
rect 24289 22594 24345 22596
rect 24369 22594 24425 22596
rect 24449 22594 24505 22596
rect 24529 22594 24585 22596
rect 24289 22542 24315 22594
rect 24315 22542 24345 22594
rect 24369 22542 24379 22594
rect 24379 22542 24425 22594
rect 24449 22542 24495 22594
rect 24495 22542 24505 22594
rect 24529 22542 24559 22594
rect 24559 22542 24585 22594
rect 24289 22540 24345 22542
rect 24369 22540 24425 22542
rect 24449 22540 24505 22542
rect 24529 22540 24585 22542
rect 24766 22336 24822 22392
rect 24674 21656 24730 21712
rect 24122 21520 24178 21576
rect 24289 21506 24345 21508
rect 24369 21506 24425 21508
rect 24449 21506 24505 21508
rect 24529 21506 24585 21508
rect 24289 21454 24315 21506
rect 24315 21454 24345 21506
rect 24369 21454 24379 21506
rect 24379 21454 24425 21506
rect 24449 21454 24495 21506
rect 24495 21454 24505 21506
rect 24529 21454 24559 21506
rect 24559 21454 24585 21506
rect 24289 21452 24345 21454
rect 24369 21452 24425 21454
rect 24449 21452 24505 21454
rect 24529 21452 24585 21454
rect 24766 21384 24822 21440
rect 23846 20724 23902 20760
rect 23846 20704 23848 20724
rect 23848 20704 23900 20724
rect 23900 20704 23902 20724
rect 23754 18120 23810 18176
rect 23662 17748 23664 17768
rect 23664 17748 23716 17768
rect 23716 17748 23718 17768
rect 23662 17712 23718 17748
rect 23662 15264 23718 15320
rect 23386 14992 23442 15048
rect 23662 14196 23718 14232
rect 23662 14176 23664 14196
rect 23664 14176 23716 14196
rect 23716 14176 23718 14196
rect 23478 6560 23534 6616
rect 23478 5336 23534 5392
rect 21546 4928 21602 4984
rect 23478 4656 23534 4712
rect 19622 4642 19678 4644
rect 19702 4642 19758 4644
rect 19782 4642 19838 4644
rect 19862 4642 19918 4644
rect 19622 4590 19648 4642
rect 19648 4590 19678 4642
rect 19702 4590 19712 4642
rect 19712 4590 19758 4642
rect 19782 4590 19828 4642
rect 19828 4590 19838 4642
rect 19862 4590 19892 4642
rect 19892 4590 19918 4642
rect 19622 4588 19678 4590
rect 19702 4588 19758 4590
rect 19782 4588 19838 4590
rect 19862 4588 19918 4590
rect 17958 4248 18014 4304
rect 5622 4098 5678 4100
rect 5702 4098 5758 4100
rect 5782 4098 5838 4100
rect 5862 4098 5918 4100
rect 5622 4046 5648 4098
rect 5648 4046 5678 4098
rect 5702 4046 5712 4098
rect 5712 4046 5758 4098
rect 5782 4046 5828 4098
rect 5828 4046 5838 4098
rect 5862 4046 5892 4098
rect 5892 4046 5918 4098
rect 5622 4044 5678 4046
rect 5702 4044 5758 4046
rect 5782 4044 5838 4046
rect 5862 4044 5918 4046
rect 14956 4098 15012 4100
rect 15036 4098 15092 4100
rect 15116 4098 15172 4100
rect 15196 4098 15252 4100
rect 14956 4046 14982 4098
rect 14982 4046 15012 4098
rect 15036 4046 15046 4098
rect 15046 4046 15092 4098
rect 15116 4046 15162 4098
rect 15162 4046 15172 4098
rect 15196 4046 15226 4098
rect 15226 4046 15252 4098
rect 14956 4044 15012 4046
rect 15036 4044 15092 4046
rect 15116 4044 15172 4046
rect 15196 4044 15252 4046
rect 10289 3554 10345 3556
rect 10369 3554 10425 3556
rect 10449 3554 10505 3556
rect 10529 3554 10585 3556
rect 10289 3502 10315 3554
rect 10315 3502 10345 3554
rect 10369 3502 10379 3554
rect 10379 3502 10425 3554
rect 10449 3502 10495 3554
rect 10495 3502 10505 3554
rect 10529 3502 10559 3554
rect 10559 3502 10585 3554
rect 10289 3500 10345 3502
rect 10369 3500 10425 3502
rect 10449 3500 10505 3502
rect 10529 3500 10585 3502
rect 19622 3554 19678 3556
rect 19702 3554 19758 3556
rect 19782 3554 19838 3556
rect 19862 3554 19918 3556
rect 19622 3502 19648 3554
rect 19648 3502 19678 3554
rect 19702 3502 19712 3554
rect 19712 3502 19758 3554
rect 19782 3502 19828 3554
rect 19828 3502 19838 3554
rect 19862 3502 19892 3554
rect 19892 3502 19918 3554
rect 19622 3500 19678 3502
rect 19702 3500 19758 3502
rect 19782 3500 19838 3502
rect 19862 3500 19918 3502
rect 5622 3010 5678 3012
rect 5702 3010 5758 3012
rect 5782 3010 5838 3012
rect 5862 3010 5918 3012
rect 5622 2958 5648 3010
rect 5648 2958 5678 3010
rect 5702 2958 5712 3010
rect 5712 2958 5758 3010
rect 5782 2958 5828 3010
rect 5828 2958 5838 3010
rect 5862 2958 5892 3010
rect 5892 2958 5918 3010
rect 5622 2956 5678 2958
rect 5702 2956 5758 2958
rect 5782 2956 5838 2958
rect 5862 2956 5918 2958
rect 14956 3010 15012 3012
rect 15036 3010 15092 3012
rect 15116 3010 15172 3012
rect 15196 3010 15252 3012
rect 14956 2958 14982 3010
rect 14982 2958 15012 3010
rect 15036 2958 15046 3010
rect 15046 2958 15092 3010
rect 15116 2958 15162 3010
rect 15162 2958 15172 3010
rect 15196 2958 15226 3010
rect 15226 2958 15252 3010
rect 14956 2956 15012 2958
rect 15036 2956 15092 2958
rect 15116 2956 15172 2958
rect 15196 2956 15252 2958
rect 10289 2466 10345 2468
rect 10369 2466 10425 2468
rect 10449 2466 10505 2468
rect 10529 2466 10585 2468
rect 10289 2414 10315 2466
rect 10315 2414 10345 2466
rect 10369 2414 10379 2466
rect 10379 2414 10425 2466
rect 10449 2414 10495 2466
rect 10495 2414 10505 2466
rect 10529 2414 10559 2466
rect 10559 2414 10585 2466
rect 10289 2412 10345 2414
rect 10369 2412 10425 2414
rect 10449 2412 10505 2414
rect 10529 2412 10585 2414
rect 19622 2466 19678 2468
rect 19702 2466 19758 2468
rect 19782 2466 19838 2468
rect 19862 2466 19918 2468
rect 19622 2414 19648 2466
rect 19648 2414 19678 2466
rect 19702 2414 19712 2466
rect 19712 2414 19758 2466
rect 19782 2414 19828 2466
rect 19828 2414 19838 2466
rect 19862 2414 19892 2466
rect 19892 2414 19918 2466
rect 19622 2412 19678 2414
rect 19702 2412 19758 2414
rect 19782 2412 19838 2414
rect 19862 2412 19918 2414
rect 23478 2344 23534 2400
rect 5622 1922 5678 1924
rect 5702 1922 5758 1924
rect 5782 1922 5838 1924
rect 5862 1922 5918 1924
rect 5622 1870 5648 1922
rect 5648 1870 5678 1922
rect 5702 1870 5712 1922
rect 5712 1870 5758 1922
rect 5782 1870 5828 1922
rect 5828 1870 5838 1922
rect 5862 1870 5892 1922
rect 5892 1870 5918 1922
rect 5622 1868 5678 1870
rect 5702 1868 5758 1870
rect 5782 1868 5838 1870
rect 5862 1868 5918 1870
rect 14956 1922 15012 1924
rect 15036 1922 15092 1924
rect 15116 1922 15172 1924
rect 15196 1922 15252 1924
rect 14956 1870 14982 1922
rect 14982 1870 15012 1922
rect 15036 1870 15046 1922
rect 15046 1870 15092 1922
rect 15116 1870 15162 1922
rect 15162 1870 15172 1922
rect 15196 1870 15226 1922
rect 15226 1870 15252 1922
rect 14956 1868 15012 1870
rect 15036 1868 15092 1870
rect 15116 1868 15172 1870
rect 15196 1868 15252 1870
rect 23662 7648 23718 7704
rect 23662 5336 23718 5392
rect 23662 4928 23718 4984
rect 23938 16796 23940 16816
rect 23940 16796 23992 16816
rect 23992 16796 23994 16816
rect 23938 16760 23994 16796
rect 24030 16488 24086 16544
rect 23938 13088 23994 13144
rect 24289 20418 24345 20420
rect 24369 20418 24425 20420
rect 24449 20418 24505 20420
rect 24529 20418 24585 20420
rect 24289 20366 24315 20418
rect 24315 20366 24345 20418
rect 24369 20366 24379 20418
rect 24379 20366 24425 20418
rect 24449 20366 24495 20418
rect 24495 20366 24505 20418
rect 24529 20366 24559 20418
rect 24559 20366 24585 20418
rect 24289 20364 24345 20366
rect 24369 20364 24425 20366
rect 24449 20364 24505 20366
rect 24529 20364 24585 20366
rect 24289 19330 24345 19332
rect 24369 19330 24425 19332
rect 24449 19330 24505 19332
rect 24529 19330 24585 19332
rect 24289 19278 24315 19330
rect 24315 19278 24345 19330
rect 24369 19278 24379 19330
rect 24379 19278 24425 19330
rect 24449 19278 24495 19330
rect 24495 19278 24505 19330
rect 24529 19278 24559 19330
rect 24559 19278 24585 19330
rect 24289 19276 24345 19278
rect 24369 19276 24425 19278
rect 24449 19276 24505 19278
rect 24529 19276 24585 19278
rect 24289 18242 24345 18244
rect 24369 18242 24425 18244
rect 24449 18242 24505 18244
rect 24529 18242 24585 18244
rect 24289 18190 24315 18242
rect 24315 18190 24345 18242
rect 24369 18190 24379 18242
rect 24379 18190 24425 18242
rect 24449 18190 24495 18242
rect 24495 18190 24505 18242
rect 24529 18190 24559 18242
rect 24559 18190 24585 18242
rect 24289 18188 24345 18190
rect 24369 18188 24425 18190
rect 24449 18188 24505 18190
rect 24529 18188 24585 18190
rect 24289 17154 24345 17156
rect 24369 17154 24425 17156
rect 24449 17154 24505 17156
rect 24529 17154 24585 17156
rect 24289 17102 24315 17154
rect 24315 17102 24345 17154
rect 24369 17102 24379 17154
rect 24379 17102 24425 17154
rect 24449 17102 24495 17154
rect 24495 17102 24505 17154
rect 24529 17102 24559 17154
rect 24559 17102 24585 17154
rect 24289 17100 24345 17102
rect 24369 17100 24425 17102
rect 24449 17100 24505 17102
rect 24529 17100 24585 17102
rect 24289 16066 24345 16068
rect 24369 16066 24425 16068
rect 24449 16066 24505 16068
rect 24529 16066 24585 16068
rect 24289 16014 24315 16066
rect 24315 16014 24345 16066
rect 24369 16014 24379 16066
rect 24379 16014 24425 16066
rect 24449 16014 24495 16066
rect 24495 16014 24505 16066
rect 24529 16014 24559 16066
rect 24559 16014 24585 16066
rect 24289 16012 24345 16014
rect 24369 16012 24425 16014
rect 24449 16012 24505 16014
rect 24529 16012 24585 16014
rect 24950 22100 24952 22120
rect 24952 22100 25004 22120
rect 25004 22100 25006 22120
rect 24950 22064 25006 22100
rect 25134 21148 25136 21168
rect 25136 21148 25188 21168
rect 25188 21148 25190 21168
rect 25134 21112 25190 21148
rect 25134 20316 25190 20352
rect 25134 20296 25136 20316
rect 25136 20296 25188 20316
rect 25188 20296 25190 20316
rect 24950 19616 25006 19672
rect 25134 19072 25190 19128
rect 24766 17848 24822 17904
rect 25502 23288 25558 23344
rect 25410 23036 25466 23072
rect 25410 23016 25412 23036
rect 25412 23016 25464 23036
rect 25464 23016 25466 23036
rect 25686 21792 25742 21848
rect 25318 20840 25374 20896
rect 25410 19616 25466 19672
rect 25594 20160 25650 20216
rect 25318 18392 25374 18448
rect 24766 16080 24822 16136
rect 24289 14978 24345 14980
rect 24369 14978 24425 14980
rect 24449 14978 24505 14980
rect 24529 14978 24585 14980
rect 24289 14926 24315 14978
rect 24315 14926 24345 14978
rect 24369 14926 24379 14978
rect 24379 14926 24425 14978
rect 24449 14926 24495 14978
rect 24495 14926 24505 14978
rect 24529 14926 24559 14978
rect 24559 14926 24585 14978
rect 24289 14924 24345 14926
rect 24369 14924 24425 14926
rect 24449 14924 24505 14926
rect 24529 14924 24585 14926
rect 24289 13890 24345 13892
rect 24369 13890 24425 13892
rect 24449 13890 24505 13892
rect 24529 13890 24585 13892
rect 24289 13838 24315 13890
rect 24315 13838 24345 13890
rect 24369 13838 24379 13890
rect 24379 13838 24425 13890
rect 24449 13838 24495 13890
rect 24495 13838 24505 13890
rect 24529 13838 24559 13890
rect 24559 13838 24585 13890
rect 24289 13836 24345 13838
rect 24369 13836 24425 13838
rect 24449 13836 24505 13838
rect 24529 13836 24585 13838
rect 24289 12802 24345 12804
rect 24369 12802 24425 12804
rect 24449 12802 24505 12804
rect 24529 12802 24585 12804
rect 24289 12750 24315 12802
rect 24315 12750 24345 12802
rect 24369 12750 24379 12802
rect 24379 12750 24425 12802
rect 24449 12750 24495 12802
rect 24495 12750 24505 12802
rect 24529 12750 24559 12802
rect 24559 12750 24585 12802
rect 24289 12748 24345 12750
rect 24369 12748 24425 12750
rect 24449 12748 24505 12750
rect 24529 12748 24585 12750
rect 24674 12564 24730 12600
rect 24674 12544 24676 12564
rect 24676 12544 24728 12564
rect 24728 12544 24730 12564
rect 24582 11864 24638 11920
rect 24289 11714 24345 11716
rect 24369 11714 24425 11716
rect 24449 11714 24505 11716
rect 24529 11714 24585 11716
rect 24289 11662 24315 11714
rect 24315 11662 24345 11714
rect 24369 11662 24379 11714
rect 24379 11662 24425 11714
rect 24449 11662 24495 11714
rect 24495 11662 24505 11714
rect 24529 11662 24559 11714
rect 24559 11662 24585 11714
rect 24289 11660 24345 11662
rect 24369 11660 24425 11662
rect 24449 11660 24505 11662
rect 24529 11660 24585 11662
rect 25410 17304 25466 17360
rect 25410 16624 25466 16680
rect 25502 15400 25558 15456
rect 25870 14876 25926 14912
rect 25870 14856 25872 14876
rect 25872 14856 25924 14876
rect 25924 14856 25926 14876
rect 25594 14312 25650 14368
rect 25226 13652 25282 13688
rect 25226 13632 25228 13652
rect 25228 13632 25280 13652
rect 25280 13632 25282 13652
rect 25042 13108 25098 13144
rect 25042 13088 25044 13108
rect 25044 13088 25096 13108
rect 25096 13088 25098 13108
rect 24030 10640 24086 10696
rect 24674 10640 24730 10696
rect 24289 10626 24345 10628
rect 24369 10626 24425 10628
rect 24449 10626 24505 10628
rect 24529 10626 24585 10628
rect 24289 10574 24315 10626
rect 24315 10574 24345 10626
rect 24369 10574 24379 10626
rect 24379 10574 24425 10626
rect 24449 10574 24495 10626
rect 24495 10574 24505 10626
rect 24529 10574 24559 10626
rect 24559 10574 24585 10626
rect 24289 10572 24345 10574
rect 24369 10572 24425 10574
rect 24449 10572 24505 10574
rect 24529 10572 24585 10574
rect 24122 10504 24178 10560
rect 24030 3160 24086 3216
rect 23754 2072 23810 2128
rect 25226 10132 25228 10152
rect 25228 10132 25280 10152
rect 25280 10132 25282 10152
rect 25226 10096 25282 10132
rect 24674 9552 24730 9608
rect 25226 9552 25282 9608
rect 24289 9538 24345 9540
rect 24369 9538 24425 9540
rect 24449 9538 24505 9540
rect 24529 9538 24585 9540
rect 24289 9486 24315 9538
rect 24315 9486 24345 9538
rect 24369 9486 24379 9538
rect 24379 9486 24425 9538
rect 24449 9486 24495 9538
rect 24495 9486 24505 9538
rect 24529 9486 24559 9538
rect 24559 9486 24585 9538
rect 24289 9484 24345 9486
rect 24369 9484 24425 9486
rect 24449 9484 24505 9486
rect 24529 9484 24585 9486
rect 24766 9316 24768 9336
rect 24768 9316 24820 9336
rect 24820 9316 24822 9336
rect 24766 9280 24822 9316
rect 24766 9008 24822 9064
rect 24490 8872 24546 8928
rect 24289 8450 24345 8452
rect 24369 8450 24425 8452
rect 24449 8450 24505 8452
rect 24529 8450 24585 8452
rect 24289 8398 24315 8450
rect 24315 8398 24345 8450
rect 24369 8398 24379 8450
rect 24379 8398 24425 8450
rect 24449 8398 24495 8450
rect 24495 8398 24505 8450
rect 24529 8398 24559 8450
rect 24559 8398 24585 8450
rect 24289 8396 24345 8398
rect 24369 8396 24425 8398
rect 24449 8396 24505 8398
rect 24529 8396 24585 8398
rect 24674 8348 24730 8384
rect 24674 8328 24676 8348
rect 24676 8328 24728 8348
rect 24728 8328 24730 8348
rect 24582 7668 24638 7704
rect 24582 7648 24584 7668
rect 24584 7648 24636 7668
rect 24636 7648 24638 7668
rect 24289 7362 24345 7364
rect 24369 7362 24425 7364
rect 24449 7362 24505 7364
rect 24529 7362 24585 7364
rect 24289 7310 24315 7362
rect 24315 7310 24345 7362
rect 24369 7310 24379 7362
rect 24379 7310 24425 7362
rect 24449 7310 24495 7362
rect 24495 7310 24505 7362
rect 24529 7310 24559 7362
rect 24559 7310 24585 7362
rect 24289 7308 24345 7310
rect 24369 7308 24425 7310
rect 24449 7308 24505 7310
rect 24529 7308 24585 7310
rect 24766 7532 24822 7568
rect 24766 7512 24768 7532
rect 24768 7512 24820 7532
rect 24820 7512 24822 7532
rect 24289 6274 24345 6276
rect 24369 6274 24425 6276
rect 24449 6274 24505 6276
rect 24529 6274 24585 6276
rect 24289 6222 24315 6274
rect 24315 6222 24345 6274
rect 24369 6222 24379 6274
rect 24379 6222 24425 6274
rect 24449 6222 24495 6274
rect 24495 6222 24505 6274
rect 24529 6222 24559 6274
rect 24559 6222 24585 6274
rect 24289 6220 24345 6222
rect 24369 6220 24425 6222
rect 24449 6220 24505 6222
rect 24529 6220 24585 6222
rect 24674 6016 24730 6072
rect 24289 5186 24345 5188
rect 24369 5186 24425 5188
rect 24449 5186 24505 5188
rect 24529 5186 24585 5188
rect 24289 5134 24315 5186
rect 24315 5134 24345 5186
rect 24369 5134 24379 5186
rect 24379 5134 24425 5186
rect 24449 5134 24495 5186
rect 24495 5134 24505 5186
rect 24529 5134 24559 5186
rect 24559 5134 24585 5186
rect 24289 5132 24345 5134
rect 24369 5132 24425 5134
rect 24449 5132 24505 5134
rect 24529 5132 24585 5134
rect 24674 4112 24730 4168
rect 24289 4098 24345 4100
rect 24369 4098 24425 4100
rect 24449 4098 24505 4100
rect 24529 4098 24585 4100
rect 24289 4046 24315 4098
rect 24315 4046 24345 4098
rect 24369 4046 24379 4098
rect 24379 4046 24425 4098
rect 24449 4046 24495 4098
rect 24495 4046 24505 4098
rect 24529 4046 24559 4098
rect 24559 4046 24585 4098
rect 24289 4044 24345 4046
rect 24369 4044 24425 4046
rect 24449 4044 24505 4046
rect 24529 4044 24585 4046
rect 26882 20160 26938 20216
rect 24766 3704 24822 3760
rect 26238 3704 26294 3760
rect 25226 3604 25228 3624
rect 25228 3604 25280 3624
rect 25280 3604 25282 3624
rect 25226 3568 25282 3604
rect 24289 3010 24345 3012
rect 24369 3010 24425 3012
rect 24449 3010 24505 3012
rect 24529 3010 24585 3012
rect 24289 2958 24315 3010
rect 24315 2958 24345 3010
rect 24369 2958 24379 3010
rect 24379 2958 24425 3010
rect 24449 2958 24495 3010
rect 24495 2958 24505 3010
rect 24529 2958 24559 3010
rect 24559 2958 24585 3010
rect 24289 2956 24345 2958
rect 24369 2956 24425 2958
rect 24449 2956 24505 2958
rect 24529 2956 24585 2958
rect 24289 1922 24345 1924
rect 24369 1922 24425 1924
rect 24449 1922 24505 1924
rect 24529 1922 24585 1924
rect 24289 1870 24315 1922
rect 24315 1870 24345 1922
rect 24369 1870 24379 1922
rect 24379 1870 24425 1922
rect 24449 1870 24495 1922
rect 24495 1870 24505 1922
rect 24529 1870 24559 1922
rect 24559 1870 24585 1922
rect 24289 1868 24345 1870
rect 24369 1868 24425 1870
rect 24449 1868 24505 1870
rect 24529 1868 24585 1870
rect 24122 1120 24178 1176
rect 23662 576 23718 632
rect 23570 32 23626 88
<< metal3 >>
rect 23197 27426 23263 27429
rect 27520 27426 28000 27456
rect 23197 27424 28000 27426
rect 23197 27368 23202 27424
rect 23258 27368 28000 27424
rect 23197 27366 28000 27368
rect 23197 27363 23263 27366
rect 27520 27336 28000 27366
rect 23565 26882 23631 26885
rect 27520 26882 28000 26912
rect 23565 26880 28000 26882
rect 23565 26824 23570 26880
rect 23626 26824 28000 26880
rect 23565 26822 28000 26824
rect 23565 26819 23631 26822
rect 27520 26792 28000 26822
rect 23381 26202 23447 26205
rect 27520 26202 28000 26232
rect 23381 26200 28000 26202
rect 23381 26144 23386 26200
rect 23442 26144 28000 26200
rect 23381 26142 28000 26144
rect 23381 26139 23447 26142
rect 27520 26112 28000 26142
rect 23289 25658 23355 25661
rect 27520 25658 28000 25688
rect 23289 25656 28000 25658
rect 23289 25600 23294 25656
rect 23350 25600 28000 25656
rect 23289 25598 28000 25600
rect 23289 25595 23355 25598
rect 27520 25568 28000 25598
rect 10277 25320 10597 25321
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 25255 10597 25256
rect 19610 25320 19930 25321
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 25255 19930 25256
rect 24761 25114 24827 25117
rect 27520 25114 28000 25144
rect 24761 25112 28000 25114
rect 24761 25056 24766 25112
rect 24822 25056 28000 25112
rect 24761 25054 28000 25056
rect 24761 25051 24827 25054
rect 27520 25024 28000 25054
rect 5610 24776 5930 24777
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5930 24776
rect 5610 24711 5930 24712
rect 14944 24776 15264 24777
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 24711 15264 24712
rect 24277 24776 24597 24777
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 24711 24597 24712
rect 13169 24570 13235 24573
rect 22829 24570 22895 24573
rect 13169 24568 22895 24570
rect 13169 24512 13174 24568
rect 13230 24512 22834 24568
rect 22890 24512 22895 24568
rect 13169 24510 22895 24512
rect 13169 24507 13235 24510
rect 22829 24507 22895 24510
rect 12525 24434 12591 24437
rect 22553 24434 22619 24437
rect 12525 24432 22619 24434
rect 12525 24376 12530 24432
rect 12586 24376 22558 24432
rect 22614 24376 22619 24432
rect 12525 24374 22619 24376
rect 12525 24371 12591 24374
rect 22553 24371 22619 24374
rect 25129 24434 25195 24437
rect 27520 24434 28000 24464
rect 25129 24432 28000 24434
rect 25129 24376 25134 24432
rect 25190 24376 28000 24432
rect 25129 24374 28000 24376
rect 25129 24371 25195 24374
rect 27520 24344 28000 24374
rect 10277 24232 10597 24233
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 10277 24167 10597 24168
rect 19610 24232 19930 24233
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 24167 19930 24168
rect 10685 24162 10751 24165
rect 18413 24162 18479 24165
rect 10685 24160 18479 24162
rect 10685 24104 10690 24160
rect 10746 24104 18418 24160
rect 18474 24104 18479 24160
rect 10685 24102 18479 24104
rect 10685 24099 10751 24102
rect 18413 24099 18479 24102
rect 9765 24026 9831 24029
rect 16113 24026 16179 24029
rect 9765 24024 16179 24026
rect 9765 23968 9770 24024
rect 9826 23968 16118 24024
rect 16174 23968 16179 24024
rect 9765 23966 16179 23968
rect 9765 23963 9831 23966
rect 16113 23963 16179 23966
rect 15101 23890 15167 23893
rect 19977 23890 20043 23893
rect 15101 23888 20043 23890
rect 15101 23832 15106 23888
rect 15162 23832 19982 23888
rect 20038 23832 20043 23888
rect 15101 23830 20043 23832
rect 15101 23827 15167 23830
rect 19977 23827 20043 23830
rect 25129 23890 25195 23893
rect 27520 23890 28000 23920
rect 25129 23888 28000 23890
rect 25129 23832 25134 23888
rect 25190 23832 28000 23888
rect 25129 23830 28000 23832
rect 25129 23827 25195 23830
rect 27520 23800 28000 23830
rect 5610 23688 5930 23689
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5930 23688
rect 5610 23623 5930 23624
rect 14944 23688 15264 23689
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 14944 23623 15264 23624
rect 24277 23688 24597 23689
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 23623 24597 23624
rect 11145 23618 11211 23621
rect 13445 23618 13511 23621
rect 11145 23616 13511 23618
rect 11145 23560 11150 23616
rect 11206 23560 13450 23616
rect 13506 23560 13511 23616
rect 11145 23558 13511 23560
rect 11145 23555 11211 23558
rect 13445 23555 13511 23558
rect 18137 23618 18203 23621
rect 18781 23618 18847 23621
rect 22093 23618 22159 23621
rect 18137 23616 22159 23618
rect 18137 23560 18142 23616
rect 18198 23560 18786 23616
rect 18842 23560 22098 23616
rect 22154 23560 22159 23616
rect 18137 23558 22159 23560
rect 18137 23555 18203 23558
rect 18781 23555 18847 23558
rect 22093 23555 22159 23558
rect 4337 23346 4403 23349
rect 22369 23346 22435 23349
rect 25497 23346 25563 23349
rect 4337 23344 22435 23346
rect 4337 23288 4342 23344
rect 4398 23288 22374 23344
rect 22430 23288 22435 23344
rect 4337 23286 22435 23288
rect 4337 23283 4403 23286
rect 22369 23283 22435 23286
rect 23982 23344 25563 23346
rect 23982 23288 25502 23344
rect 25558 23288 25563 23344
rect 23982 23286 25563 23288
rect 10277 23144 10597 23145
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 23079 10597 23080
rect 19610 23144 19930 23145
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 19610 23079 19930 23080
rect 12157 23074 12223 23077
rect 14825 23074 14891 23077
rect 15193 23074 15259 23077
rect 12157 23072 15259 23074
rect 12157 23016 12162 23072
rect 12218 23016 14830 23072
rect 14886 23016 15198 23072
rect 15254 23016 15259 23072
rect 12157 23014 15259 23016
rect 12157 23011 12223 23014
rect 14825 23011 14891 23014
rect 15193 23011 15259 23014
rect 3417 22802 3483 22805
rect 11237 22802 11303 22805
rect 12709 22802 12775 22805
rect 3417 22800 12775 22802
rect 3417 22744 3422 22800
rect 3478 22744 11242 22800
rect 11298 22744 12714 22800
rect 12770 22744 12775 22800
rect 3417 22742 12775 22744
rect 3417 22739 3483 22742
rect 11237 22739 11303 22742
rect 12709 22739 12775 22742
rect 13721 22802 13787 22805
rect 16389 22802 16455 22805
rect 23841 22802 23907 22805
rect 13721 22800 16314 22802
rect 13721 22744 13726 22800
rect 13782 22744 16314 22800
rect 13721 22742 16314 22744
rect 13721 22739 13787 22742
rect 16254 22666 16314 22742
rect 16389 22800 23907 22802
rect 16389 22744 16394 22800
rect 16450 22744 23846 22800
rect 23902 22744 23907 22800
rect 16389 22742 23907 22744
rect 16389 22739 16455 22742
rect 23841 22739 23907 22742
rect 22277 22666 22343 22669
rect 16254 22664 22343 22666
rect 16254 22608 22282 22664
rect 22338 22608 22343 22664
rect 16254 22606 22343 22608
rect 22277 22603 22343 22606
rect 23841 22666 23907 22669
rect 23982 22666 24042 23286
rect 25497 23283 25563 23286
rect 27520 23210 28000 23240
rect 25454 23150 28000 23210
rect 25454 23077 25514 23150
rect 27520 23120 28000 23150
rect 25405 23072 25514 23077
rect 25405 23016 25410 23072
rect 25466 23016 25514 23072
rect 25405 23014 25514 23016
rect 25405 23011 25471 23014
rect 23841 22664 24042 22666
rect 23841 22608 23846 22664
rect 23902 22608 24042 22664
rect 23841 22606 24042 22608
rect 24669 22666 24735 22669
rect 27520 22666 28000 22696
rect 24669 22664 28000 22666
rect 24669 22608 24674 22664
rect 24730 22608 28000 22664
rect 24669 22606 28000 22608
rect 23841 22603 23907 22606
rect 24669 22603 24735 22606
rect 5610 22600 5930 22601
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5930 22600
rect 5610 22535 5930 22536
rect 14944 22600 15264 22601
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 22535 15264 22536
rect 24277 22600 24597 22601
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 27520 22576 28000 22606
rect 24277 22535 24597 22536
rect 18137 22530 18203 22533
rect 20989 22530 21055 22533
rect 18137 22528 21055 22530
rect 18137 22472 18142 22528
rect 18198 22472 20994 22528
rect 21050 22472 21055 22528
rect 18137 22470 21055 22472
rect 18137 22467 18203 22470
rect 20989 22467 21055 22470
rect 21357 22530 21423 22533
rect 23933 22530 23999 22533
rect 21357 22528 23999 22530
rect 21357 22472 21362 22528
rect 21418 22472 23938 22528
rect 23994 22472 23999 22528
rect 21357 22470 23999 22472
rect 21357 22467 21423 22470
rect 23933 22467 23999 22470
rect 7741 22394 7807 22397
rect 24761 22394 24827 22397
rect 7741 22392 24827 22394
rect 7741 22336 7746 22392
rect 7802 22336 24766 22392
rect 24822 22336 24827 22392
rect 7741 22334 24827 22336
rect 7741 22331 7807 22334
rect 24761 22331 24827 22334
rect 4981 22258 5047 22261
rect 20713 22258 20779 22261
rect 4981 22256 20779 22258
rect 4981 22200 4986 22256
rect 5042 22200 20718 22256
rect 20774 22200 20779 22256
rect 4981 22198 20779 22200
rect 4981 22195 5047 22198
rect 20713 22195 20779 22198
rect 13721 22122 13787 22125
rect 13997 22122 14063 22125
rect 18413 22122 18479 22125
rect 13721 22120 18479 22122
rect 13721 22064 13726 22120
rect 13782 22064 14002 22120
rect 14058 22064 18418 22120
rect 18474 22064 18479 22120
rect 13721 22062 18479 22064
rect 13721 22059 13787 22062
rect 13997 22059 14063 22062
rect 18413 22059 18479 22062
rect 24945 22122 25011 22125
rect 27520 22122 28000 22152
rect 24945 22120 28000 22122
rect 24945 22064 24950 22120
rect 25006 22064 28000 22120
rect 24945 22062 28000 22064
rect 24945 22059 25011 22062
rect 10277 22056 10597 22057
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 10277 21991 10597 21992
rect 19610 22056 19930 22057
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 27520 22032 28000 22062
rect 19610 21991 19930 21992
rect 18321 21850 18387 21853
rect 25681 21850 25747 21853
rect 18321 21848 25747 21850
rect 18321 21792 18326 21848
rect 18382 21792 25686 21848
rect 25742 21792 25747 21848
rect 18321 21790 25747 21792
rect 18321 21787 18387 21790
rect 25681 21787 25747 21790
rect 14273 21714 14339 21717
rect 18321 21714 18387 21717
rect 22921 21714 22987 21717
rect 24669 21714 24735 21717
rect 14273 21712 18200 21714
rect 14273 21656 14278 21712
rect 14334 21656 18200 21712
rect 14273 21654 18200 21656
rect 14273 21651 14339 21654
rect 6361 21578 6427 21581
rect 11513 21578 11579 21581
rect 6361 21576 11579 21578
rect 6361 21520 6366 21576
rect 6422 21520 11518 21576
rect 11574 21520 11579 21576
rect 6361 21518 11579 21520
rect 18140 21578 18200 21654
rect 18321 21712 22754 21714
rect 18321 21656 18326 21712
rect 18382 21656 22754 21712
rect 18321 21654 22754 21656
rect 18321 21651 18387 21654
rect 22694 21578 22754 21654
rect 22921 21712 24735 21714
rect 22921 21656 22926 21712
rect 22982 21656 24674 21712
rect 24730 21656 24735 21712
rect 22921 21654 24735 21656
rect 22921 21651 22987 21654
rect 24669 21651 24735 21654
rect 24117 21578 24183 21581
rect 18140 21518 22570 21578
rect 22694 21576 24183 21578
rect 22694 21520 24122 21576
rect 24178 21520 24183 21576
rect 22694 21518 24183 21520
rect 6361 21515 6427 21518
rect 11513 21515 11579 21518
rect 5610 21512 5930 21513
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5930 21512
rect 5610 21447 5930 21448
rect 14944 21512 15264 21513
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 21447 15264 21448
rect 7097 21442 7163 21445
rect 22510 21442 22570 21518
rect 24117 21515 24183 21518
rect 24277 21512 24597 21513
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 24277 21447 24597 21448
rect 23657 21442 23723 21445
rect 7097 21440 14842 21442
rect 7097 21384 7102 21440
rect 7158 21384 14842 21440
rect 7097 21382 14842 21384
rect 22510 21440 23723 21442
rect 22510 21384 23662 21440
rect 23718 21384 23723 21440
rect 22510 21382 23723 21384
rect 7097 21379 7163 21382
rect 14782 21306 14842 21382
rect 23657 21379 23723 21382
rect 24761 21442 24827 21445
rect 27520 21442 28000 21472
rect 24761 21440 28000 21442
rect 24761 21384 24766 21440
rect 24822 21384 28000 21440
rect 24761 21382 28000 21384
rect 24761 21379 24827 21382
rect 27520 21352 28000 21382
rect 18321 21306 18387 21309
rect 14782 21304 18387 21306
rect 14782 21248 18326 21304
rect 18382 21248 18387 21304
rect 14782 21246 18387 21248
rect 18321 21243 18387 21246
rect 9121 21170 9187 21173
rect 13537 21170 13603 21173
rect 25129 21170 25195 21173
rect 9121 21168 13370 21170
rect 9121 21112 9126 21168
rect 9182 21112 13370 21168
rect 9121 21110 13370 21112
rect 9121 21107 9187 21110
rect 13310 21034 13370 21110
rect 13537 21168 25195 21170
rect 13537 21112 13542 21168
rect 13598 21112 25134 21168
rect 25190 21112 25195 21168
rect 13537 21110 25195 21112
rect 13537 21107 13603 21110
rect 25129 21107 25195 21110
rect 15837 21034 15903 21037
rect 13310 21032 15903 21034
rect 13310 20976 15842 21032
rect 15898 20976 15903 21032
rect 13310 20974 15903 20976
rect 15837 20971 15903 20974
rect 10277 20968 10597 20969
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 20903 10597 20904
rect 19610 20968 19930 20969
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 20903 19930 20904
rect 14641 20898 14707 20901
rect 17033 20898 17099 20901
rect 14641 20896 17099 20898
rect 14641 20840 14646 20896
rect 14702 20840 17038 20896
rect 17094 20840 17099 20896
rect 14641 20838 17099 20840
rect 14641 20835 14707 20838
rect 17033 20835 17099 20838
rect 25313 20898 25379 20901
rect 27520 20898 28000 20928
rect 25313 20896 28000 20898
rect 25313 20840 25318 20896
rect 25374 20840 28000 20896
rect 25313 20838 28000 20840
rect 25313 20835 25379 20838
rect 27520 20808 28000 20838
rect 0 20762 480 20792
rect 3417 20762 3483 20765
rect 0 20760 3483 20762
rect 0 20704 3422 20760
rect 3478 20704 3483 20760
rect 0 20702 3483 20704
rect 0 20672 480 20702
rect 3417 20699 3483 20702
rect 5993 20762 6059 20765
rect 17953 20762 18019 20765
rect 5993 20760 18019 20762
rect 5993 20704 5998 20760
rect 6054 20704 17958 20760
rect 18014 20704 18019 20760
rect 5993 20702 18019 20704
rect 5993 20699 6059 20702
rect 17953 20699 18019 20702
rect 20897 20762 20963 20765
rect 23841 20762 23907 20765
rect 20897 20760 23907 20762
rect 20897 20704 20902 20760
rect 20958 20704 23846 20760
rect 23902 20704 23907 20760
rect 20897 20702 23907 20704
rect 20897 20699 20963 20702
rect 23841 20699 23907 20702
rect 15561 20626 15627 20629
rect 23657 20626 23723 20629
rect 15561 20624 23723 20626
rect 15561 20568 15566 20624
rect 15622 20568 23662 20624
rect 23718 20568 23723 20624
rect 15561 20566 23723 20568
rect 15561 20563 15627 20566
rect 23657 20563 23723 20566
rect 13537 20490 13603 20493
rect 14549 20490 14615 20493
rect 13537 20488 14615 20490
rect 13537 20432 13542 20488
rect 13598 20432 14554 20488
rect 14610 20432 14615 20488
rect 13537 20430 14615 20432
rect 13537 20427 13603 20430
rect 14549 20427 14615 20430
rect 5610 20424 5930 20425
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5930 20424
rect 5610 20359 5930 20360
rect 14944 20424 15264 20425
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 14944 20359 15264 20360
rect 24277 20424 24597 20425
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 24277 20359 24597 20360
rect 25129 20354 25195 20357
rect 27520 20354 28000 20384
rect 25129 20352 28000 20354
rect 25129 20296 25134 20352
rect 25190 20296 28000 20352
rect 25129 20294 28000 20296
rect 25129 20291 25195 20294
rect 27520 20264 28000 20294
rect 25589 20218 25655 20221
rect 26877 20218 26943 20221
rect 25589 20216 26943 20218
rect 25589 20160 25594 20216
rect 25650 20160 26882 20216
rect 26938 20160 26943 20216
rect 25589 20158 26943 20160
rect 25589 20155 25655 20158
rect 26877 20155 26943 20158
rect 10869 20082 10935 20085
rect 17585 20082 17651 20085
rect 10869 20080 17651 20082
rect 10869 20024 10874 20080
rect 10930 20024 17590 20080
rect 17646 20024 17651 20080
rect 10869 20022 17651 20024
rect 10869 20019 10935 20022
rect 17585 20019 17651 20022
rect 10277 19880 10597 19881
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 19815 10597 19816
rect 19610 19880 19930 19881
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 19815 19930 19816
rect 18965 19674 19031 19677
rect 24945 19674 25011 19677
rect 18965 19672 25011 19674
rect 18965 19616 18970 19672
rect 19026 19616 24950 19672
rect 25006 19616 25011 19672
rect 18965 19614 25011 19616
rect 18965 19611 19031 19614
rect 24945 19611 25011 19614
rect 25405 19674 25471 19677
rect 27520 19674 28000 19704
rect 25405 19672 28000 19674
rect 25405 19616 25410 19672
rect 25466 19616 28000 19672
rect 25405 19614 28000 19616
rect 25405 19611 25471 19614
rect 27520 19584 28000 19614
rect 5610 19336 5930 19337
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5930 19336
rect 5610 19271 5930 19272
rect 14944 19336 15264 19337
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 19271 15264 19272
rect 24277 19336 24597 19337
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 24277 19271 24597 19272
rect 16389 19266 16455 19269
rect 16849 19266 16915 19269
rect 21541 19266 21607 19269
rect 16389 19264 21607 19266
rect 16389 19208 16394 19264
rect 16450 19208 16854 19264
rect 16910 19208 21546 19264
rect 21602 19208 21607 19264
rect 16389 19206 21607 19208
rect 16389 19203 16455 19206
rect 16849 19203 16915 19206
rect 21541 19203 21607 19206
rect 3693 19130 3759 19133
rect 22093 19130 22159 19133
rect 3693 19128 22159 19130
rect 3693 19072 3698 19128
rect 3754 19072 22098 19128
rect 22154 19072 22159 19128
rect 3693 19070 22159 19072
rect 3693 19067 3759 19070
rect 22093 19067 22159 19070
rect 25129 19130 25195 19133
rect 27520 19130 28000 19160
rect 25129 19128 28000 19130
rect 25129 19072 25134 19128
rect 25190 19072 28000 19128
rect 25129 19070 28000 19072
rect 25129 19067 25195 19070
rect 27520 19040 28000 19070
rect 8385 18994 8451 18997
rect 13445 18994 13511 18997
rect 8385 18992 13511 18994
rect 8385 18936 8390 18992
rect 8446 18936 13450 18992
rect 13506 18936 13511 18992
rect 8385 18934 13511 18936
rect 8385 18931 8451 18934
rect 13445 18931 13511 18934
rect 13629 18858 13695 18861
rect 15745 18858 15811 18861
rect 13629 18856 15811 18858
rect 13629 18800 13634 18856
rect 13690 18800 15750 18856
rect 15806 18800 15811 18856
rect 13629 18798 15811 18800
rect 13629 18795 13695 18798
rect 15745 18795 15811 18798
rect 21633 18858 21699 18861
rect 23289 18858 23355 18861
rect 21633 18856 23355 18858
rect 21633 18800 21638 18856
rect 21694 18800 23294 18856
rect 23350 18800 23355 18856
rect 21633 18798 23355 18800
rect 21633 18795 21699 18798
rect 23289 18795 23355 18798
rect 10277 18792 10597 18793
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 18727 10597 18728
rect 19610 18792 19930 18793
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 19610 18727 19930 18728
rect 2957 18450 3023 18453
rect 20713 18450 20779 18453
rect 2957 18448 20779 18450
rect 2957 18392 2962 18448
rect 3018 18392 20718 18448
rect 20774 18392 20779 18448
rect 2957 18390 20779 18392
rect 2957 18387 3023 18390
rect 20713 18387 20779 18390
rect 25313 18450 25379 18453
rect 27520 18450 28000 18480
rect 25313 18448 28000 18450
rect 25313 18392 25318 18448
rect 25374 18392 28000 18448
rect 25313 18390 28000 18392
rect 25313 18387 25379 18390
rect 27520 18360 28000 18390
rect 5610 18248 5930 18249
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5930 18248
rect 5610 18183 5930 18184
rect 14944 18248 15264 18249
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 18183 15264 18184
rect 24277 18248 24597 18249
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 24277 18183 24597 18184
rect 15377 18178 15443 18181
rect 23749 18178 23815 18181
rect 15377 18176 23815 18178
rect 15377 18120 15382 18176
rect 15438 18120 23754 18176
rect 23810 18120 23815 18176
rect 15377 18118 23815 18120
rect 15377 18115 15443 18118
rect 23749 18115 23815 18118
rect 2313 17906 2379 17909
rect 16389 17906 16455 17909
rect 2313 17904 16455 17906
rect 2313 17848 2318 17904
rect 2374 17848 16394 17904
rect 16450 17848 16455 17904
rect 2313 17846 16455 17848
rect 2313 17843 2379 17846
rect 16389 17843 16455 17846
rect 24761 17906 24827 17909
rect 27520 17906 28000 17936
rect 24761 17904 28000 17906
rect 24761 17848 24766 17904
rect 24822 17848 28000 17904
rect 24761 17846 28000 17848
rect 24761 17843 24827 17846
rect 27520 17816 28000 17846
rect 21817 17770 21883 17773
rect 23657 17770 23723 17773
rect 21817 17768 23723 17770
rect 21817 17712 21822 17768
rect 21878 17712 23662 17768
rect 23718 17712 23723 17768
rect 21817 17710 23723 17712
rect 21817 17707 21883 17710
rect 23657 17707 23723 17710
rect 10277 17704 10597 17705
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 17639 10597 17640
rect 19610 17704 19930 17705
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 19610 17639 19930 17640
rect 16481 17634 16547 17637
rect 18505 17634 18571 17637
rect 16481 17632 18571 17634
rect 16481 17576 16486 17632
rect 16542 17576 18510 17632
rect 18566 17576 18571 17632
rect 16481 17574 18571 17576
rect 16481 17571 16547 17574
rect 18505 17571 18571 17574
rect 18413 17498 18479 17501
rect 21725 17498 21791 17501
rect 18413 17496 21791 17498
rect 18413 17440 18418 17496
rect 18474 17440 21730 17496
rect 21786 17440 21791 17496
rect 18413 17438 21791 17440
rect 18413 17435 18479 17438
rect 21725 17435 21791 17438
rect 933 17362 999 17365
rect 21173 17362 21239 17365
rect 933 17360 21239 17362
rect 933 17304 938 17360
rect 994 17304 21178 17360
rect 21234 17304 21239 17360
rect 933 17302 21239 17304
rect 933 17299 999 17302
rect 21173 17299 21239 17302
rect 25405 17362 25471 17365
rect 27520 17362 28000 17392
rect 25405 17360 28000 17362
rect 25405 17304 25410 17360
rect 25466 17304 28000 17360
rect 25405 17302 28000 17304
rect 25405 17299 25471 17302
rect 27520 17272 28000 17302
rect 5610 17160 5930 17161
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5930 17160
rect 5610 17095 5930 17096
rect 14944 17160 15264 17161
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 17095 15264 17096
rect 24277 17160 24597 17161
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 24277 17095 24597 17096
rect 11789 16954 11855 16957
rect 18413 16954 18479 16957
rect 11789 16952 18479 16954
rect 11789 16896 11794 16952
rect 11850 16896 18418 16952
rect 18474 16896 18479 16952
rect 11789 16894 18479 16896
rect 11789 16891 11855 16894
rect 18413 16891 18479 16894
rect 1577 16818 1643 16821
rect 14181 16818 14247 16821
rect 1577 16816 14247 16818
rect 1577 16760 1582 16816
rect 1638 16760 14186 16816
rect 14242 16760 14247 16816
rect 1577 16758 14247 16760
rect 1577 16755 1643 16758
rect 14181 16755 14247 16758
rect 18689 16818 18755 16821
rect 23933 16818 23999 16821
rect 18689 16816 23999 16818
rect 18689 16760 18694 16816
rect 18750 16760 23938 16816
rect 23994 16760 23999 16816
rect 18689 16758 23999 16760
rect 18689 16755 18755 16758
rect 23933 16755 23999 16758
rect 25405 16682 25471 16685
rect 27520 16682 28000 16712
rect 25405 16680 28000 16682
rect 25405 16624 25410 16680
rect 25466 16624 28000 16680
rect 25405 16622 28000 16624
rect 25405 16619 25471 16622
rect 10277 16616 10597 16617
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 16551 10597 16552
rect 19610 16616 19930 16617
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 27520 16592 28000 16622
rect 19610 16551 19930 16552
rect 21909 16546 21975 16549
rect 24025 16546 24091 16549
rect 21909 16544 24091 16546
rect 21909 16488 21914 16544
rect 21970 16488 24030 16544
rect 24086 16488 24091 16544
rect 21909 16486 24091 16488
rect 21909 16483 21975 16486
rect 24025 16483 24091 16486
rect 19057 16410 19123 16413
rect 22185 16410 22251 16413
rect 19057 16408 22251 16410
rect 19057 16352 19062 16408
rect 19118 16352 22190 16408
rect 22246 16352 22251 16408
rect 19057 16350 22251 16352
rect 19057 16347 19123 16350
rect 22185 16347 22251 16350
rect 24761 16138 24827 16141
rect 27520 16138 28000 16168
rect 24761 16136 28000 16138
rect 24761 16080 24766 16136
rect 24822 16080 28000 16136
rect 24761 16078 28000 16080
rect 24761 16075 24827 16078
rect 5610 16072 5930 16073
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5930 16072
rect 5610 16007 5930 16008
rect 14944 16072 15264 16073
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 16007 15264 16008
rect 24277 16072 24597 16073
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 27520 16048 28000 16078
rect 24277 16007 24597 16008
rect 18689 15730 18755 15733
rect 18416 15728 18755 15730
rect 18416 15672 18694 15728
rect 18750 15672 18755 15728
rect 18416 15670 18755 15672
rect 18416 15597 18476 15670
rect 18689 15667 18755 15670
rect 15653 15594 15719 15597
rect 18413 15594 18479 15597
rect 15653 15592 18479 15594
rect 15653 15536 15658 15592
rect 15714 15536 18418 15592
rect 18474 15536 18479 15592
rect 15653 15534 18479 15536
rect 15653 15531 15719 15534
rect 18413 15531 18479 15534
rect 10277 15528 10597 15529
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 15463 10597 15464
rect 19610 15528 19930 15529
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 15463 19930 15464
rect 13905 15458 13971 15461
rect 16389 15458 16455 15461
rect 13905 15456 16455 15458
rect 13905 15400 13910 15456
rect 13966 15400 16394 15456
rect 16450 15400 16455 15456
rect 13905 15398 16455 15400
rect 13905 15395 13971 15398
rect 16389 15395 16455 15398
rect 25497 15458 25563 15461
rect 27520 15458 28000 15488
rect 25497 15456 28000 15458
rect 25497 15400 25502 15456
rect 25558 15400 28000 15456
rect 25497 15398 28000 15400
rect 25497 15395 25563 15398
rect 27520 15368 28000 15398
rect 13905 15322 13971 15325
rect 23657 15322 23723 15325
rect 13905 15320 23723 15322
rect 13905 15264 13910 15320
rect 13966 15264 23662 15320
rect 23718 15264 23723 15320
rect 13905 15262 23723 15264
rect 13905 15259 13971 15262
rect 23657 15259 23723 15262
rect 16297 15050 16363 15053
rect 21357 15050 21423 15053
rect 23381 15050 23447 15053
rect 16297 15048 23447 15050
rect 16297 14992 16302 15048
rect 16358 14992 21362 15048
rect 21418 14992 23386 15048
rect 23442 14992 23447 15048
rect 16297 14990 23447 14992
rect 16297 14987 16363 14990
rect 21357 14987 21423 14990
rect 23381 14987 23447 14990
rect 5610 14984 5930 14985
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5930 14984
rect 5610 14919 5930 14920
rect 14944 14984 15264 14985
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 14919 15264 14920
rect 24277 14984 24597 14985
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 14919 24597 14920
rect 25865 14914 25931 14917
rect 27520 14914 28000 14944
rect 25865 14912 28000 14914
rect 25865 14856 25870 14912
rect 25926 14856 28000 14912
rect 25865 14854 28000 14856
rect 25865 14851 25931 14854
rect 27520 14824 28000 14854
rect 15929 14778 15995 14781
rect 19057 14778 19123 14781
rect 20713 14778 20779 14781
rect 15929 14776 20779 14778
rect 15929 14720 15934 14776
rect 15990 14720 19062 14776
rect 19118 14720 20718 14776
rect 20774 14720 20779 14776
rect 15929 14718 20779 14720
rect 15929 14715 15995 14718
rect 19057 14715 19123 14718
rect 20713 14715 20779 14718
rect 10277 14440 10597 14441
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 14375 10597 14376
rect 19610 14440 19930 14441
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 14375 19930 14376
rect 25589 14370 25655 14373
rect 27520 14370 28000 14400
rect 25589 14368 28000 14370
rect 25589 14312 25594 14368
rect 25650 14312 28000 14368
rect 25589 14310 28000 14312
rect 25589 14307 25655 14310
rect 27520 14280 28000 14310
rect 18689 14234 18755 14237
rect 23657 14234 23723 14237
rect 18689 14232 23723 14234
rect 18689 14176 18694 14232
rect 18750 14176 23662 14232
rect 23718 14176 23723 14232
rect 18689 14174 23723 14176
rect 18689 14171 18755 14174
rect 23657 14171 23723 14174
rect 5610 13896 5930 13897
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5930 13896
rect 5610 13831 5930 13832
rect 14944 13896 15264 13897
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 13831 15264 13832
rect 24277 13896 24597 13897
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 13831 24597 13832
rect 16389 13826 16455 13829
rect 20253 13826 20319 13829
rect 16389 13824 20319 13826
rect 16389 13768 16394 13824
rect 16450 13768 20258 13824
rect 20314 13768 20319 13824
rect 16389 13766 20319 13768
rect 16389 13763 16455 13766
rect 20253 13763 20319 13766
rect 18873 13690 18939 13693
rect 20897 13690 20963 13693
rect 18873 13688 20963 13690
rect 18873 13632 18878 13688
rect 18934 13632 20902 13688
rect 20958 13632 20963 13688
rect 18873 13630 20963 13632
rect 18873 13627 18939 13630
rect 20897 13627 20963 13630
rect 25221 13690 25287 13693
rect 27520 13690 28000 13720
rect 25221 13688 28000 13690
rect 25221 13632 25226 13688
rect 25282 13632 28000 13688
rect 25221 13630 28000 13632
rect 25221 13627 25287 13630
rect 27520 13600 28000 13630
rect 10277 13352 10597 13353
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 13287 10597 13288
rect 19610 13352 19930 13353
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 13287 19930 13288
rect 19241 13146 19307 13149
rect 23933 13146 23999 13149
rect 19241 13144 23999 13146
rect 19241 13088 19246 13144
rect 19302 13088 23938 13144
rect 23994 13088 23999 13144
rect 19241 13086 23999 13088
rect 19241 13083 19307 13086
rect 23933 13083 23999 13086
rect 25037 13146 25103 13149
rect 27520 13146 28000 13176
rect 25037 13144 28000 13146
rect 25037 13088 25042 13144
rect 25098 13088 28000 13144
rect 25037 13086 28000 13088
rect 25037 13083 25103 13086
rect 27520 13056 28000 13086
rect 5610 12808 5930 12809
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5930 12808
rect 5610 12743 5930 12744
rect 14944 12808 15264 12809
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 12743 15264 12744
rect 24277 12808 24597 12809
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 12743 24597 12744
rect 24669 12602 24735 12605
rect 27520 12602 28000 12632
rect 24669 12600 28000 12602
rect 24669 12544 24674 12600
rect 24730 12544 28000 12600
rect 24669 12542 28000 12544
rect 24669 12539 24735 12542
rect 27520 12512 28000 12542
rect 10277 12264 10597 12265
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 12199 10597 12200
rect 19610 12264 19930 12265
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 12199 19930 12200
rect 24577 11922 24643 11925
rect 27520 11922 28000 11952
rect 24577 11920 28000 11922
rect 24577 11864 24582 11920
rect 24638 11864 28000 11920
rect 24577 11862 28000 11864
rect 24577 11859 24643 11862
rect 27520 11832 28000 11862
rect 5610 11720 5930 11721
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5930 11720
rect 5610 11655 5930 11656
rect 14944 11720 15264 11721
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 11655 15264 11656
rect 24277 11720 24597 11721
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 11655 24597 11656
rect 19241 11514 19307 11517
rect 21449 11514 21515 11517
rect 19241 11512 21515 11514
rect 19241 11456 19246 11512
rect 19302 11456 21454 11512
rect 21510 11456 21515 11512
rect 19241 11454 21515 11456
rect 19241 11451 19307 11454
rect 21449 11451 21515 11454
rect 3417 11378 3483 11381
rect 10133 11378 10199 11381
rect 3417 11376 10199 11378
rect 3417 11320 3422 11376
rect 3478 11320 10138 11376
rect 10194 11320 10199 11376
rect 3417 11318 10199 11320
rect 3417 11315 3483 11318
rect 10133 11315 10199 11318
rect 21173 11378 21239 11381
rect 27520 11378 28000 11408
rect 21173 11376 28000 11378
rect 21173 11320 21178 11376
rect 21234 11320 28000 11376
rect 21173 11318 28000 11320
rect 21173 11315 21239 11318
rect 27520 11288 28000 11318
rect 10277 11176 10597 11177
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 11111 10597 11112
rect 19610 11176 19930 11177
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 11111 19930 11112
rect 473 10970 539 10973
rect 13537 10970 13603 10973
rect 473 10968 13603 10970
rect 473 10912 478 10968
rect 534 10912 13542 10968
rect 13598 10912 13603 10968
rect 473 10910 13603 10912
rect 473 10907 539 10910
rect 13537 10907 13603 10910
rect 22921 10698 22987 10701
rect 24025 10698 24091 10701
rect 22921 10696 24091 10698
rect 22921 10640 22926 10696
rect 22982 10640 24030 10696
rect 24086 10640 24091 10696
rect 22921 10638 24091 10640
rect 22921 10635 22987 10638
rect 24025 10635 24091 10638
rect 24669 10698 24735 10701
rect 27520 10698 28000 10728
rect 24669 10696 28000 10698
rect 24669 10640 24674 10696
rect 24730 10640 28000 10696
rect 24669 10638 28000 10640
rect 24669 10635 24735 10638
rect 5610 10632 5930 10633
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5930 10632
rect 5610 10567 5930 10568
rect 14944 10632 15264 10633
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 10567 15264 10568
rect 24277 10632 24597 10633
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 27520 10608 28000 10638
rect 24277 10567 24597 10568
rect 22001 10562 22067 10565
rect 24117 10562 24183 10565
rect 22001 10560 24183 10562
rect 22001 10504 22006 10560
rect 22062 10504 24122 10560
rect 24178 10504 24183 10560
rect 22001 10502 24183 10504
rect 22001 10499 22067 10502
rect 24117 10499 24183 10502
rect 25221 10154 25287 10157
rect 27520 10154 28000 10184
rect 25221 10152 28000 10154
rect 25221 10096 25226 10152
rect 25282 10096 28000 10152
rect 25221 10094 28000 10096
rect 25221 10091 25287 10094
rect 10277 10088 10597 10089
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 10023 10597 10024
rect 19610 10088 19930 10089
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 27520 10064 28000 10094
rect 19610 10023 19930 10024
rect 24669 9610 24735 9613
rect 25221 9610 25287 9613
rect 27520 9610 28000 9640
rect 24669 9608 28000 9610
rect 24669 9552 24674 9608
rect 24730 9552 25226 9608
rect 25282 9552 28000 9608
rect 24669 9550 28000 9552
rect 24669 9547 24735 9550
rect 25221 9547 25287 9550
rect 5610 9544 5930 9545
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5930 9544
rect 5610 9479 5930 9480
rect 14944 9544 15264 9545
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 9479 15264 9480
rect 24277 9544 24597 9545
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 27520 9520 28000 9550
rect 24277 9479 24597 9480
rect 20437 9338 20503 9341
rect 24761 9338 24827 9341
rect 20437 9336 24827 9338
rect 20437 9280 20442 9336
rect 20498 9280 24766 9336
rect 24822 9280 24827 9336
rect 20437 9278 24827 9280
rect 20437 9275 20503 9278
rect 24761 9275 24827 9278
rect 20621 9066 20687 9069
rect 24761 9066 24827 9069
rect 20621 9064 24827 9066
rect 20621 9008 20626 9064
rect 20682 9008 24766 9064
rect 24822 9008 24827 9064
rect 20621 9006 24827 9008
rect 20621 9003 20687 9006
rect 24761 9003 24827 9006
rect 10277 9000 10597 9001
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 8935 10597 8936
rect 19610 9000 19930 9001
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 8935 19930 8936
rect 24485 8930 24551 8933
rect 27520 8930 28000 8960
rect 24485 8928 28000 8930
rect 24485 8872 24490 8928
rect 24546 8872 28000 8928
rect 24485 8870 28000 8872
rect 24485 8867 24551 8870
rect 27520 8840 28000 8870
rect 5610 8456 5930 8457
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5930 8456
rect 5610 8391 5930 8392
rect 14944 8456 15264 8457
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 8391 15264 8392
rect 24277 8456 24597 8457
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 8391 24597 8392
rect 24669 8386 24735 8389
rect 27520 8386 28000 8416
rect 24669 8384 28000 8386
rect 24669 8328 24674 8384
rect 24730 8328 28000 8384
rect 24669 8326 28000 8328
rect 24669 8323 24735 8326
rect 27520 8296 28000 8326
rect 10277 7912 10597 7913
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 7847 10597 7848
rect 19610 7912 19930 7913
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 19610 7847 19930 7848
rect 15653 7706 15719 7709
rect 23657 7706 23723 7709
rect 15653 7704 23723 7706
rect 15653 7648 15658 7704
rect 15714 7648 23662 7704
rect 23718 7648 23723 7704
rect 15653 7646 23723 7648
rect 15653 7643 15719 7646
rect 23657 7643 23723 7646
rect 24577 7706 24643 7709
rect 27520 7706 28000 7736
rect 24577 7704 28000 7706
rect 24577 7648 24582 7704
rect 24638 7648 28000 7704
rect 24577 7646 28000 7648
rect 24577 7643 24643 7646
rect 27520 7616 28000 7646
rect 19149 7570 19215 7573
rect 24761 7570 24827 7573
rect 19149 7568 24827 7570
rect 19149 7512 19154 7568
rect 19210 7512 24766 7568
rect 24822 7512 24827 7568
rect 19149 7510 24827 7512
rect 19149 7507 19215 7510
rect 24761 7507 24827 7510
rect 5610 7368 5930 7369
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5930 7368
rect 5610 7303 5930 7304
rect 14944 7368 15264 7369
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 7303 15264 7304
rect 24277 7368 24597 7369
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 24277 7303 24597 7304
rect 17769 7298 17835 7301
rect 18689 7298 18755 7301
rect 17769 7296 18755 7298
rect 17769 7240 17774 7296
rect 17830 7240 18694 7296
rect 18750 7240 18755 7296
rect 17769 7238 18755 7240
rect 17769 7235 17835 7238
rect 18689 7235 18755 7238
rect 18229 7162 18295 7165
rect 27520 7162 28000 7192
rect 18229 7160 28000 7162
rect 18229 7104 18234 7160
rect 18290 7104 28000 7160
rect 18229 7102 28000 7104
rect 18229 7099 18295 7102
rect 27520 7072 28000 7102
rect 10277 6824 10597 6825
rect 0 6754 480 6784
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 6759 10597 6760
rect 19610 6824 19930 6825
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 19610 6759 19930 6760
rect 3417 6754 3483 6757
rect 0 6752 3483 6754
rect 0 6696 3422 6752
rect 3478 6696 3483 6752
rect 0 6694 3483 6696
rect 0 6664 480 6694
rect 3417 6691 3483 6694
rect 23473 6618 23539 6621
rect 27520 6618 28000 6648
rect 23473 6616 28000 6618
rect 23473 6560 23478 6616
rect 23534 6560 28000 6616
rect 23473 6558 28000 6560
rect 23473 6555 23539 6558
rect 27520 6528 28000 6558
rect 5610 6280 5930 6281
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5930 6280
rect 5610 6215 5930 6216
rect 14944 6280 15264 6281
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 6215 15264 6216
rect 24277 6280 24597 6281
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 24277 6215 24597 6216
rect 13169 6074 13235 6077
rect 24669 6074 24735 6077
rect 13169 6072 24735 6074
rect 13169 6016 13174 6072
rect 13230 6016 24674 6072
rect 24730 6016 24735 6072
rect 13169 6014 24735 6016
rect 13169 6011 13235 6014
rect 24669 6011 24735 6014
rect 16849 5938 16915 5941
rect 27520 5938 28000 5968
rect 16849 5936 28000 5938
rect 16849 5880 16854 5936
rect 16910 5880 28000 5936
rect 16849 5878 28000 5880
rect 16849 5875 16915 5878
rect 27520 5848 28000 5878
rect 10277 5736 10597 5737
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 5671 10597 5672
rect 19610 5736 19930 5737
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 19610 5671 19930 5672
rect 19241 5394 19307 5397
rect 23473 5394 23539 5397
rect 19241 5392 23539 5394
rect 19241 5336 19246 5392
rect 19302 5336 23478 5392
rect 23534 5336 23539 5392
rect 19241 5334 23539 5336
rect 19241 5331 19307 5334
rect 23473 5331 23539 5334
rect 23657 5394 23723 5397
rect 27520 5394 28000 5424
rect 23657 5392 28000 5394
rect 23657 5336 23662 5392
rect 23718 5336 28000 5392
rect 23657 5334 28000 5336
rect 23657 5331 23723 5334
rect 27520 5304 28000 5334
rect 5610 5192 5930 5193
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5930 5192
rect 5610 5127 5930 5128
rect 14944 5192 15264 5193
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 5127 15264 5128
rect 24277 5192 24597 5193
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 5127 24597 5128
rect 21541 4986 21607 4989
rect 23657 4986 23723 4989
rect 21541 4984 23723 4986
rect 21541 4928 21546 4984
rect 21602 4928 23662 4984
rect 23718 4928 23723 4984
rect 21541 4926 23723 4928
rect 21541 4923 21607 4926
rect 23657 4923 23723 4926
rect 15929 4850 15995 4853
rect 27520 4850 28000 4880
rect 15929 4848 28000 4850
rect 15929 4792 15934 4848
rect 15990 4792 28000 4848
rect 15929 4790 28000 4792
rect 15929 4787 15995 4790
rect 27520 4760 28000 4790
rect 23473 4714 23539 4717
rect 20118 4712 23539 4714
rect 20118 4656 23478 4712
rect 23534 4656 23539 4712
rect 20118 4654 23539 4656
rect 10277 4648 10597 4649
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 4583 10597 4584
rect 19610 4648 19930 4649
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 4583 19930 4584
rect 17953 4306 18019 4309
rect 20118 4306 20178 4654
rect 23473 4651 23539 4654
rect 17953 4304 20178 4306
rect 17953 4248 17958 4304
rect 18014 4248 20178 4304
rect 17953 4246 20178 4248
rect 17953 4243 18019 4246
rect 24669 4170 24735 4173
rect 27520 4170 28000 4200
rect 24669 4168 28000 4170
rect 24669 4112 24674 4168
rect 24730 4112 28000 4168
rect 24669 4110 28000 4112
rect 24669 4107 24735 4110
rect 5610 4104 5930 4105
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5930 4104
rect 5610 4039 5930 4040
rect 14944 4104 15264 4105
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 4039 15264 4040
rect 24277 4104 24597 4105
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 27520 4080 28000 4110
rect 24277 4039 24597 4040
rect 24761 3762 24827 3765
rect 26233 3762 26299 3765
rect 24761 3760 26299 3762
rect 24761 3704 24766 3760
rect 24822 3704 26238 3760
rect 26294 3704 26299 3760
rect 24761 3702 26299 3704
rect 24761 3699 24827 3702
rect 26233 3699 26299 3702
rect 25221 3626 25287 3629
rect 27520 3626 28000 3656
rect 25221 3624 28000 3626
rect 25221 3568 25226 3624
rect 25282 3568 28000 3624
rect 25221 3566 28000 3568
rect 25221 3563 25287 3566
rect 10277 3560 10597 3561
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 3495 10597 3496
rect 19610 3560 19930 3561
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 27520 3536 28000 3566
rect 19610 3495 19930 3496
rect 24025 3218 24091 3221
rect 24025 3216 24778 3218
rect 24025 3160 24030 3216
rect 24086 3160 24778 3216
rect 24025 3158 24778 3160
rect 24025 3155 24091 3158
rect 5610 3016 5930 3017
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5930 3016
rect 5610 2951 5930 2952
rect 14944 3016 15264 3017
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 2951 15264 2952
rect 24277 3016 24597 3017
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 2951 24597 2952
rect 24718 2946 24778 3158
rect 27520 2946 28000 2976
rect 24718 2886 28000 2946
rect 27520 2856 28000 2886
rect 10277 2472 10597 2473
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 2407 10597 2408
rect 19610 2472 19930 2473
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 2407 19930 2408
rect 23473 2402 23539 2405
rect 27520 2402 28000 2432
rect 23473 2400 28000 2402
rect 23473 2344 23478 2400
rect 23534 2344 28000 2400
rect 23473 2342 28000 2344
rect 23473 2339 23539 2342
rect 27520 2312 28000 2342
rect 23749 2130 23815 2133
rect 23749 2128 25698 2130
rect 23749 2072 23754 2128
rect 23810 2072 25698 2128
rect 23749 2070 25698 2072
rect 23749 2067 23815 2070
rect 5610 1928 5930 1929
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5930 1928
rect 5610 1863 5930 1864
rect 14944 1928 15264 1929
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1863 15264 1864
rect 24277 1928 24597 1929
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1863 24597 1864
rect 25638 1858 25698 2070
rect 27520 1858 28000 1888
rect 25638 1798 28000 1858
rect 27520 1768 28000 1798
rect 24117 1178 24183 1181
rect 27520 1178 28000 1208
rect 24117 1176 28000 1178
rect 24117 1120 24122 1176
rect 24178 1120 28000 1176
rect 24117 1118 28000 1120
rect 24117 1115 24183 1118
rect 27520 1088 28000 1118
rect 23657 634 23723 637
rect 27520 634 28000 664
rect 23657 632 28000 634
rect 23657 576 23662 632
rect 23718 576 28000 632
rect 23657 574 28000 576
rect 23657 571 23723 574
rect 27520 544 28000 574
rect 23565 90 23631 93
rect 27520 90 28000 120
rect 23565 88 28000 90
rect 23565 32 23570 88
rect 23626 32 28000 88
rect 23565 30 28000 32
rect 23565 27 23631 30
rect 27520 0 28000 30
<< via3 >>
rect 10285 25316 10349 25320
rect 10285 25260 10289 25316
rect 10289 25260 10345 25316
rect 10345 25260 10349 25316
rect 10285 25256 10349 25260
rect 10365 25316 10429 25320
rect 10365 25260 10369 25316
rect 10369 25260 10425 25316
rect 10425 25260 10429 25316
rect 10365 25256 10429 25260
rect 10445 25316 10509 25320
rect 10445 25260 10449 25316
rect 10449 25260 10505 25316
rect 10505 25260 10509 25316
rect 10445 25256 10509 25260
rect 10525 25316 10589 25320
rect 10525 25260 10529 25316
rect 10529 25260 10585 25316
rect 10585 25260 10589 25316
rect 10525 25256 10589 25260
rect 19618 25316 19682 25320
rect 19618 25260 19622 25316
rect 19622 25260 19678 25316
rect 19678 25260 19682 25316
rect 19618 25256 19682 25260
rect 19698 25316 19762 25320
rect 19698 25260 19702 25316
rect 19702 25260 19758 25316
rect 19758 25260 19762 25316
rect 19698 25256 19762 25260
rect 19778 25316 19842 25320
rect 19778 25260 19782 25316
rect 19782 25260 19838 25316
rect 19838 25260 19842 25316
rect 19778 25256 19842 25260
rect 19858 25316 19922 25320
rect 19858 25260 19862 25316
rect 19862 25260 19918 25316
rect 19918 25260 19922 25316
rect 19858 25256 19922 25260
rect 5618 24772 5682 24776
rect 5618 24716 5622 24772
rect 5622 24716 5678 24772
rect 5678 24716 5682 24772
rect 5618 24712 5682 24716
rect 5698 24772 5762 24776
rect 5698 24716 5702 24772
rect 5702 24716 5758 24772
rect 5758 24716 5762 24772
rect 5698 24712 5762 24716
rect 5778 24772 5842 24776
rect 5778 24716 5782 24772
rect 5782 24716 5838 24772
rect 5838 24716 5842 24772
rect 5778 24712 5842 24716
rect 5858 24772 5922 24776
rect 5858 24716 5862 24772
rect 5862 24716 5918 24772
rect 5918 24716 5922 24772
rect 5858 24712 5922 24716
rect 14952 24772 15016 24776
rect 14952 24716 14956 24772
rect 14956 24716 15012 24772
rect 15012 24716 15016 24772
rect 14952 24712 15016 24716
rect 15032 24772 15096 24776
rect 15032 24716 15036 24772
rect 15036 24716 15092 24772
rect 15092 24716 15096 24772
rect 15032 24712 15096 24716
rect 15112 24772 15176 24776
rect 15112 24716 15116 24772
rect 15116 24716 15172 24772
rect 15172 24716 15176 24772
rect 15112 24712 15176 24716
rect 15192 24772 15256 24776
rect 15192 24716 15196 24772
rect 15196 24716 15252 24772
rect 15252 24716 15256 24772
rect 15192 24712 15256 24716
rect 24285 24772 24349 24776
rect 24285 24716 24289 24772
rect 24289 24716 24345 24772
rect 24345 24716 24349 24772
rect 24285 24712 24349 24716
rect 24365 24772 24429 24776
rect 24365 24716 24369 24772
rect 24369 24716 24425 24772
rect 24425 24716 24429 24772
rect 24365 24712 24429 24716
rect 24445 24772 24509 24776
rect 24445 24716 24449 24772
rect 24449 24716 24505 24772
rect 24505 24716 24509 24772
rect 24445 24712 24509 24716
rect 24525 24772 24589 24776
rect 24525 24716 24529 24772
rect 24529 24716 24585 24772
rect 24585 24716 24589 24772
rect 24525 24712 24589 24716
rect 10285 24228 10349 24232
rect 10285 24172 10289 24228
rect 10289 24172 10345 24228
rect 10345 24172 10349 24228
rect 10285 24168 10349 24172
rect 10365 24228 10429 24232
rect 10365 24172 10369 24228
rect 10369 24172 10425 24228
rect 10425 24172 10429 24228
rect 10365 24168 10429 24172
rect 10445 24228 10509 24232
rect 10445 24172 10449 24228
rect 10449 24172 10505 24228
rect 10505 24172 10509 24228
rect 10445 24168 10509 24172
rect 10525 24228 10589 24232
rect 10525 24172 10529 24228
rect 10529 24172 10585 24228
rect 10585 24172 10589 24228
rect 10525 24168 10589 24172
rect 19618 24228 19682 24232
rect 19618 24172 19622 24228
rect 19622 24172 19678 24228
rect 19678 24172 19682 24228
rect 19618 24168 19682 24172
rect 19698 24228 19762 24232
rect 19698 24172 19702 24228
rect 19702 24172 19758 24228
rect 19758 24172 19762 24228
rect 19698 24168 19762 24172
rect 19778 24228 19842 24232
rect 19778 24172 19782 24228
rect 19782 24172 19838 24228
rect 19838 24172 19842 24228
rect 19778 24168 19842 24172
rect 19858 24228 19922 24232
rect 19858 24172 19862 24228
rect 19862 24172 19918 24228
rect 19918 24172 19922 24228
rect 19858 24168 19922 24172
rect 5618 23684 5682 23688
rect 5618 23628 5622 23684
rect 5622 23628 5678 23684
rect 5678 23628 5682 23684
rect 5618 23624 5682 23628
rect 5698 23684 5762 23688
rect 5698 23628 5702 23684
rect 5702 23628 5758 23684
rect 5758 23628 5762 23684
rect 5698 23624 5762 23628
rect 5778 23684 5842 23688
rect 5778 23628 5782 23684
rect 5782 23628 5838 23684
rect 5838 23628 5842 23684
rect 5778 23624 5842 23628
rect 5858 23684 5922 23688
rect 5858 23628 5862 23684
rect 5862 23628 5918 23684
rect 5918 23628 5922 23684
rect 5858 23624 5922 23628
rect 14952 23684 15016 23688
rect 14952 23628 14956 23684
rect 14956 23628 15012 23684
rect 15012 23628 15016 23684
rect 14952 23624 15016 23628
rect 15032 23684 15096 23688
rect 15032 23628 15036 23684
rect 15036 23628 15092 23684
rect 15092 23628 15096 23684
rect 15032 23624 15096 23628
rect 15112 23684 15176 23688
rect 15112 23628 15116 23684
rect 15116 23628 15172 23684
rect 15172 23628 15176 23684
rect 15112 23624 15176 23628
rect 15192 23684 15256 23688
rect 15192 23628 15196 23684
rect 15196 23628 15252 23684
rect 15252 23628 15256 23684
rect 15192 23624 15256 23628
rect 24285 23684 24349 23688
rect 24285 23628 24289 23684
rect 24289 23628 24345 23684
rect 24345 23628 24349 23684
rect 24285 23624 24349 23628
rect 24365 23684 24429 23688
rect 24365 23628 24369 23684
rect 24369 23628 24425 23684
rect 24425 23628 24429 23684
rect 24365 23624 24429 23628
rect 24445 23684 24509 23688
rect 24445 23628 24449 23684
rect 24449 23628 24505 23684
rect 24505 23628 24509 23684
rect 24445 23624 24509 23628
rect 24525 23684 24589 23688
rect 24525 23628 24529 23684
rect 24529 23628 24585 23684
rect 24585 23628 24589 23684
rect 24525 23624 24589 23628
rect 10285 23140 10349 23144
rect 10285 23084 10289 23140
rect 10289 23084 10345 23140
rect 10345 23084 10349 23140
rect 10285 23080 10349 23084
rect 10365 23140 10429 23144
rect 10365 23084 10369 23140
rect 10369 23084 10425 23140
rect 10425 23084 10429 23140
rect 10365 23080 10429 23084
rect 10445 23140 10509 23144
rect 10445 23084 10449 23140
rect 10449 23084 10505 23140
rect 10505 23084 10509 23140
rect 10445 23080 10509 23084
rect 10525 23140 10589 23144
rect 10525 23084 10529 23140
rect 10529 23084 10585 23140
rect 10585 23084 10589 23140
rect 10525 23080 10589 23084
rect 19618 23140 19682 23144
rect 19618 23084 19622 23140
rect 19622 23084 19678 23140
rect 19678 23084 19682 23140
rect 19618 23080 19682 23084
rect 19698 23140 19762 23144
rect 19698 23084 19702 23140
rect 19702 23084 19758 23140
rect 19758 23084 19762 23140
rect 19698 23080 19762 23084
rect 19778 23140 19842 23144
rect 19778 23084 19782 23140
rect 19782 23084 19838 23140
rect 19838 23084 19842 23140
rect 19778 23080 19842 23084
rect 19858 23140 19922 23144
rect 19858 23084 19862 23140
rect 19862 23084 19918 23140
rect 19918 23084 19922 23140
rect 19858 23080 19922 23084
rect 5618 22596 5682 22600
rect 5618 22540 5622 22596
rect 5622 22540 5678 22596
rect 5678 22540 5682 22596
rect 5618 22536 5682 22540
rect 5698 22596 5762 22600
rect 5698 22540 5702 22596
rect 5702 22540 5758 22596
rect 5758 22540 5762 22596
rect 5698 22536 5762 22540
rect 5778 22596 5842 22600
rect 5778 22540 5782 22596
rect 5782 22540 5838 22596
rect 5838 22540 5842 22596
rect 5778 22536 5842 22540
rect 5858 22596 5922 22600
rect 5858 22540 5862 22596
rect 5862 22540 5918 22596
rect 5918 22540 5922 22596
rect 5858 22536 5922 22540
rect 14952 22596 15016 22600
rect 14952 22540 14956 22596
rect 14956 22540 15012 22596
rect 15012 22540 15016 22596
rect 14952 22536 15016 22540
rect 15032 22596 15096 22600
rect 15032 22540 15036 22596
rect 15036 22540 15092 22596
rect 15092 22540 15096 22596
rect 15032 22536 15096 22540
rect 15112 22596 15176 22600
rect 15112 22540 15116 22596
rect 15116 22540 15172 22596
rect 15172 22540 15176 22596
rect 15112 22536 15176 22540
rect 15192 22596 15256 22600
rect 15192 22540 15196 22596
rect 15196 22540 15252 22596
rect 15252 22540 15256 22596
rect 15192 22536 15256 22540
rect 24285 22596 24349 22600
rect 24285 22540 24289 22596
rect 24289 22540 24345 22596
rect 24345 22540 24349 22596
rect 24285 22536 24349 22540
rect 24365 22596 24429 22600
rect 24365 22540 24369 22596
rect 24369 22540 24425 22596
rect 24425 22540 24429 22596
rect 24365 22536 24429 22540
rect 24445 22596 24509 22600
rect 24445 22540 24449 22596
rect 24449 22540 24505 22596
rect 24505 22540 24509 22596
rect 24445 22536 24509 22540
rect 24525 22596 24589 22600
rect 24525 22540 24529 22596
rect 24529 22540 24585 22596
rect 24585 22540 24589 22596
rect 24525 22536 24589 22540
rect 10285 22052 10349 22056
rect 10285 21996 10289 22052
rect 10289 21996 10345 22052
rect 10345 21996 10349 22052
rect 10285 21992 10349 21996
rect 10365 22052 10429 22056
rect 10365 21996 10369 22052
rect 10369 21996 10425 22052
rect 10425 21996 10429 22052
rect 10365 21992 10429 21996
rect 10445 22052 10509 22056
rect 10445 21996 10449 22052
rect 10449 21996 10505 22052
rect 10505 21996 10509 22052
rect 10445 21992 10509 21996
rect 10525 22052 10589 22056
rect 10525 21996 10529 22052
rect 10529 21996 10585 22052
rect 10585 21996 10589 22052
rect 10525 21992 10589 21996
rect 19618 22052 19682 22056
rect 19618 21996 19622 22052
rect 19622 21996 19678 22052
rect 19678 21996 19682 22052
rect 19618 21992 19682 21996
rect 19698 22052 19762 22056
rect 19698 21996 19702 22052
rect 19702 21996 19758 22052
rect 19758 21996 19762 22052
rect 19698 21992 19762 21996
rect 19778 22052 19842 22056
rect 19778 21996 19782 22052
rect 19782 21996 19838 22052
rect 19838 21996 19842 22052
rect 19778 21992 19842 21996
rect 19858 22052 19922 22056
rect 19858 21996 19862 22052
rect 19862 21996 19918 22052
rect 19918 21996 19922 22052
rect 19858 21992 19922 21996
rect 5618 21508 5682 21512
rect 5618 21452 5622 21508
rect 5622 21452 5678 21508
rect 5678 21452 5682 21508
rect 5618 21448 5682 21452
rect 5698 21508 5762 21512
rect 5698 21452 5702 21508
rect 5702 21452 5758 21508
rect 5758 21452 5762 21508
rect 5698 21448 5762 21452
rect 5778 21508 5842 21512
rect 5778 21452 5782 21508
rect 5782 21452 5838 21508
rect 5838 21452 5842 21508
rect 5778 21448 5842 21452
rect 5858 21508 5922 21512
rect 5858 21452 5862 21508
rect 5862 21452 5918 21508
rect 5918 21452 5922 21508
rect 5858 21448 5922 21452
rect 14952 21508 15016 21512
rect 14952 21452 14956 21508
rect 14956 21452 15012 21508
rect 15012 21452 15016 21508
rect 14952 21448 15016 21452
rect 15032 21508 15096 21512
rect 15032 21452 15036 21508
rect 15036 21452 15092 21508
rect 15092 21452 15096 21508
rect 15032 21448 15096 21452
rect 15112 21508 15176 21512
rect 15112 21452 15116 21508
rect 15116 21452 15172 21508
rect 15172 21452 15176 21508
rect 15112 21448 15176 21452
rect 15192 21508 15256 21512
rect 15192 21452 15196 21508
rect 15196 21452 15252 21508
rect 15252 21452 15256 21508
rect 15192 21448 15256 21452
rect 24285 21508 24349 21512
rect 24285 21452 24289 21508
rect 24289 21452 24345 21508
rect 24345 21452 24349 21508
rect 24285 21448 24349 21452
rect 24365 21508 24429 21512
rect 24365 21452 24369 21508
rect 24369 21452 24425 21508
rect 24425 21452 24429 21508
rect 24365 21448 24429 21452
rect 24445 21508 24509 21512
rect 24445 21452 24449 21508
rect 24449 21452 24505 21508
rect 24505 21452 24509 21508
rect 24445 21448 24509 21452
rect 24525 21508 24589 21512
rect 24525 21452 24529 21508
rect 24529 21452 24585 21508
rect 24585 21452 24589 21508
rect 24525 21448 24589 21452
rect 10285 20964 10349 20968
rect 10285 20908 10289 20964
rect 10289 20908 10345 20964
rect 10345 20908 10349 20964
rect 10285 20904 10349 20908
rect 10365 20964 10429 20968
rect 10365 20908 10369 20964
rect 10369 20908 10425 20964
rect 10425 20908 10429 20964
rect 10365 20904 10429 20908
rect 10445 20964 10509 20968
rect 10445 20908 10449 20964
rect 10449 20908 10505 20964
rect 10505 20908 10509 20964
rect 10445 20904 10509 20908
rect 10525 20964 10589 20968
rect 10525 20908 10529 20964
rect 10529 20908 10585 20964
rect 10585 20908 10589 20964
rect 10525 20904 10589 20908
rect 19618 20964 19682 20968
rect 19618 20908 19622 20964
rect 19622 20908 19678 20964
rect 19678 20908 19682 20964
rect 19618 20904 19682 20908
rect 19698 20964 19762 20968
rect 19698 20908 19702 20964
rect 19702 20908 19758 20964
rect 19758 20908 19762 20964
rect 19698 20904 19762 20908
rect 19778 20964 19842 20968
rect 19778 20908 19782 20964
rect 19782 20908 19838 20964
rect 19838 20908 19842 20964
rect 19778 20904 19842 20908
rect 19858 20964 19922 20968
rect 19858 20908 19862 20964
rect 19862 20908 19918 20964
rect 19918 20908 19922 20964
rect 19858 20904 19922 20908
rect 5618 20420 5682 20424
rect 5618 20364 5622 20420
rect 5622 20364 5678 20420
rect 5678 20364 5682 20420
rect 5618 20360 5682 20364
rect 5698 20420 5762 20424
rect 5698 20364 5702 20420
rect 5702 20364 5758 20420
rect 5758 20364 5762 20420
rect 5698 20360 5762 20364
rect 5778 20420 5842 20424
rect 5778 20364 5782 20420
rect 5782 20364 5838 20420
rect 5838 20364 5842 20420
rect 5778 20360 5842 20364
rect 5858 20420 5922 20424
rect 5858 20364 5862 20420
rect 5862 20364 5918 20420
rect 5918 20364 5922 20420
rect 5858 20360 5922 20364
rect 14952 20420 15016 20424
rect 14952 20364 14956 20420
rect 14956 20364 15012 20420
rect 15012 20364 15016 20420
rect 14952 20360 15016 20364
rect 15032 20420 15096 20424
rect 15032 20364 15036 20420
rect 15036 20364 15092 20420
rect 15092 20364 15096 20420
rect 15032 20360 15096 20364
rect 15112 20420 15176 20424
rect 15112 20364 15116 20420
rect 15116 20364 15172 20420
rect 15172 20364 15176 20420
rect 15112 20360 15176 20364
rect 15192 20420 15256 20424
rect 15192 20364 15196 20420
rect 15196 20364 15252 20420
rect 15252 20364 15256 20420
rect 15192 20360 15256 20364
rect 24285 20420 24349 20424
rect 24285 20364 24289 20420
rect 24289 20364 24345 20420
rect 24345 20364 24349 20420
rect 24285 20360 24349 20364
rect 24365 20420 24429 20424
rect 24365 20364 24369 20420
rect 24369 20364 24425 20420
rect 24425 20364 24429 20420
rect 24365 20360 24429 20364
rect 24445 20420 24509 20424
rect 24445 20364 24449 20420
rect 24449 20364 24505 20420
rect 24505 20364 24509 20420
rect 24445 20360 24509 20364
rect 24525 20420 24589 20424
rect 24525 20364 24529 20420
rect 24529 20364 24585 20420
rect 24585 20364 24589 20420
rect 24525 20360 24589 20364
rect 10285 19876 10349 19880
rect 10285 19820 10289 19876
rect 10289 19820 10345 19876
rect 10345 19820 10349 19876
rect 10285 19816 10349 19820
rect 10365 19876 10429 19880
rect 10365 19820 10369 19876
rect 10369 19820 10425 19876
rect 10425 19820 10429 19876
rect 10365 19816 10429 19820
rect 10445 19876 10509 19880
rect 10445 19820 10449 19876
rect 10449 19820 10505 19876
rect 10505 19820 10509 19876
rect 10445 19816 10509 19820
rect 10525 19876 10589 19880
rect 10525 19820 10529 19876
rect 10529 19820 10585 19876
rect 10585 19820 10589 19876
rect 10525 19816 10589 19820
rect 19618 19876 19682 19880
rect 19618 19820 19622 19876
rect 19622 19820 19678 19876
rect 19678 19820 19682 19876
rect 19618 19816 19682 19820
rect 19698 19876 19762 19880
rect 19698 19820 19702 19876
rect 19702 19820 19758 19876
rect 19758 19820 19762 19876
rect 19698 19816 19762 19820
rect 19778 19876 19842 19880
rect 19778 19820 19782 19876
rect 19782 19820 19838 19876
rect 19838 19820 19842 19876
rect 19778 19816 19842 19820
rect 19858 19876 19922 19880
rect 19858 19820 19862 19876
rect 19862 19820 19918 19876
rect 19918 19820 19922 19876
rect 19858 19816 19922 19820
rect 5618 19332 5682 19336
rect 5618 19276 5622 19332
rect 5622 19276 5678 19332
rect 5678 19276 5682 19332
rect 5618 19272 5682 19276
rect 5698 19332 5762 19336
rect 5698 19276 5702 19332
rect 5702 19276 5758 19332
rect 5758 19276 5762 19332
rect 5698 19272 5762 19276
rect 5778 19332 5842 19336
rect 5778 19276 5782 19332
rect 5782 19276 5838 19332
rect 5838 19276 5842 19332
rect 5778 19272 5842 19276
rect 5858 19332 5922 19336
rect 5858 19276 5862 19332
rect 5862 19276 5918 19332
rect 5918 19276 5922 19332
rect 5858 19272 5922 19276
rect 14952 19332 15016 19336
rect 14952 19276 14956 19332
rect 14956 19276 15012 19332
rect 15012 19276 15016 19332
rect 14952 19272 15016 19276
rect 15032 19332 15096 19336
rect 15032 19276 15036 19332
rect 15036 19276 15092 19332
rect 15092 19276 15096 19332
rect 15032 19272 15096 19276
rect 15112 19332 15176 19336
rect 15112 19276 15116 19332
rect 15116 19276 15172 19332
rect 15172 19276 15176 19332
rect 15112 19272 15176 19276
rect 15192 19332 15256 19336
rect 15192 19276 15196 19332
rect 15196 19276 15252 19332
rect 15252 19276 15256 19332
rect 15192 19272 15256 19276
rect 24285 19332 24349 19336
rect 24285 19276 24289 19332
rect 24289 19276 24345 19332
rect 24345 19276 24349 19332
rect 24285 19272 24349 19276
rect 24365 19332 24429 19336
rect 24365 19276 24369 19332
rect 24369 19276 24425 19332
rect 24425 19276 24429 19332
rect 24365 19272 24429 19276
rect 24445 19332 24509 19336
rect 24445 19276 24449 19332
rect 24449 19276 24505 19332
rect 24505 19276 24509 19332
rect 24445 19272 24509 19276
rect 24525 19332 24589 19336
rect 24525 19276 24529 19332
rect 24529 19276 24585 19332
rect 24585 19276 24589 19332
rect 24525 19272 24589 19276
rect 10285 18788 10349 18792
rect 10285 18732 10289 18788
rect 10289 18732 10345 18788
rect 10345 18732 10349 18788
rect 10285 18728 10349 18732
rect 10365 18788 10429 18792
rect 10365 18732 10369 18788
rect 10369 18732 10425 18788
rect 10425 18732 10429 18788
rect 10365 18728 10429 18732
rect 10445 18788 10509 18792
rect 10445 18732 10449 18788
rect 10449 18732 10505 18788
rect 10505 18732 10509 18788
rect 10445 18728 10509 18732
rect 10525 18788 10589 18792
rect 10525 18732 10529 18788
rect 10529 18732 10585 18788
rect 10585 18732 10589 18788
rect 10525 18728 10589 18732
rect 19618 18788 19682 18792
rect 19618 18732 19622 18788
rect 19622 18732 19678 18788
rect 19678 18732 19682 18788
rect 19618 18728 19682 18732
rect 19698 18788 19762 18792
rect 19698 18732 19702 18788
rect 19702 18732 19758 18788
rect 19758 18732 19762 18788
rect 19698 18728 19762 18732
rect 19778 18788 19842 18792
rect 19778 18732 19782 18788
rect 19782 18732 19838 18788
rect 19838 18732 19842 18788
rect 19778 18728 19842 18732
rect 19858 18788 19922 18792
rect 19858 18732 19862 18788
rect 19862 18732 19918 18788
rect 19918 18732 19922 18788
rect 19858 18728 19922 18732
rect 5618 18244 5682 18248
rect 5618 18188 5622 18244
rect 5622 18188 5678 18244
rect 5678 18188 5682 18244
rect 5618 18184 5682 18188
rect 5698 18244 5762 18248
rect 5698 18188 5702 18244
rect 5702 18188 5758 18244
rect 5758 18188 5762 18244
rect 5698 18184 5762 18188
rect 5778 18244 5842 18248
rect 5778 18188 5782 18244
rect 5782 18188 5838 18244
rect 5838 18188 5842 18244
rect 5778 18184 5842 18188
rect 5858 18244 5922 18248
rect 5858 18188 5862 18244
rect 5862 18188 5918 18244
rect 5918 18188 5922 18244
rect 5858 18184 5922 18188
rect 14952 18244 15016 18248
rect 14952 18188 14956 18244
rect 14956 18188 15012 18244
rect 15012 18188 15016 18244
rect 14952 18184 15016 18188
rect 15032 18244 15096 18248
rect 15032 18188 15036 18244
rect 15036 18188 15092 18244
rect 15092 18188 15096 18244
rect 15032 18184 15096 18188
rect 15112 18244 15176 18248
rect 15112 18188 15116 18244
rect 15116 18188 15172 18244
rect 15172 18188 15176 18244
rect 15112 18184 15176 18188
rect 15192 18244 15256 18248
rect 15192 18188 15196 18244
rect 15196 18188 15252 18244
rect 15252 18188 15256 18244
rect 15192 18184 15256 18188
rect 24285 18244 24349 18248
rect 24285 18188 24289 18244
rect 24289 18188 24345 18244
rect 24345 18188 24349 18244
rect 24285 18184 24349 18188
rect 24365 18244 24429 18248
rect 24365 18188 24369 18244
rect 24369 18188 24425 18244
rect 24425 18188 24429 18244
rect 24365 18184 24429 18188
rect 24445 18244 24509 18248
rect 24445 18188 24449 18244
rect 24449 18188 24505 18244
rect 24505 18188 24509 18244
rect 24445 18184 24509 18188
rect 24525 18244 24589 18248
rect 24525 18188 24529 18244
rect 24529 18188 24585 18244
rect 24585 18188 24589 18244
rect 24525 18184 24589 18188
rect 10285 17700 10349 17704
rect 10285 17644 10289 17700
rect 10289 17644 10345 17700
rect 10345 17644 10349 17700
rect 10285 17640 10349 17644
rect 10365 17700 10429 17704
rect 10365 17644 10369 17700
rect 10369 17644 10425 17700
rect 10425 17644 10429 17700
rect 10365 17640 10429 17644
rect 10445 17700 10509 17704
rect 10445 17644 10449 17700
rect 10449 17644 10505 17700
rect 10505 17644 10509 17700
rect 10445 17640 10509 17644
rect 10525 17700 10589 17704
rect 10525 17644 10529 17700
rect 10529 17644 10585 17700
rect 10585 17644 10589 17700
rect 10525 17640 10589 17644
rect 19618 17700 19682 17704
rect 19618 17644 19622 17700
rect 19622 17644 19678 17700
rect 19678 17644 19682 17700
rect 19618 17640 19682 17644
rect 19698 17700 19762 17704
rect 19698 17644 19702 17700
rect 19702 17644 19758 17700
rect 19758 17644 19762 17700
rect 19698 17640 19762 17644
rect 19778 17700 19842 17704
rect 19778 17644 19782 17700
rect 19782 17644 19838 17700
rect 19838 17644 19842 17700
rect 19778 17640 19842 17644
rect 19858 17700 19922 17704
rect 19858 17644 19862 17700
rect 19862 17644 19918 17700
rect 19918 17644 19922 17700
rect 19858 17640 19922 17644
rect 5618 17156 5682 17160
rect 5618 17100 5622 17156
rect 5622 17100 5678 17156
rect 5678 17100 5682 17156
rect 5618 17096 5682 17100
rect 5698 17156 5762 17160
rect 5698 17100 5702 17156
rect 5702 17100 5758 17156
rect 5758 17100 5762 17156
rect 5698 17096 5762 17100
rect 5778 17156 5842 17160
rect 5778 17100 5782 17156
rect 5782 17100 5838 17156
rect 5838 17100 5842 17156
rect 5778 17096 5842 17100
rect 5858 17156 5922 17160
rect 5858 17100 5862 17156
rect 5862 17100 5918 17156
rect 5918 17100 5922 17156
rect 5858 17096 5922 17100
rect 14952 17156 15016 17160
rect 14952 17100 14956 17156
rect 14956 17100 15012 17156
rect 15012 17100 15016 17156
rect 14952 17096 15016 17100
rect 15032 17156 15096 17160
rect 15032 17100 15036 17156
rect 15036 17100 15092 17156
rect 15092 17100 15096 17156
rect 15032 17096 15096 17100
rect 15112 17156 15176 17160
rect 15112 17100 15116 17156
rect 15116 17100 15172 17156
rect 15172 17100 15176 17156
rect 15112 17096 15176 17100
rect 15192 17156 15256 17160
rect 15192 17100 15196 17156
rect 15196 17100 15252 17156
rect 15252 17100 15256 17156
rect 15192 17096 15256 17100
rect 24285 17156 24349 17160
rect 24285 17100 24289 17156
rect 24289 17100 24345 17156
rect 24345 17100 24349 17156
rect 24285 17096 24349 17100
rect 24365 17156 24429 17160
rect 24365 17100 24369 17156
rect 24369 17100 24425 17156
rect 24425 17100 24429 17156
rect 24365 17096 24429 17100
rect 24445 17156 24509 17160
rect 24445 17100 24449 17156
rect 24449 17100 24505 17156
rect 24505 17100 24509 17156
rect 24445 17096 24509 17100
rect 24525 17156 24589 17160
rect 24525 17100 24529 17156
rect 24529 17100 24585 17156
rect 24585 17100 24589 17156
rect 24525 17096 24589 17100
rect 10285 16612 10349 16616
rect 10285 16556 10289 16612
rect 10289 16556 10345 16612
rect 10345 16556 10349 16612
rect 10285 16552 10349 16556
rect 10365 16612 10429 16616
rect 10365 16556 10369 16612
rect 10369 16556 10425 16612
rect 10425 16556 10429 16612
rect 10365 16552 10429 16556
rect 10445 16612 10509 16616
rect 10445 16556 10449 16612
rect 10449 16556 10505 16612
rect 10505 16556 10509 16612
rect 10445 16552 10509 16556
rect 10525 16612 10589 16616
rect 10525 16556 10529 16612
rect 10529 16556 10585 16612
rect 10585 16556 10589 16612
rect 10525 16552 10589 16556
rect 19618 16612 19682 16616
rect 19618 16556 19622 16612
rect 19622 16556 19678 16612
rect 19678 16556 19682 16612
rect 19618 16552 19682 16556
rect 19698 16612 19762 16616
rect 19698 16556 19702 16612
rect 19702 16556 19758 16612
rect 19758 16556 19762 16612
rect 19698 16552 19762 16556
rect 19778 16612 19842 16616
rect 19778 16556 19782 16612
rect 19782 16556 19838 16612
rect 19838 16556 19842 16612
rect 19778 16552 19842 16556
rect 19858 16612 19922 16616
rect 19858 16556 19862 16612
rect 19862 16556 19918 16612
rect 19918 16556 19922 16612
rect 19858 16552 19922 16556
rect 5618 16068 5682 16072
rect 5618 16012 5622 16068
rect 5622 16012 5678 16068
rect 5678 16012 5682 16068
rect 5618 16008 5682 16012
rect 5698 16068 5762 16072
rect 5698 16012 5702 16068
rect 5702 16012 5758 16068
rect 5758 16012 5762 16068
rect 5698 16008 5762 16012
rect 5778 16068 5842 16072
rect 5778 16012 5782 16068
rect 5782 16012 5838 16068
rect 5838 16012 5842 16068
rect 5778 16008 5842 16012
rect 5858 16068 5922 16072
rect 5858 16012 5862 16068
rect 5862 16012 5918 16068
rect 5918 16012 5922 16068
rect 5858 16008 5922 16012
rect 14952 16068 15016 16072
rect 14952 16012 14956 16068
rect 14956 16012 15012 16068
rect 15012 16012 15016 16068
rect 14952 16008 15016 16012
rect 15032 16068 15096 16072
rect 15032 16012 15036 16068
rect 15036 16012 15092 16068
rect 15092 16012 15096 16068
rect 15032 16008 15096 16012
rect 15112 16068 15176 16072
rect 15112 16012 15116 16068
rect 15116 16012 15172 16068
rect 15172 16012 15176 16068
rect 15112 16008 15176 16012
rect 15192 16068 15256 16072
rect 15192 16012 15196 16068
rect 15196 16012 15252 16068
rect 15252 16012 15256 16068
rect 15192 16008 15256 16012
rect 24285 16068 24349 16072
rect 24285 16012 24289 16068
rect 24289 16012 24345 16068
rect 24345 16012 24349 16068
rect 24285 16008 24349 16012
rect 24365 16068 24429 16072
rect 24365 16012 24369 16068
rect 24369 16012 24425 16068
rect 24425 16012 24429 16068
rect 24365 16008 24429 16012
rect 24445 16068 24509 16072
rect 24445 16012 24449 16068
rect 24449 16012 24505 16068
rect 24505 16012 24509 16068
rect 24445 16008 24509 16012
rect 24525 16068 24589 16072
rect 24525 16012 24529 16068
rect 24529 16012 24585 16068
rect 24585 16012 24589 16068
rect 24525 16008 24589 16012
rect 10285 15524 10349 15528
rect 10285 15468 10289 15524
rect 10289 15468 10345 15524
rect 10345 15468 10349 15524
rect 10285 15464 10349 15468
rect 10365 15524 10429 15528
rect 10365 15468 10369 15524
rect 10369 15468 10425 15524
rect 10425 15468 10429 15524
rect 10365 15464 10429 15468
rect 10445 15524 10509 15528
rect 10445 15468 10449 15524
rect 10449 15468 10505 15524
rect 10505 15468 10509 15524
rect 10445 15464 10509 15468
rect 10525 15524 10589 15528
rect 10525 15468 10529 15524
rect 10529 15468 10585 15524
rect 10585 15468 10589 15524
rect 10525 15464 10589 15468
rect 19618 15524 19682 15528
rect 19618 15468 19622 15524
rect 19622 15468 19678 15524
rect 19678 15468 19682 15524
rect 19618 15464 19682 15468
rect 19698 15524 19762 15528
rect 19698 15468 19702 15524
rect 19702 15468 19758 15524
rect 19758 15468 19762 15524
rect 19698 15464 19762 15468
rect 19778 15524 19842 15528
rect 19778 15468 19782 15524
rect 19782 15468 19838 15524
rect 19838 15468 19842 15524
rect 19778 15464 19842 15468
rect 19858 15524 19922 15528
rect 19858 15468 19862 15524
rect 19862 15468 19918 15524
rect 19918 15468 19922 15524
rect 19858 15464 19922 15468
rect 5618 14980 5682 14984
rect 5618 14924 5622 14980
rect 5622 14924 5678 14980
rect 5678 14924 5682 14980
rect 5618 14920 5682 14924
rect 5698 14980 5762 14984
rect 5698 14924 5702 14980
rect 5702 14924 5758 14980
rect 5758 14924 5762 14980
rect 5698 14920 5762 14924
rect 5778 14980 5842 14984
rect 5778 14924 5782 14980
rect 5782 14924 5838 14980
rect 5838 14924 5842 14980
rect 5778 14920 5842 14924
rect 5858 14980 5922 14984
rect 5858 14924 5862 14980
rect 5862 14924 5918 14980
rect 5918 14924 5922 14980
rect 5858 14920 5922 14924
rect 14952 14980 15016 14984
rect 14952 14924 14956 14980
rect 14956 14924 15012 14980
rect 15012 14924 15016 14980
rect 14952 14920 15016 14924
rect 15032 14980 15096 14984
rect 15032 14924 15036 14980
rect 15036 14924 15092 14980
rect 15092 14924 15096 14980
rect 15032 14920 15096 14924
rect 15112 14980 15176 14984
rect 15112 14924 15116 14980
rect 15116 14924 15172 14980
rect 15172 14924 15176 14980
rect 15112 14920 15176 14924
rect 15192 14980 15256 14984
rect 15192 14924 15196 14980
rect 15196 14924 15252 14980
rect 15252 14924 15256 14980
rect 15192 14920 15256 14924
rect 24285 14980 24349 14984
rect 24285 14924 24289 14980
rect 24289 14924 24345 14980
rect 24345 14924 24349 14980
rect 24285 14920 24349 14924
rect 24365 14980 24429 14984
rect 24365 14924 24369 14980
rect 24369 14924 24425 14980
rect 24425 14924 24429 14980
rect 24365 14920 24429 14924
rect 24445 14980 24509 14984
rect 24445 14924 24449 14980
rect 24449 14924 24505 14980
rect 24505 14924 24509 14980
rect 24445 14920 24509 14924
rect 24525 14980 24589 14984
rect 24525 14924 24529 14980
rect 24529 14924 24585 14980
rect 24585 14924 24589 14980
rect 24525 14920 24589 14924
rect 10285 14436 10349 14440
rect 10285 14380 10289 14436
rect 10289 14380 10345 14436
rect 10345 14380 10349 14436
rect 10285 14376 10349 14380
rect 10365 14436 10429 14440
rect 10365 14380 10369 14436
rect 10369 14380 10425 14436
rect 10425 14380 10429 14436
rect 10365 14376 10429 14380
rect 10445 14436 10509 14440
rect 10445 14380 10449 14436
rect 10449 14380 10505 14436
rect 10505 14380 10509 14436
rect 10445 14376 10509 14380
rect 10525 14436 10589 14440
rect 10525 14380 10529 14436
rect 10529 14380 10585 14436
rect 10585 14380 10589 14436
rect 10525 14376 10589 14380
rect 19618 14436 19682 14440
rect 19618 14380 19622 14436
rect 19622 14380 19678 14436
rect 19678 14380 19682 14436
rect 19618 14376 19682 14380
rect 19698 14436 19762 14440
rect 19698 14380 19702 14436
rect 19702 14380 19758 14436
rect 19758 14380 19762 14436
rect 19698 14376 19762 14380
rect 19778 14436 19842 14440
rect 19778 14380 19782 14436
rect 19782 14380 19838 14436
rect 19838 14380 19842 14436
rect 19778 14376 19842 14380
rect 19858 14436 19922 14440
rect 19858 14380 19862 14436
rect 19862 14380 19918 14436
rect 19918 14380 19922 14436
rect 19858 14376 19922 14380
rect 5618 13892 5682 13896
rect 5618 13836 5622 13892
rect 5622 13836 5678 13892
rect 5678 13836 5682 13892
rect 5618 13832 5682 13836
rect 5698 13892 5762 13896
rect 5698 13836 5702 13892
rect 5702 13836 5758 13892
rect 5758 13836 5762 13892
rect 5698 13832 5762 13836
rect 5778 13892 5842 13896
rect 5778 13836 5782 13892
rect 5782 13836 5838 13892
rect 5838 13836 5842 13892
rect 5778 13832 5842 13836
rect 5858 13892 5922 13896
rect 5858 13836 5862 13892
rect 5862 13836 5918 13892
rect 5918 13836 5922 13892
rect 5858 13832 5922 13836
rect 14952 13892 15016 13896
rect 14952 13836 14956 13892
rect 14956 13836 15012 13892
rect 15012 13836 15016 13892
rect 14952 13832 15016 13836
rect 15032 13892 15096 13896
rect 15032 13836 15036 13892
rect 15036 13836 15092 13892
rect 15092 13836 15096 13892
rect 15032 13832 15096 13836
rect 15112 13892 15176 13896
rect 15112 13836 15116 13892
rect 15116 13836 15172 13892
rect 15172 13836 15176 13892
rect 15112 13832 15176 13836
rect 15192 13892 15256 13896
rect 15192 13836 15196 13892
rect 15196 13836 15252 13892
rect 15252 13836 15256 13892
rect 15192 13832 15256 13836
rect 24285 13892 24349 13896
rect 24285 13836 24289 13892
rect 24289 13836 24345 13892
rect 24345 13836 24349 13892
rect 24285 13832 24349 13836
rect 24365 13892 24429 13896
rect 24365 13836 24369 13892
rect 24369 13836 24425 13892
rect 24425 13836 24429 13892
rect 24365 13832 24429 13836
rect 24445 13892 24509 13896
rect 24445 13836 24449 13892
rect 24449 13836 24505 13892
rect 24505 13836 24509 13892
rect 24445 13832 24509 13836
rect 24525 13892 24589 13896
rect 24525 13836 24529 13892
rect 24529 13836 24585 13892
rect 24585 13836 24589 13892
rect 24525 13832 24589 13836
rect 10285 13348 10349 13352
rect 10285 13292 10289 13348
rect 10289 13292 10345 13348
rect 10345 13292 10349 13348
rect 10285 13288 10349 13292
rect 10365 13348 10429 13352
rect 10365 13292 10369 13348
rect 10369 13292 10425 13348
rect 10425 13292 10429 13348
rect 10365 13288 10429 13292
rect 10445 13348 10509 13352
rect 10445 13292 10449 13348
rect 10449 13292 10505 13348
rect 10505 13292 10509 13348
rect 10445 13288 10509 13292
rect 10525 13348 10589 13352
rect 10525 13292 10529 13348
rect 10529 13292 10585 13348
rect 10585 13292 10589 13348
rect 10525 13288 10589 13292
rect 19618 13348 19682 13352
rect 19618 13292 19622 13348
rect 19622 13292 19678 13348
rect 19678 13292 19682 13348
rect 19618 13288 19682 13292
rect 19698 13348 19762 13352
rect 19698 13292 19702 13348
rect 19702 13292 19758 13348
rect 19758 13292 19762 13348
rect 19698 13288 19762 13292
rect 19778 13348 19842 13352
rect 19778 13292 19782 13348
rect 19782 13292 19838 13348
rect 19838 13292 19842 13348
rect 19778 13288 19842 13292
rect 19858 13348 19922 13352
rect 19858 13292 19862 13348
rect 19862 13292 19918 13348
rect 19918 13292 19922 13348
rect 19858 13288 19922 13292
rect 5618 12804 5682 12808
rect 5618 12748 5622 12804
rect 5622 12748 5678 12804
rect 5678 12748 5682 12804
rect 5618 12744 5682 12748
rect 5698 12804 5762 12808
rect 5698 12748 5702 12804
rect 5702 12748 5758 12804
rect 5758 12748 5762 12804
rect 5698 12744 5762 12748
rect 5778 12804 5842 12808
rect 5778 12748 5782 12804
rect 5782 12748 5838 12804
rect 5838 12748 5842 12804
rect 5778 12744 5842 12748
rect 5858 12804 5922 12808
rect 5858 12748 5862 12804
rect 5862 12748 5918 12804
rect 5918 12748 5922 12804
rect 5858 12744 5922 12748
rect 14952 12804 15016 12808
rect 14952 12748 14956 12804
rect 14956 12748 15012 12804
rect 15012 12748 15016 12804
rect 14952 12744 15016 12748
rect 15032 12804 15096 12808
rect 15032 12748 15036 12804
rect 15036 12748 15092 12804
rect 15092 12748 15096 12804
rect 15032 12744 15096 12748
rect 15112 12804 15176 12808
rect 15112 12748 15116 12804
rect 15116 12748 15172 12804
rect 15172 12748 15176 12804
rect 15112 12744 15176 12748
rect 15192 12804 15256 12808
rect 15192 12748 15196 12804
rect 15196 12748 15252 12804
rect 15252 12748 15256 12804
rect 15192 12744 15256 12748
rect 24285 12804 24349 12808
rect 24285 12748 24289 12804
rect 24289 12748 24345 12804
rect 24345 12748 24349 12804
rect 24285 12744 24349 12748
rect 24365 12804 24429 12808
rect 24365 12748 24369 12804
rect 24369 12748 24425 12804
rect 24425 12748 24429 12804
rect 24365 12744 24429 12748
rect 24445 12804 24509 12808
rect 24445 12748 24449 12804
rect 24449 12748 24505 12804
rect 24505 12748 24509 12804
rect 24445 12744 24509 12748
rect 24525 12804 24589 12808
rect 24525 12748 24529 12804
rect 24529 12748 24585 12804
rect 24585 12748 24589 12804
rect 24525 12744 24589 12748
rect 10285 12260 10349 12264
rect 10285 12204 10289 12260
rect 10289 12204 10345 12260
rect 10345 12204 10349 12260
rect 10285 12200 10349 12204
rect 10365 12260 10429 12264
rect 10365 12204 10369 12260
rect 10369 12204 10425 12260
rect 10425 12204 10429 12260
rect 10365 12200 10429 12204
rect 10445 12260 10509 12264
rect 10445 12204 10449 12260
rect 10449 12204 10505 12260
rect 10505 12204 10509 12260
rect 10445 12200 10509 12204
rect 10525 12260 10589 12264
rect 10525 12204 10529 12260
rect 10529 12204 10585 12260
rect 10585 12204 10589 12260
rect 10525 12200 10589 12204
rect 19618 12260 19682 12264
rect 19618 12204 19622 12260
rect 19622 12204 19678 12260
rect 19678 12204 19682 12260
rect 19618 12200 19682 12204
rect 19698 12260 19762 12264
rect 19698 12204 19702 12260
rect 19702 12204 19758 12260
rect 19758 12204 19762 12260
rect 19698 12200 19762 12204
rect 19778 12260 19842 12264
rect 19778 12204 19782 12260
rect 19782 12204 19838 12260
rect 19838 12204 19842 12260
rect 19778 12200 19842 12204
rect 19858 12260 19922 12264
rect 19858 12204 19862 12260
rect 19862 12204 19918 12260
rect 19918 12204 19922 12260
rect 19858 12200 19922 12204
rect 5618 11716 5682 11720
rect 5618 11660 5622 11716
rect 5622 11660 5678 11716
rect 5678 11660 5682 11716
rect 5618 11656 5682 11660
rect 5698 11716 5762 11720
rect 5698 11660 5702 11716
rect 5702 11660 5758 11716
rect 5758 11660 5762 11716
rect 5698 11656 5762 11660
rect 5778 11716 5842 11720
rect 5778 11660 5782 11716
rect 5782 11660 5838 11716
rect 5838 11660 5842 11716
rect 5778 11656 5842 11660
rect 5858 11716 5922 11720
rect 5858 11660 5862 11716
rect 5862 11660 5918 11716
rect 5918 11660 5922 11716
rect 5858 11656 5922 11660
rect 14952 11716 15016 11720
rect 14952 11660 14956 11716
rect 14956 11660 15012 11716
rect 15012 11660 15016 11716
rect 14952 11656 15016 11660
rect 15032 11716 15096 11720
rect 15032 11660 15036 11716
rect 15036 11660 15092 11716
rect 15092 11660 15096 11716
rect 15032 11656 15096 11660
rect 15112 11716 15176 11720
rect 15112 11660 15116 11716
rect 15116 11660 15172 11716
rect 15172 11660 15176 11716
rect 15112 11656 15176 11660
rect 15192 11716 15256 11720
rect 15192 11660 15196 11716
rect 15196 11660 15252 11716
rect 15252 11660 15256 11716
rect 15192 11656 15256 11660
rect 24285 11716 24349 11720
rect 24285 11660 24289 11716
rect 24289 11660 24345 11716
rect 24345 11660 24349 11716
rect 24285 11656 24349 11660
rect 24365 11716 24429 11720
rect 24365 11660 24369 11716
rect 24369 11660 24425 11716
rect 24425 11660 24429 11716
rect 24365 11656 24429 11660
rect 24445 11716 24509 11720
rect 24445 11660 24449 11716
rect 24449 11660 24505 11716
rect 24505 11660 24509 11716
rect 24445 11656 24509 11660
rect 24525 11716 24589 11720
rect 24525 11660 24529 11716
rect 24529 11660 24585 11716
rect 24585 11660 24589 11716
rect 24525 11656 24589 11660
rect 10285 11172 10349 11176
rect 10285 11116 10289 11172
rect 10289 11116 10345 11172
rect 10345 11116 10349 11172
rect 10285 11112 10349 11116
rect 10365 11172 10429 11176
rect 10365 11116 10369 11172
rect 10369 11116 10425 11172
rect 10425 11116 10429 11172
rect 10365 11112 10429 11116
rect 10445 11172 10509 11176
rect 10445 11116 10449 11172
rect 10449 11116 10505 11172
rect 10505 11116 10509 11172
rect 10445 11112 10509 11116
rect 10525 11172 10589 11176
rect 10525 11116 10529 11172
rect 10529 11116 10585 11172
rect 10585 11116 10589 11172
rect 10525 11112 10589 11116
rect 19618 11172 19682 11176
rect 19618 11116 19622 11172
rect 19622 11116 19678 11172
rect 19678 11116 19682 11172
rect 19618 11112 19682 11116
rect 19698 11172 19762 11176
rect 19698 11116 19702 11172
rect 19702 11116 19758 11172
rect 19758 11116 19762 11172
rect 19698 11112 19762 11116
rect 19778 11172 19842 11176
rect 19778 11116 19782 11172
rect 19782 11116 19838 11172
rect 19838 11116 19842 11172
rect 19778 11112 19842 11116
rect 19858 11172 19922 11176
rect 19858 11116 19862 11172
rect 19862 11116 19918 11172
rect 19918 11116 19922 11172
rect 19858 11112 19922 11116
rect 5618 10628 5682 10632
rect 5618 10572 5622 10628
rect 5622 10572 5678 10628
rect 5678 10572 5682 10628
rect 5618 10568 5682 10572
rect 5698 10628 5762 10632
rect 5698 10572 5702 10628
rect 5702 10572 5758 10628
rect 5758 10572 5762 10628
rect 5698 10568 5762 10572
rect 5778 10628 5842 10632
rect 5778 10572 5782 10628
rect 5782 10572 5838 10628
rect 5838 10572 5842 10628
rect 5778 10568 5842 10572
rect 5858 10628 5922 10632
rect 5858 10572 5862 10628
rect 5862 10572 5918 10628
rect 5918 10572 5922 10628
rect 5858 10568 5922 10572
rect 14952 10628 15016 10632
rect 14952 10572 14956 10628
rect 14956 10572 15012 10628
rect 15012 10572 15016 10628
rect 14952 10568 15016 10572
rect 15032 10628 15096 10632
rect 15032 10572 15036 10628
rect 15036 10572 15092 10628
rect 15092 10572 15096 10628
rect 15032 10568 15096 10572
rect 15112 10628 15176 10632
rect 15112 10572 15116 10628
rect 15116 10572 15172 10628
rect 15172 10572 15176 10628
rect 15112 10568 15176 10572
rect 15192 10628 15256 10632
rect 15192 10572 15196 10628
rect 15196 10572 15252 10628
rect 15252 10572 15256 10628
rect 15192 10568 15256 10572
rect 24285 10628 24349 10632
rect 24285 10572 24289 10628
rect 24289 10572 24345 10628
rect 24345 10572 24349 10628
rect 24285 10568 24349 10572
rect 24365 10628 24429 10632
rect 24365 10572 24369 10628
rect 24369 10572 24425 10628
rect 24425 10572 24429 10628
rect 24365 10568 24429 10572
rect 24445 10628 24509 10632
rect 24445 10572 24449 10628
rect 24449 10572 24505 10628
rect 24505 10572 24509 10628
rect 24445 10568 24509 10572
rect 24525 10628 24589 10632
rect 24525 10572 24529 10628
rect 24529 10572 24585 10628
rect 24585 10572 24589 10628
rect 24525 10568 24589 10572
rect 10285 10084 10349 10088
rect 10285 10028 10289 10084
rect 10289 10028 10345 10084
rect 10345 10028 10349 10084
rect 10285 10024 10349 10028
rect 10365 10084 10429 10088
rect 10365 10028 10369 10084
rect 10369 10028 10425 10084
rect 10425 10028 10429 10084
rect 10365 10024 10429 10028
rect 10445 10084 10509 10088
rect 10445 10028 10449 10084
rect 10449 10028 10505 10084
rect 10505 10028 10509 10084
rect 10445 10024 10509 10028
rect 10525 10084 10589 10088
rect 10525 10028 10529 10084
rect 10529 10028 10585 10084
rect 10585 10028 10589 10084
rect 10525 10024 10589 10028
rect 19618 10084 19682 10088
rect 19618 10028 19622 10084
rect 19622 10028 19678 10084
rect 19678 10028 19682 10084
rect 19618 10024 19682 10028
rect 19698 10084 19762 10088
rect 19698 10028 19702 10084
rect 19702 10028 19758 10084
rect 19758 10028 19762 10084
rect 19698 10024 19762 10028
rect 19778 10084 19842 10088
rect 19778 10028 19782 10084
rect 19782 10028 19838 10084
rect 19838 10028 19842 10084
rect 19778 10024 19842 10028
rect 19858 10084 19922 10088
rect 19858 10028 19862 10084
rect 19862 10028 19918 10084
rect 19918 10028 19922 10084
rect 19858 10024 19922 10028
rect 5618 9540 5682 9544
rect 5618 9484 5622 9540
rect 5622 9484 5678 9540
rect 5678 9484 5682 9540
rect 5618 9480 5682 9484
rect 5698 9540 5762 9544
rect 5698 9484 5702 9540
rect 5702 9484 5758 9540
rect 5758 9484 5762 9540
rect 5698 9480 5762 9484
rect 5778 9540 5842 9544
rect 5778 9484 5782 9540
rect 5782 9484 5838 9540
rect 5838 9484 5842 9540
rect 5778 9480 5842 9484
rect 5858 9540 5922 9544
rect 5858 9484 5862 9540
rect 5862 9484 5918 9540
rect 5918 9484 5922 9540
rect 5858 9480 5922 9484
rect 14952 9540 15016 9544
rect 14952 9484 14956 9540
rect 14956 9484 15012 9540
rect 15012 9484 15016 9540
rect 14952 9480 15016 9484
rect 15032 9540 15096 9544
rect 15032 9484 15036 9540
rect 15036 9484 15092 9540
rect 15092 9484 15096 9540
rect 15032 9480 15096 9484
rect 15112 9540 15176 9544
rect 15112 9484 15116 9540
rect 15116 9484 15172 9540
rect 15172 9484 15176 9540
rect 15112 9480 15176 9484
rect 15192 9540 15256 9544
rect 15192 9484 15196 9540
rect 15196 9484 15252 9540
rect 15252 9484 15256 9540
rect 15192 9480 15256 9484
rect 24285 9540 24349 9544
rect 24285 9484 24289 9540
rect 24289 9484 24345 9540
rect 24345 9484 24349 9540
rect 24285 9480 24349 9484
rect 24365 9540 24429 9544
rect 24365 9484 24369 9540
rect 24369 9484 24425 9540
rect 24425 9484 24429 9540
rect 24365 9480 24429 9484
rect 24445 9540 24509 9544
rect 24445 9484 24449 9540
rect 24449 9484 24505 9540
rect 24505 9484 24509 9540
rect 24445 9480 24509 9484
rect 24525 9540 24589 9544
rect 24525 9484 24529 9540
rect 24529 9484 24585 9540
rect 24585 9484 24589 9540
rect 24525 9480 24589 9484
rect 10285 8996 10349 9000
rect 10285 8940 10289 8996
rect 10289 8940 10345 8996
rect 10345 8940 10349 8996
rect 10285 8936 10349 8940
rect 10365 8996 10429 9000
rect 10365 8940 10369 8996
rect 10369 8940 10425 8996
rect 10425 8940 10429 8996
rect 10365 8936 10429 8940
rect 10445 8996 10509 9000
rect 10445 8940 10449 8996
rect 10449 8940 10505 8996
rect 10505 8940 10509 8996
rect 10445 8936 10509 8940
rect 10525 8996 10589 9000
rect 10525 8940 10529 8996
rect 10529 8940 10585 8996
rect 10585 8940 10589 8996
rect 10525 8936 10589 8940
rect 19618 8996 19682 9000
rect 19618 8940 19622 8996
rect 19622 8940 19678 8996
rect 19678 8940 19682 8996
rect 19618 8936 19682 8940
rect 19698 8996 19762 9000
rect 19698 8940 19702 8996
rect 19702 8940 19758 8996
rect 19758 8940 19762 8996
rect 19698 8936 19762 8940
rect 19778 8996 19842 9000
rect 19778 8940 19782 8996
rect 19782 8940 19838 8996
rect 19838 8940 19842 8996
rect 19778 8936 19842 8940
rect 19858 8996 19922 9000
rect 19858 8940 19862 8996
rect 19862 8940 19918 8996
rect 19918 8940 19922 8996
rect 19858 8936 19922 8940
rect 5618 8452 5682 8456
rect 5618 8396 5622 8452
rect 5622 8396 5678 8452
rect 5678 8396 5682 8452
rect 5618 8392 5682 8396
rect 5698 8452 5762 8456
rect 5698 8396 5702 8452
rect 5702 8396 5758 8452
rect 5758 8396 5762 8452
rect 5698 8392 5762 8396
rect 5778 8452 5842 8456
rect 5778 8396 5782 8452
rect 5782 8396 5838 8452
rect 5838 8396 5842 8452
rect 5778 8392 5842 8396
rect 5858 8452 5922 8456
rect 5858 8396 5862 8452
rect 5862 8396 5918 8452
rect 5918 8396 5922 8452
rect 5858 8392 5922 8396
rect 14952 8452 15016 8456
rect 14952 8396 14956 8452
rect 14956 8396 15012 8452
rect 15012 8396 15016 8452
rect 14952 8392 15016 8396
rect 15032 8452 15096 8456
rect 15032 8396 15036 8452
rect 15036 8396 15092 8452
rect 15092 8396 15096 8452
rect 15032 8392 15096 8396
rect 15112 8452 15176 8456
rect 15112 8396 15116 8452
rect 15116 8396 15172 8452
rect 15172 8396 15176 8452
rect 15112 8392 15176 8396
rect 15192 8452 15256 8456
rect 15192 8396 15196 8452
rect 15196 8396 15252 8452
rect 15252 8396 15256 8452
rect 15192 8392 15256 8396
rect 24285 8452 24349 8456
rect 24285 8396 24289 8452
rect 24289 8396 24345 8452
rect 24345 8396 24349 8452
rect 24285 8392 24349 8396
rect 24365 8452 24429 8456
rect 24365 8396 24369 8452
rect 24369 8396 24425 8452
rect 24425 8396 24429 8452
rect 24365 8392 24429 8396
rect 24445 8452 24509 8456
rect 24445 8396 24449 8452
rect 24449 8396 24505 8452
rect 24505 8396 24509 8452
rect 24445 8392 24509 8396
rect 24525 8452 24589 8456
rect 24525 8396 24529 8452
rect 24529 8396 24585 8452
rect 24585 8396 24589 8452
rect 24525 8392 24589 8396
rect 10285 7908 10349 7912
rect 10285 7852 10289 7908
rect 10289 7852 10345 7908
rect 10345 7852 10349 7908
rect 10285 7848 10349 7852
rect 10365 7908 10429 7912
rect 10365 7852 10369 7908
rect 10369 7852 10425 7908
rect 10425 7852 10429 7908
rect 10365 7848 10429 7852
rect 10445 7908 10509 7912
rect 10445 7852 10449 7908
rect 10449 7852 10505 7908
rect 10505 7852 10509 7908
rect 10445 7848 10509 7852
rect 10525 7908 10589 7912
rect 10525 7852 10529 7908
rect 10529 7852 10585 7908
rect 10585 7852 10589 7908
rect 10525 7848 10589 7852
rect 19618 7908 19682 7912
rect 19618 7852 19622 7908
rect 19622 7852 19678 7908
rect 19678 7852 19682 7908
rect 19618 7848 19682 7852
rect 19698 7908 19762 7912
rect 19698 7852 19702 7908
rect 19702 7852 19758 7908
rect 19758 7852 19762 7908
rect 19698 7848 19762 7852
rect 19778 7908 19842 7912
rect 19778 7852 19782 7908
rect 19782 7852 19838 7908
rect 19838 7852 19842 7908
rect 19778 7848 19842 7852
rect 19858 7908 19922 7912
rect 19858 7852 19862 7908
rect 19862 7852 19918 7908
rect 19918 7852 19922 7908
rect 19858 7848 19922 7852
rect 5618 7364 5682 7368
rect 5618 7308 5622 7364
rect 5622 7308 5678 7364
rect 5678 7308 5682 7364
rect 5618 7304 5682 7308
rect 5698 7364 5762 7368
rect 5698 7308 5702 7364
rect 5702 7308 5758 7364
rect 5758 7308 5762 7364
rect 5698 7304 5762 7308
rect 5778 7364 5842 7368
rect 5778 7308 5782 7364
rect 5782 7308 5838 7364
rect 5838 7308 5842 7364
rect 5778 7304 5842 7308
rect 5858 7364 5922 7368
rect 5858 7308 5862 7364
rect 5862 7308 5918 7364
rect 5918 7308 5922 7364
rect 5858 7304 5922 7308
rect 14952 7364 15016 7368
rect 14952 7308 14956 7364
rect 14956 7308 15012 7364
rect 15012 7308 15016 7364
rect 14952 7304 15016 7308
rect 15032 7364 15096 7368
rect 15032 7308 15036 7364
rect 15036 7308 15092 7364
rect 15092 7308 15096 7364
rect 15032 7304 15096 7308
rect 15112 7364 15176 7368
rect 15112 7308 15116 7364
rect 15116 7308 15172 7364
rect 15172 7308 15176 7364
rect 15112 7304 15176 7308
rect 15192 7364 15256 7368
rect 15192 7308 15196 7364
rect 15196 7308 15252 7364
rect 15252 7308 15256 7364
rect 15192 7304 15256 7308
rect 24285 7364 24349 7368
rect 24285 7308 24289 7364
rect 24289 7308 24345 7364
rect 24345 7308 24349 7364
rect 24285 7304 24349 7308
rect 24365 7364 24429 7368
rect 24365 7308 24369 7364
rect 24369 7308 24425 7364
rect 24425 7308 24429 7364
rect 24365 7304 24429 7308
rect 24445 7364 24509 7368
rect 24445 7308 24449 7364
rect 24449 7308 24505 7364
rect 24505 7308 24509 7364
rect 24445 7304 24509 7308
rect 24525 7364 24589 7368
rect 24525 7308 24529 7364
rect 24529 7308 24585 7364
rect 24585 7308 24589 7364
rect 24525 7304 24589 7308
rect 10285 6820 10349 6824
rect 10285 6764 10289 6820
rect 10289 6764 10345 6820
rect 10345 6764 10349 6820
rect 10285 6760 10349 6764
rect 10365 6820 10429 6824
rect 10365 6764 10369 6820
rect 10369 6764 10425 6820
rect 10425 6764 10429 6820
rect 10365 6760 10429 6764
rect 10445 6820 10509 6824
rect 10445 6764 10449 6820
rect 10449 6764 10505 6820
rect 10505 6764 10509 6820
rect 10445 6760 10509 6764
rect 10525 6820 10589 6824
rect 10525 6764 10529 6820
rect 10529 6764 10585 6820
rect 10585 6764 10589 6820
rect 10525 6760 10589 6764
rect 19618 6820 19682 6824
rect 19618 6764 19622 6820
rect 19622 6764 19678 6820
rect 19678 6764 19682 6820
rect 19618 6760 19682 6764
rect 19698 6820 19762 6824
rect 19698 6764 19702 6820
rect 19702 6764 19758 6820
rect 19758 6764 19762 6820
rect 19698 6760 19762 6764
rect 19778 6820 19842 6824
rect 19778 6764 19782 6820
rect 19782 6764 19838 6820
rect 19838 6764 19842 6820
rect 19778 6760 19842 6764
rect 19858 6820 19922 6824
rect 19858 6764 19862 6820
rect 19862 6764 19918 6820
rect 19918 6764 19922 6820
rect 19858 6760 19922 6764
rect 5618 6276 5682 6280
rect 5618 6220 5622 6276
rect 5622 6220 5678 6276
rect 5678 6220 5682 6276
rect 5618 6216 5682 6220
rect 5698 6276 5762 6280
rect 5698 6220 5702 6276
rect 5702 6220 5758 6276
rect 5758 6220 5762 6276
rect 5698 6216 5762 6220
rect 5778 6276 5842 6280
rect 5778 6220 5782 6276
rect 5782 6220 5838 6276
rect 5838 6220 5842 6276
rect 5778 6216 5842 6220
rect 5858 6276 5922 6280
rect 5858 6220 5862 6276
rect 5862 6220 5918 6276
rect 5918 6220 5922 6276
rect 5858 6216 5922 6220
rect 14952 6276 15016 6280
rect 14952 6220 14956 6276
rect 14956 6220 15012 6276
rect 15012 6220 15016 6276
rect 14952 6216 15016 6220
rect 15032 6276 15096 6280
rect 15032 6220 15036 6276
rect 15036 6220 15092 6276
rect 15092 6220 15096 6276
rect 15032 6216 15096 6220
rect 15112 6276 15176 6280
rect 15112 6220 15116 6276
rect 15116 6220 15172 6276
rect 15172 6220 15176 6276
rect 15112 6216 15176 6220
rect 15192 6276 15256 6280
rect 15192 6220 15196 6276
rect 15196 6220 15252 6276
rect 15252 6220 15256 6276
rect 15192 6216 15256 6220
rect 24285 6276 24349 6280
rect 24285 6220 24289 6276
rect 24289 6220 24345 6276
rect 24345 6220 24349 6276
rect 24285 6216 24349 6220
rect 24365 6276 24429 6280
rect 24365 6220 24369 6276
rect 24369 6220 24425 6276
rect 24425 6220 24429 6276
rect 24365 6216 24429 6220
rect 24445 6276 24509 6280
rect 24445 6220 24449 6276
rect 24449 6220 24505 6276
rect 24505 6220 24509 6276
rect 24445 6216 24509 6220
rect 24525 6276 24589 6280
rect 24525 6220 24529 6276
rect 24529 6220 24585 6276
rect 24585 6220 24589 6276
rect 24525 6216 24589 6220
rect 10285 5732 10349 5736
rect 10285 5676 10289 5732
rect 10289 5676 10345 5732
rect 10345 5676 10349 5732
rect 10285 5672 10349 5676
rect 10365 5732 10429 5736
rect 10365 5676 10369 5732
rect 10369 5676 10425 5732
rect 10425 5676 10429 5732
rect 10365 5672 10429 5676
rect 10445 5732 10509 5736
rect 10445 5676 10449 5732
rect 10449 5676 10505 5732
rect 10505 5676 10509 5732
rect 10445 5672 10509 5676
rect 10525 5732 10589 5736
rect 10525 5676 10529 5732
rect 10529 5676 10585 5732
rect 10585 5676 10589 5732
rect 10525 5672 10589 5676
rect 19618 5732 19682 5736
rect 19618 5676 19622 5732
rect 19622 5676 19678 5732
rect 19678 5676 19682 5732
rect 19618 5672 19682 5676
rect 19698 5732 19762 5736
rect 19698 5676 19702 5732
rect 19702 5676 19758 5732
rect 19758 5676 19762 5732
rect 19698 5672 19762 5676
rect 19778 5732 19842 5736
rect 19778 5676 19782 5732
rect 19782 5676 19838 5732
rect 19838 5676 19842 5732
rect 19778 5672 19842 5676
rect 19858 5732 19922 5736
rect 19858 5676 19862 5732
rect 19862 5676 19918 5732
rect 19918 5676 19922 5732
rect 19858 5672 19922 5676
rect 5618 5188 5682 5192
rect 5618 5132 5622 5188
rect 5622 5132 5678 5188
rect 5678 5132 5682 5188
rect 5618 5128 5682 5132
rect 5698 5188 5762 5192
rect 5698 5132 5702 5188
rect 5702 5132 5758 5188
rect 5758 5132 5762 5188
rect 5698 5128 5762 5132
rect 5778 5188 5842 5192
rect 5778 5132 5782 5188
rect 5782 5132 5838 5188
rect 5838 5132 5842 5188
rect 5778 5128 5842 5132
rect 5858 5188 5922 5192
rect 5858 5132 5862 5188
rect 5862 5132 5918 5188
rect 5918 5132 5922 5188
rect 5858 5128 5922 5132
rect 14952 5188 15016 5192
rect 14952 5132 14956 5188
rect 14956 5132 15012 5188
rect 15012 5132 15016 5188
rect 14952 5128 15016 5132
rect 15032 5188 15096 5192
rect 15032 5132 15036 5188
rect 15036 5132 15092 5188
rect 15092 5132 15096 5188
rect 15032 5128 15096 5132
rect 15112 5188 15176 5192
rect 15112 5132 15116 5188
rect 15116 5132 15172 5188
rect 15172 5132 15176 5188
rect 15112 5128 15176 5132
rect 15192 5188 15256 5192
rect 15192 5132 15196 5188
rect 15196 5132 15252 5188
rect 15252 5132 15256 5188
rect 15192 5128 15256 5132
rect 24285 5188 24349 5192
rect 24285 5132 24289 5188
rect 24289 5132 24345 5188
rect 24345 5132 24349 5188
rect 24285 5128 24349 5132
rect 24365 5188 24429 5192
rect 24365 5132 24369 5188
rect 24369 5132 24425 5188
rect 24425 5132 24429 5188
rect 24365 5128 24429 5132
rect 24445 5188 24509 5192
rect 24445 5132 24449 5188
rect 24449 5132 24505 5188
rect 24505 5132 24509 5188
rect 24445 5128 24509 5132
rect 24525 5188 24589 5192
rect 24525 5132 24529 5188
rect 24529 5132 24585 5188
rect 24585 5132 24589 5188
rect 24525 5128 24589 5132
rect 10285 4644 10349 4648
rect 10285 4588 10289 4644
rect 10289 4588 10345 4644
rect 10345 4588 10349 4644
rect 10285 4584 10349 4588
rect 10365 4644 10429 4648
rect 10365 4588 10369 4644
rect 10369 4588 10425 4644
rect 10425 4588 10429 4644
rect 10365 4584 10429 4588
rect 10445 4644 10509 4648
rect 10445 4588 10449 4644
rect 10449 4588 10505 4644
rect 10505 4588 10509 4644
rect 10445 4584 10509 4588
rect 10525 4644 10589 4648
rect 10525 4588 10529 4644
rect 10529 4588 10585 4644
rect 10585 4588 10589 4644
rect 10525 4584 10589 4588
rect 19618 4644 19682 4648
rect 19618 4588 19622 4644
rect 19622 4588 19678 4644
rect 19678 4588 19682 4644
rect 19618 4584 19682 4588
rect 19698 4644 19762 4648
rect 19698 4588 19702 4644
rect 19702 4588 19758 4644
rect 19758 4588 19762 4644
rect 19698 4584 19762 4588
rect 19778 4644 19842 4648
rect 19778 4588 19782 4644
rect 19782 4588 19838 4644
rect 19838 4588 19842 4644
rect 19778 4584 19842 4588
rect 19858 4644 19922 4648
rect 19858 4588 19862 4644
rect 19862 4588 19918 4644
rect 19918 4588 19922 4644
rect 19858 4584 19922 4588
rect 5618 4100 5682 4104
rect 5618 4044 5622 4100
rect 5622 4044 5678 4100
rect 5678 4044 5682 4100
rect 5618 4040 5682 4044
rect 5698 4100 5762 4104
rect 5698 4044 5702 4100
rect 5702 4044 5758 4100
rect 5758 4044 5762 4100
rect 5698 4040 5762 4044
rect 5778 4100 5842 4104
rect 5778 4044 5782 4100
rect 5782 4044 5838 4100
rect 5838 4044 5842 4100
rect 5778 4040 5842 4044
rect 5858 4100 5922 4104
rect 5858 4044 5862 4100
rect 5862 4044 5918 4100
rect 5918 4044 5922 4100
rect 5858 4040 5922 4044
rect 14952 4100 15016 4104
rect 14952 4044 14956 4100
rect 14956 4044 15012 4100
rect 15012 4044 15016 4100
rect 14952 4040 15016 4044
rect 15032 4100 15096 4104
rect 15032 4044 15036 4100
rect 15036 4044 15092 4100
rect 15092 4044 15096 4100
rect 15032 4040 15096 4044
rect 15112 4100 15176 4104
rect 15112 4044 15116 4100
rect 15116 4044 15172 4100
rect 15172 4044 15176 4100
rect 15112 4040 15176 4044
rect 15192 4100 15256 4104
rect 15192 4044 15196 4100
rect 15196 4044 15252 4100
rect 15252 4044 15256 4100
rect 15192 4040 15256 4044
rect 24285 4100 24349 4104
rect 24285 4044 24289 4100
rect 24289 4044 24345 4100
rect 24345 4044 24349 4100
rect 24285 4040 24349 4044
rect 24365 4100 24429 4104
rect 24365 4044 24369 4100
rect 24369 4044 24425 4100
rect 24425 4044 24429 4100
rect 24365 4040 24429 4044
rect 24445 4100 24509 4104
rect 24445 4044 24449 4100
rect 24449 4044 24505 4100
rect 24505 4044 24509 4100
rect 24445 4040 24509 4044
rect 24525 4100 24589 4104
rect 24525 4044 24529 4100
rect 24529 4044 24585 4100
rect 24585 4044 24589 4100
rect 24525 4040 24589 4044
rect 10285 3556 10349 3560
rect 10285 3500 10289 3556
rect 10289 3500 10345 3556
rect 10345 3500 10349 3556
rect 10285 3496 10349 3500
rect 10365 3556 10429 3560
rect 10365 3500 10369 3556
rect 10369 3500 10425 3556
rect 10425 3500 10429 3556
rect 10365 3496 10429 3500
rect 10445 3556 10509 3560
rect 10445 3500 10449 3556
rect 10449 3500 10505 3556
rect 10505 3500 10509 3556
rect 10445 3496 10509 3500
rect 10525 3556 10589 3560
rect 10525 3500 10529 3556
rect 10529 3500 10585 3556
rect 10585 3500 10589 3556
rect 10525 3496 10589 3500
rect 19618 3556 19682 3560
rect 19618 3500 19622 3556
rect 19622 3500 19678 3556
rect 19678 3500 19682 3556
rect 19618 3496 19682 3500
rect 19698 3556 19762 3560
rect 19698 3500 19702 3556
rect 19702 3500 19758 3556
rect 19758 3500 19762 3556
rect 19698 3496 19762 3500
rect 19778 3556 19842 3560
rect 19778 3500 19782 3556
rect 19782 3500 19838 3556
rect 19838 3500 19842 3556
rect 19778 3496 19842 3500
rect 19858 3556 19922 3560
rect 19858 3500 19862 3556
rect 19862 3500 19918 3556
rect 19918 3500 19922 3556
rect 19858 3496 19922 3500
rect 5618 3012 5682 3016
rect 5618 2956 5622 3012
rect 5622 2956 5678 3012
rect 5678 2956 5682 3012
rect 5618 2952 5682 2956
rect 5698 3012 5762 3016
rect 5698 2956 5702 3012
rect 5702 2956 5758 3012
rect 5758 2956 5762 3012
rect 5698 2952 5762 2956
rect 5778 3012 5842 3016
rect 5778 2956 5782 3012
rect 5782 2956 5838 3012
rect 5838 2956 5842 3012
rect 5778 2952 5842 2956
rect 5858 3012 5922 3016
rect 5858 2956 5862 3012
rect 5862 2956 5918 3012
rect 5918 2956 5922 3012
rect 5858 2952 5922 2956
rect 14952 3012 15016 3016
rect 14952 2956 14956 3012
rect 14956 2956 15012 3012
rect 15012 2956 15016 3012
rect 14952 2952 15016 2956
rect 15032 3012 15096 3016
rect 15032 2956 15036 3012
rect 15036 2956 15092 3012
rect 15092 2956 15096 3012
rect 15032 2952 15096 2956
rect 15112 3012 15176 3016
rect 15112 2956 15116 3012
rect 15116 2956 15172 3012
rect 15172 2956 15176 3012
rect 15112 2952 15176 2956
rect 15192 3012 15256 3016
rect 15192 2956 15196 3012
rect 15196 2956 15252 3012
rect 15252 2956 15256 3012
rect 15192 2952 15256 2956
rect 24285 3012 24349 3016
rect 24285 2956 24289 3012
rect 24289 2956 24345 3012
rect 24345 2956 24349 3012
rect 24285 2952 24349 2956
rect 24365 3012 24429 3016
rect 24365 2956 24369 3012
rect 24369 2956 24425 3012
rect 24425 2956 24429 3012
rect 24365 2952 24429 2956
rect 24445 3012 24509 3016
rect 24445 2956 24449 3012
rect 24449 2956 24505 3012
rect 24505 2956 24509 3012
rect 24445 2952 24509 2956
rect 24525 3012 24589 3016
rect 24525 2956 24529 3012
rect 24529 2956 24585 3012
rect 24585 2956 24589 3012
rect 24525 2952 24589 2956
rect 10285 2468 10349 2472
rect 10285 2412 10289 2468
rect 10289 2412 10345 2468
rect 10345 2412 10349 2468
rect 10285 2408 10349 2412
rect 10365 2468 10429 2472
rect 10365 2412 10369 2468
rect 10369 2412 10425 2468
rect 10425 2412 10429 2468
rect 10365 2408 10429 2412
rect 10445 2468 10509 2472
rect 10445 2412 10449 2468
rect 10449 2412 10505 2468
rect 10505 2412 10509 2468
rect 10445 2408 10509 2412
rect 10525 2468 10589 2472
rect 10525 2412 10529 2468
rect 10529 2412 10585 2468
rect 10585 2412 10589 2468
rect 10525 2408 10589 2412
rect 19618 2468 19682 2472
rect 19618 2412 19622 2468
rect 19622 2412 19678 2468
rect 19678 2412 19682 2468
rect 19618 2408 19682 2412
rect 19698 2468 19762 2472
rect 19698 2412 19702 2468
rect 19702 2412 19758 2468
rect 19758 2412 19762 2468
rect 19698 2408 19762 2412
rect 19778 2468 19842 2472
rect 19778 2412 19782 2468
rect 19782 2412 19838 2468
rect 19838 2412 19842 2468
rect 19778 2408 19842 2412
rect 19858 2468 19922 2472
rect 19858 2412 19862 2468
rect 19862 2412 19918 2468
rect 19918 2412 19922 2468
rect 19858 2408 19922 2412
rect 5618 1924 5682 1928
rect 5618 1868 5622 1924
rect 5622 1868 5678 1924
rect 5678 1868 5682 1924
rect 5618 1864 5682 1868
rect 5698 1924 5762 1928
rect 5698 1868 5702 1924
rect 5702 1868 5758 1924
rect 5758 1868 5762 1924
rect 5698 1864 5762 1868
rect 5778 1924 5842 1928
rect 5778 1868 5782 1924
rect 5782 1868 5838 1924
rect 5838 1868 5842 1924
rect 5778 1864 5842 1868
rect 5858 1924 5922 1928
rect 5858 1868 5862 1924
rect 5862 1868 5918 1924
rect 5918 1868 5922 1924
rect 5858 1864 5922 1868
rect 14952 1924 15016 1928
rect 14952 1868 14956 1924
rect 14956 1868 15012 1924
rect 15012 1868 15016 1924
rect 14952 1864 15016 1868
rect 15032 1924 15096 1928
rect 15032 1868 15036 1924
rect 15036 1868 15092 1924
rect 15092 1868 15096 1924
rect 15032 1864 15096 1868
rect 15112 1924 15176 1928
rect 15112 1868 15116 1924
rect 15116 1868 15172 1924
rect 15172 1868 15176 1924
rect 15112 1864 15176 1868
rect 15192 1924 15256 1928
rect 15192 1868 15196 1924
rect 15196 1868 15252 1924
rect 15252 1868 15256 1924
rect 15192 1864 15256 1868
rect 24285 1924 24349 1928
rect 24285 1868 24289 1924
rect 24289 1868 24345 1924
rect 24345 1868 24349 1924
rect 24285 1864 24349 1868
rect 24365 1924 24429 1928
rect 24365 1868 24369 1924
rect 24369 1868 24425 1924
rect 24425 1868 24429 1924
rect 24365 1864 24429 1868
rect 24445 1924 24509 1928
rect 24445 1868 24449 1924
rect 24449 1868 24505 1924
rect 24505 1868 24509 1924
rect 24445 1864 24509 1868
rect 24525 1924 24589 1928
rect 24525 1868 24529 1924
rect 24529 1868 24585 1924
rect 24585 1868 24589 1924
rect 24525 1864 24589 1868
<< metal4 >>
rect 5610 24776 5931 25336
rect 5610 24712 5618 24776
rect 5682 24712 5698 24776
rect 5762 24712 5778 24776
rect 5842 24712 5858 24776
rect 5922 24712 5931 24776
rect 5610 23688 5931 24712
rect 5610 23624 5618 23688
rect 5682 23624 5698 23688
rect 5762 23624 5778 23688
rect 5842 23624 5858 23688
rect 5922 23624 5931 23688
rect 5610 22600 5931 23624
rect 5610 22536 5618 22600
rect 5682 22536 5698 22600
rect 5762 22536 5778 22600
rect 5842 22536 5858 22600
rect 5922 22536 5931 22600
rect 5610 21512 5931 22536
rect 5610 21448 5618 21512
rect 5682 21448 5698 21512
rect 5762 21448 5778 21512
rect 5842 21448 5858 21512
rect 5922 21448 5931 21512
rect 5610 20424 5931 21448
rect 5610 20360 5618 20424
rect 5682 20360 5698 20424
rect 5762 20360 5778 20424
rect 5842 20360 5858 20424
rect 5922 20360 5931 20424
rect 5610 19336 5931 20360
rect 5610 19272 5618 19336
rect 5682 19272 5698 19336
rect 5762 19272 5778 19336
rect 5842 19272 5858 19336
rect 5922 19272 5931 19336
rect 5610 18248 5931 19272
rect 5610 18184 5618 18248
rect 5682 18184 5698 18248
rect 5762 18184 5778 18248
rect 5842 18184 5858 18248
rect 5922 18184 5931 18248
rect 5610 17160 5931 18184
rect 5610 17096 5618 17160
rect 5682 17096 5698 17160
rect 5762 17096 5778 17160
rect 5842 17096 5858 17160
rect 5922 17096 5931 17160
rect 5610 16072 5931 17096
rect 5610 16008 5618 16072
rect 5682 16008 5698 16072
rect 5762 16008 5778 16072
rect 5842 16008 5858 16072
rect 5922 16008 5931 16072
rect 5610 14984 5931 16008
rect 5610 14920 5618 14984
rect 5682 14920 5698 14984
rect 5762 14920 5778 14984
rect 5842 14920 5858 14984
rect 5922 14920 5931 14984
rect 5610 13896 5931 14920
rect 5610 13832 5618 13896
rect 5682 13832 5698 13896
rect 5762 13832 5778 13896
rect 5842 13832 5858 13896
rect 5922 13832 5931 13896
rect 5610 12808 5931 13832
rect 5610 12744 5618 12808
rect 5682 12744 5698 12808
rect 5762 12744 5778 12808
rect 5842 12744 5858 12808
rect 5922 12744 5931 12808
rect 5610 11720 5931 12744
rect 5610 11656 5618 11720
rect 5682 11656 5698 11720
rect 5762 11656 5778 11720
rect 5842 11656 5858 11720
rect 5922 11656 5931 11720
rect 5610 10632 5931 11656
rect 5610 10568 5618 10632
rect 5682 10568 5698 10632
rect 5762 10568 5778 10632
rect 5842 10568 5858 10632
rect 5922 10568 5931 10632
rect 5610 9544 5931 10568
rect 5610 9480 5618 9544
rect 5682 9480 5698 9544
rect 5762 9480 5778 9544
rect 5842 9480 5858 9544
rect 5922 9480 5931 9544
rect 5610 8456 5931 9480
rect 5610 8392 5618 8456
rect 5682 8392 5698 8456
rect 5762 8392 5778 8456
rect 5842 8392 5858 8456
rect 5922 8392 5931 8456
rect 5610 7368 5931 8392
rect 5610 7304 5618 7368
rect 5682 7304 5698 7368
rect 5762 7304 5778 7368
rect 5842 7304 5858 7368
rect 5922 7304 5931 7368
rect 5610 6280 5931 7304
rect 5610 6216 5618 6280
rect 5682 6216 5698 6280
rect 5762 6216 5778 6280
rect 5842 6216 5858 6280
rect 5922 6216 5931 6280
rect 5610 5192 5931 6216
rect 5610 5128 5618 5192
rect 5682 5128 5698 5192
rect 5762 5128 5778 5192
rect 5842 5128 5858 5192
rect 5922 5128 5931 5192
rect 5610 4104 5931 5128
rect 5610 4040 5618 4104
rect 5682 4040 5698 4104
rect 5762 4040 5778 4104
rect 5842 4040 5858 4104
rect 5922 4040 5931 4104
rect 5610 3016 5931 4040
rect 5610 2952 5618 3016
rect 5682 2952 5698 3016
rect 5762 2952 5778 3016
rect 5842 2952 5858 3016
rect 5922 2952 5931 3016
rect 5610 1928 5931 2952
rect 5610 1864 5618 1928
rect 5682 1864 5698 1928
rect 5762 1864 5778 1928
rect 5842 1864 5858 1928
rect 5922 1864 5931 1928
rect 5610 1848 5931 1864
rect 10277 25320 10597 25336
rect 10277 25256 10285 25320
rect 10349 25256 10365 25320
rect 10429 25256 10445 25320
rect 10509 25256 10525 25320
rect 10589 25256 10597 25320
rect 10277 24232 10597 25256
rect 10277 24168 10285 24232
rect 10349 24168 10365 24232
rect 10429 24168 10445 24232
rect 10509 24168 10525 24232
rect 10589 24168 10597 24232
rect 10277 23144 10597 24168
rect 10277 23080 10285 23144
rect 10349 23080 10365 23144
rect 10429 23080 10445 23144
rect 10509 23080 10525 23144
rect 10589 23080 10597 23144
rect 10277 22056 10597 23080
rect 10277 21992 10285 22056
rect 10349 21992 10365 22056
rect 10429 21992 10445 22056
rect 10509 21992 10525 22056
rect 10589 21992 10597 22056
rect 10277 20968 10597 21992
rect 10277 20904 10285 20968
rect 10349 20904 10365 20968
rect 10429 20904 10445 20968
rect 10509 20904 10525 20968
rect 10589 20904 10597 20968
rect 10277 19880 10597 20904
rect 10277 19816 10285 19880
rect 10349 19816 10365 19880
rect 10429 19816 10445 19880
rect 10509 19816 10525 19880
rect 10589 19816 10597 19880
rect 10277 18792 10597 19816
rect 10277 18728 10285 18792
rect 10349 18728 10365 18792
rect 10429 18728 10445 18792
rect 10509 18728 10525 18792
rect 10589 18728 10597 18792
rect 10277 17704 10597 18728
rect 10277 17640 10285 17704
rect 10349 17640 10365 17704
rect 10429 17640 10445 17704
rect 10509 17640 10525 17704
rect 10589 17640 10597 17704
rect 10277 16616 10597 17640
rect 10277 16552 10285 16616
rect 10349 16552 10365 16616
rect 10429 16552 10445 16616
rect 10509 16552 10525 16616
rect 10589 16552 10597 16616
rect 10277 15528 10597 16552
rect 10277 15464 10285 15528
rect 10349 15464 10365 15528
rect 10429 15464 10445 15528
rect 10509 15464 10525 15528
rect 10589 15464 10597 15528
rect 10277 14440 10597 15464
rect 10277 14376 10285 14440
rect 10349 14376 10365 14440
rect 10429 14376 10445 14440
rect 10509 14376 10525 14440
rect 10589 14376 10597 14440
rect 10277 13352 10597 14376
rect 10277 13288 10285 13352
rect 10349 13288 10365 13352
rect 10429 13288 10445 13352
rect 10509 13288 10525 13352
rect 10589 13288 10597 13352
rect 10277 12264 10597 13288
rect 10277 12200 10285 12264
rect 10349 12200 10365 12264
rect 10429 12200 10445 12264
rect 10509 12200 10525 12264
rect 10589 12200 10597 12264
rect 10277 11176 10597 12200
rect 10277 11112 10285 11176
rect 10349 11112 10365 11176
rect 10429 11112 10445 11176
rect 10509 11112 10525 11176
rect 10589 11112 10597 11176
rect 10277 10088 10597 11112
rect 10277 10024 10285 10088
rect 10349 10024 10365 10088
rect 10429 10024 10445 10088
rect 10509 10024 10525 10088
rect 10589 10024 10597 10088
rect 10277 9000 10597 10024
rect 10277 8936 10285 9000
rect 10349 8936 10365 9000
rect 10429 8936 10445 9000
rect 10509 8936 10525 9000
rect 10589 8936 10597 9000
rect 10277 7912 10597 8936
rect 10277 7848 10285 7912
rect 10349 7848 10365 7912
rect 10429 7848 10445 7912
rect 10509 7848 10525 7912
rect 10589 7848 10597 7912
rect 10277 6824 10597 7848
rect 10277 6760 10285 6824
rect 10349 6760 10365 6824
rect 10429 6760 10445 6824
rect 10509 6760 10525 6824
rect 10589 6760 10597 6824
rect 10277 5736 10597 6760
rect 10277 5672 10285 5736
rect 10349 5672 10365 5736
rect 10429 5672 10445 5736
rect 10509 5672 10525 5736
rect 10589 5672 10597 5736
rect 10277 4648 10597 5672
rect 10277 4584 10285 4648
rect 10349 4584 10365 4648
rect 10429 4584 10445 4648
rect 10509 4584 10525 4648
rect 10589 4584 10597 4648
rect 10277 3560 10597 4584
rect 10277 3496 10285 3560
rect 10349 3496 10365 3560
rect 10429 3496 10445 3560
rect 10509 3496 10525 3560
rect 10589 3496 10597 3560
rect 10277 2472 10597 3496
rect 10277 2408 10285 2472
rect 10349 2408 10365 2472
rect 10429 2408 10445 2472
rect 10509 2408 10525 2472
rect 10589 2408 10597 2472
rect 10277 1848 10597 2408
rect 14944 24776 15264 25336
rect 14944 24712 14952 24776
rect 15016 24712 15032 24776
rect 15096 24712 15112 24776
rect 15176 24712 15192 24776
rect 15256 24712 15264 24776
rect 14944 23688 15264 24712
rect 14944 23624 14952 23688
rect 15016 23624 15032 23688
rect 15096 23624 15112 23688
rect 15176 23624 15192 23688
rect 15256 23624 15264 23688
rect 14944 22600 15264 23624
rect 14944 22536 14952 22600
rect 15016 22536 15032 22600
rect 15096 22536 15112 22600
rect 15176 22536 15192 22600
rect 15256 22536 15264 22600
rect 14944 21512 15264 22536
rect 14944 21448 14952 21512
rect 15016 21448 15032 21512
rect 15096 21448 15112 21512
rect 15176 21448 15192 21512
rect 15256 21448 15264 21512
rect 14944 20424 15264 21448
rect 14944 20360 14952 20424
rect 15016 20360 15032 20424
rect 15096 20360 15112 20424
rect 15176 20360 15192 20424
rect 15256 20360 15264 20424
rect 14944 19336 15264 20360
rect 14944 19272 14952 19336
rect 15016 19272 15032 19336
rect 15096 19272 15112 19336
rect 15176 19272 15192 19336
rect 15256 19272 15264 19336
rect 14944 18248 15264 19272
rect 14944 18184 14952 18248
rect 15016 18184 15032 18248
rect 15096 18184 15112 18248
rect 15176 18184 15192 18248
rect 15256 18184 15264 18248
rect 14944 17160 15264 18184
rect 14944 17096 14952 17160
rect 15016 17096 15032 17160
rect 15096 17096 15112 17160
rect 15176 17096 15192 17160
rect 15256 17096 15264 17160
rect 14944 16072 15264 17096
rect 14944 16008 14952 16072
rect 15016 16008 15032 16072
rect 15096 16008 15112 16072
rect 15176 16008 15192 16072
rect 15256 16008 15264 16072
rect 14944 14984 15264 16008
rect 14944 14920 14952 14984
rect 15016 14920 15032 14984
rect 15096 14920 15112 14984
rect 15176 14920 15192 14984
rect 15256 14920 15264 14984
rect 14944 13896 15264 14920
rect 14944 13832 14952 13896
rect 15016 13832 15032 13896
rect 15096 13832 15112 13896
rect 15176 13832 15192 13896
rect 15256 13832 15264 13896
rect 14944 12808 15264 13832
rect 14944 12744 14952 12808
rect 15016 12744 15032 12808
rect 15096 12744 15112 12808
rect 15176 12744 15192 12808
rect 15256 12744 15264 12808
rect 14944 11720 15264 12744
rect 14944 11656 14952 11720
rect 15016 11656 15032 11720
rect 15096 11656 15112 11720
rect 15176 11656 15192 11720
rect 15256 11656 15264 11720
rect 14944 10632 15264 11656
rect 14944 10568 14952 10632
rect 15016 10568 15032 10632
rect 15096 10568 15112 10632
rect 15176 10568 15192 10632
rect 15256 10568 15264 10632
rect 14944 9544 15264 10568
rect 14944 9480 14952 9544
rect 15016 9480 15032 9544
rect 15096 9480 15112 9544
rect 15176 9480 15192 9544
rect 15256 9480 15264 9544
rect 14944 8456 15264 9480
rect 14944 8392 14952 8456
rect 15016 8392 15032 8456
rect 15096 8392 15112 8456
rect 15176 8392 15192 8456
rect 15256 8392 15264 8456
rect 14944 7368 15264 8392
rect 14944 7304 14952 7368
rect 15016 7304 15032 7368
rect 15096 7304 15112 7368
rect 15176 7304 15192 7368
rect 15256 7304 15264 7368
rect 14944 6280 15264 7304
rect 14944 6216 14952 6280
rect 15016 6216 15032 6280
rect 15096 6216 15112 6280
rect 15176 6216 15192 6280
rect 15256 6216 15264 6280
rect 14944 5192 15264 6216
rect 14944 5128 14952 5192
rect 15016 5128 15032 5192
rect 15096 5128 15112 5192
rect 15176 5128 15192 5192
rect 15256 5128 15264 5192
rect 14944 4104 15264 5128
rect 14944 4040 14952 4104
rect 15016 4040 15032 4104
rect 15096 4040 15112 4104
rect 15176 4040 15192 4104
rect 15256 4040 15264 4104
rect 14944 3016 15264 4040
rect 14944 2952 14952 3016
rect 15016 2952 15032 3016
rect 15096 2952 15112 3016
rect 15176 2952 15192 3016
rect 15256 2952 15264 3016
rect 14944 1928 15264 2952
rect 14944 1864 14952 1928
rect 15016 1864 15032 1928
rect 15096 1864 15112 1928
rect 15176 1864 15192 1928
rect 15256 1864 15264 1928
rect 14944 1848 15264 1864
rect 19610 25320 19930 25336
rect 19610 25256 19618 25320
rect 19682 25256 19698 25320
rect 19762 25256 19778 25320
rect 19842 25256 19858 25320
rect 19922 25256 19930 25320
rect 19610 24232 19930 25256
rect 19610 24168 19618 24232
rect 19682 24168 19698 24232
rect 19762 24168 19778 24232
rect 19842 24168 19858 24232
rect 19922 24168 19930 24232
rect 19610 23144 19930 24168
rect 19610 23080 19618 23144
rect 19682 23080 19698 23144
rect 19762 23080 19778 23144
rect 19842 23080 19858 23144
rect 19922 23080 19930 23144
rect 19610 22056 19930 23080
rect 19610 21992 19618 22056
rect 19682 21992 19698 22056
rect 19762 21992 19778 22056
rect 19842 21992 19858 22056
rect 19922 21992 19930 22056
rect 19610 20968 19930 21992
rect 19610 20904 19618 20968
rect 19682 20904 19698 20968
rect 19762 20904 19778 20968
rect 19842 20904 19858 20968
rect 19922 20904 19930 20968
rect 19610 19880 19930 20904
rect 19610 19816 19618 19880
rect 19682 19816 19698 19880
rect 19762 19816 19778 19880
rect 19842 19816 19858 19880
rect 19922 19816 19930 19880
rect 19610 18792 19930 19816
rect 19610 18728 19618 18792
rect 19682 18728 19698 18792
rect 19762 18728 19778 18792
rect 19842 18728 19858 18792
rect 19922 18728 19930 18792
rect 19610 17704 19930 18728
rect 19610 17640 19618 17704
rect 19682 17640 19698 17704
rect 19762 17640 19778 17704
rect 19842 17640 19858 17704
rect 19922 17640 19930 17704
rect 19610 16616 19930 17640
rect 19610 16552 19618 16616
rect 19682 16552 19698 16616
rect 19762 16552 19778 16616
rect 19842 16552 19858 16616
rect 19922 16552 19930 16616
rect 19610 15528 19930 16552
rect 19610 15464 19618 15528
rect 19682 15464 19698 15528
rect 19762 15464 19778 15528
rect 19842 15464 19858 15528
rect 19922 15464 19930 15528
rect 19610 14440 19930 15464
rect 19610 14376 19618 14440
rect 19682 14376 19698 14440
rect 19762 14376 19778 14440
rect 19842 14376 19858 14440
rect 19922 14376 19930 14440
rect 19610 13352 19930 14376
rect 19610 13288 19618 13352
rect 19682 13288 19698 13352
rect 19762 13288 19778 13352
rect 19842 13288 19858 13352
rect 19922 13288 19930 13352
rect 19610 12264 19930 13288
rect 19610 12200 19618 12264
rect 19682 12200 19698 12264
rect 19762 12200 19778 12264
rect 19842 12200 19858 12264
rect 19922 12200 19930 12264
rect 19610 11176 19930 12200
rect 19610 11112 19618 11176
rect 19682 11112 19698 11176
rect 19762 11112 19778 11176
rect 19842 11112 19858 11176
rect 19922 11112 19930 11176
rect 19610 10088 19930 11112
rect 19610 10024 19618 10088
rect 19682 10024 19698 10088
rect 19762 10024 19778 10088
rect 19842 10024 19858 10088
rect 19922 10024 19930 10088
rect 19610 9000 19930 10024
rect 19610 8936 19618 9000
rect 19682 8936 19698 9000
rect 19762 8936 19778 9000
rect 19842 8936 19858 9000
rect 19922 8936 19930 9000
rect 19610 7912 19930 8936
rect 19610 7848 19618 7912
rect 19682 7848 19698 7912
rect 19762 7848 19778 7912
rect 19842 7848 19858 7912
rect 19922 7848 19930 7912
rect 19610 6824 19930 7848
rect 19610 6760 19618 6824
rect 19682 6760 19698 6824
rect 19762 6760 19778 6824
rect 19842 6760 19858 6824
rect 19922 6760 19930 6824
rect 19610 5736 19930 6760
rect 19610 5672 19618 5736
rect 19682 5672 19698 5736
rect 19762 5672 19778 5736
rect 19842 5672 19858 5736
rect 19922 5672 19930 5736
rect 19610 4648 19930 5672
rect 19610 4584 19618 4648
rect 19682 4584 19698 4648
rect 19762 4584 19778 4648
rect 19842 4584 19858 4648
rect 19922 4584 19930 4648
rect 19610 3560 19930 4584
rect 19610 3496 19618 3560
rect 19682 3496 19698 3560
rect 19762 3496 19778 3560
rect 19842 3496 19858 3560
rect 19922 3496 19930 3560
rect 19610 2472 19930 3496
rect 19610 2408 19618 2472
rect 19682 2408 19698 2472
rect 19762 2408 19778 2472
rect 19842 2408 19858 2472
rect 19922 2408 19930 2472
rect 19610 1848 19930 2408
rect 24277 24776 24597 25336
rect 24277 24712 24285 24776
rect 24349 24712 24365 24776
rect 24429 24712 24445 24776
rect 24509 24712 24525 24776
rect 24589 24712 24597 24776
rect 24277 23688 24597 24712
rect 24277 23624 24285 23688
rect 24349 23624 24365 23688
rect 24429 23624 24445 23688
rect 24509 23624 24525 23688
rect 24589 23624 24597 23688
rect 24277 22600 24597 23624
rect 24277 22536 24285 22600
rect 24349 22536 24365 22600
rect 24429 22536 24445 22600
rect 24509 22536 24525 22600
rect 24589 22536 24597 22600
rect 24277 21512 24597 22536
rect 24277 21448 24285 21512
rect 24349 21448 24365 21512
rect 24429 21448 24445 21512
rect 24509 21448 24525 21512
rect 24589 21448 24597 21512
rect 24277 20424 24597 21448
rect 24277 20360 24285 20424
rect 24349 20360 24365 20424
rect 24429 20360 24445 20424
rect 24509 20360 24525 20424
rect 24589 20360 24597 20424
rect 24277 19336 24597 20360
rect 24277 19272 24285 19336
rect 24349 19272 24365 19336
rect 24429 19272 24445 19336
rect 24509 19272 24525 19336
rect 24589 19272 24597 19336
rect 24277 18248 24597 19272
rect 24277 18184 24285 18248
rect 24349 18184 24365 18248
rect 24429 18184 24445 18248
rect 24509 18184 24525 18248
rect 24589 18184 24597 18248
rect 24277 17160 24597 18184
rect 24277 17096 24285 17160
rect 24349 17096 24365 17160
rect 24429 17096 24445 17160
rect 24509 17096 24525 17160
rect 24589 17096 24597 17160
rect 24277 16072 24597 17096
rect 24277 16008 24285 16072
rect 24349 16008 24365 16072
rect 24429 16008 24445 16072
rect 24509 16008 24525 16072
rect 24589 16008 24597 16072
rect 24277 14984 24597 16008
rect 24277 14920 24285 14984
rect 24349 14920 24365 14984
rect 24429 14920 24445 14984
rect 24509 14920 24525 14984
rect 24589 14920 24597 14984
rect 24277 13896 24597 14920
rect 24277 13832 24285 13896
rect 24349 13832 24365 13896
rect 24429 13832 24445 13896
rect 24509 13832 24525 13896
rect 24589 13832 24597 13896
rect 24277 12808 24597 13832
rect 24277 12744 24285 12808
rect 24349 12744 24365 12808
rect 24429 12744 24445 12808
rect 24509 12744 24525 12808
rect 24589 12744 24597 12808
rect 24277 11720 24597 12744
rect 24277 11656 24285 11720
rect 24349 11656 24365 11720
rect 24429 11656 24445 11720
rect 24509 11656 24525 11720
rect 24589 11656 24597 11720
rect 24277 10632 24597 11656
rect 24277 10568 24285 10632
rect 24349 10568 24365 10632
rect 24429 10568 24445 10632
rect 24509 10568 24525 10632
rect 24589 10568 24597 10632
rect 24277 9544 24597 10568
rect 24277 9480 24285 9544
rect 24349 9480 24365 9544
rect 24429 9480 24445 9544
rect 24509 9480 24525 9544
rect 24589 9480 24597 9544
rect 24277 8456 24597 9480
rect 24277 8392 24285 8456
rect 24349 8392 24365 8456
rect 24429 8392 24445 8456
rect 24509 8392 24525 8456
rect 24589 8392 24597 8456
rect 24277 7368 24597 8392
rect 24277 7304 24285 7368
rect 24349 7304 24365 7368
rect 24429 7304 24445 7368
rect 24509 7304 24525 7368
rect 24589 7304 24597 7368
rect 24277 6280 24597 7304
rect 24277 6216 24285 6280
rect 24349 6216 24365 6280
rect 24429 6216 24445 6280
rect 24509 6216 24525 6280
rect 24589 6216 24597 6280
rect 24277 5192 24597 6216
rect 24277 5128 24285 5192
rect 24349 5128 24365 5192
rect 24429 5128 24445 5192
rect 24509 5128 24525 5192
rect 24589 5128 24597 5192
rect 24277 4104 24597 5128
rect 24277 4040 24285 4104
rect 24349 4040 24365 4104
rect 24429 4040 24445 4104
rect 24509 4040 24525 4104
rect 24589 4040 24597 4104
rect 24277 3016 24597 4040
rect 24277 2952 24285 3016
rect 24349 2952 24365 3016
rect 24429 2952 24445 3016
rect 24509 2952 24525 3016
rect 24589 2952 24597 3016
rect 24277 1928 24597 2952
rect 24277 1864 24285 1928
rect 24349 1864 24365 1928
rect 24429 1864 24445 1928
rect 24509 1864 24525 1928
rect 24589 1864 24597 1928
rect 24277 1848 24597 1864
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1604681595
transform 1 0 4048 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1604681595
transform 1 0 5152 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1604681595
transform 1 0 6256 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1604681595
transform 1 0 7360 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1604681595
transform 1 0 8464 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1604681595
transform 1 0 9660 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1604681595
transform 1 0 10764 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1604681595
transform 1 0 12972 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1604681595
transform 1 0 14076 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1604681595
transform 1 0 16376 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1604681595
transform 1 0 19688 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_215
timestamp 1604681595
transform 1 0 20884 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_239
timestamp 1604681595
transform 1 0 23092 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_263
timestamp 1604681595
transform 1 0 25300 0 1 2440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 1 2440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1604681595
transform 1 0 4692 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 -1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1604681595
transform 1 0 6808 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1604681595
transform 1 0 7912 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1604681595
transform 1 0 9016 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1604681595
transform 1 0 10120 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1604681595
transform 1 0 11224 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1604681595
transform 1 0 12420 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1604681595
transform 1 0 13524 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1604681595
transform 1 0 14628 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1604681595
transform 1 0 15732 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1604681595
transform 1 0 19136 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_220
timestamp 1604681595
transform 1 0 21344 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_232
timestamp 1604681595
transform 1 0 22448 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 -1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_245
timestamp 1604681595
transform 1 0 23644 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_257
timestamp 1604681595
transform 1 0 24748 0 -1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_269
timestamp 1604681595
transform 1 0 25852 0 -1 3528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1604681595
transform 1 0 4048 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1604681595
transform 1 0 5152 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1604681595
transform 1 0 6256 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1604681595
transform 1 0 7360 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1604681595
transform 1 0 8464 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1604681595
transform 1 0 9660 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1604681595
transform 1 0 10764 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1604681595
transform 1 0 12972 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1604681595
transform 1 0 14076 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1604681595
transform 1 0 15272 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1604681595
transform 1 0 16376 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1604681595
transform 1 0 17480 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1604681595
transform 1 0 18584 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1604681595
transform 1 0 19688 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_227
timestamp 1604681595
transform 1 0 21988 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_239
timestamp 1604681595
transform 1 0 23092 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1604681595
transform 1 0 24196 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 1 3528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25116 0 1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_259
timestamp 1604681595
transform 1 0 24932 0 1 3528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_263
timestamp 1604681595
transform 1 0 25300 0 1 3528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1604681595
transform 1 0 4692 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1604681595
transform 1 0 5796 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1604681595
transform 1 0 6532 0 -1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1604681595
transform 1 0 13524 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1604681595
transform 1 0 14628 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1604681595
transform 1 0 15732 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1604681595
transform 1 0 16836 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1604681595
transform 1 0 18032 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1604681595
transform 1 0 19136 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1604681595
transform 1 0 20240 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_220
timestamp 1604681595
transform 1 0 21344 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_232
timestamp 1604681595
transform 1 0 22448 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 -1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1604681595
transform 1 0 23644 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_257
timestamp 1604681595
transform 1 0 24748 0 -1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_269
timestamp 1604681595
transform 1 0 25852 0 -1 4616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1604681595
transform 1 0 4048 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1604681595
transform 1 0 7360 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1604681595
transform 1 0 8464 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1604681595
transform 1 0 9660 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1604681595
transform 1 0 10764 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1604681595
transform 1 0 11868 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 15272 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 15824 0 1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_162
timestamp 1604681595
transform 1 0 16008 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_174
timestamp 1604681595
transform 1 0 17112 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_186
timestamp 1604681595
transform 1 0 18216 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_198
timestamp 1604681595
transform 1 0 19320 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_227
timestamp 1604681595
transform 1 0 21988 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_239
timestamp 1604681595
transform 1 0 23092 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_251
timestamp 1604681595
transform 1 0 24196 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_263
timestamp 1604681595
transform 1 0 25300 0 1 4616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1604681595
transform 1 0 4048 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1604681595
transform 1 0 4692 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1604681595
transform 1 0 5152 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1604681595
transform 1 0 5796 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1604681595
transform 1 0 6532 0 -1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1604681595
transform 1 0 6808 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1604681595
transform 1 0 7912 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1604681595
transform 1 0 7360 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1604681595
transform 1 0 8464 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1604681595
transform 1 0 9016 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1604681595
transform 1 0 9660 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1604681595
transform 1 0 12420 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1604681595
transform 1 0 12972 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1604681595
transform 1 0 14628 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1604681595
transform 1 0 14076 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 16192 0 1 5704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1604681595
transform 1 0 15732 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_154
timestamp 1604681595
transform 1 0 15272 0 1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_168
timestamp 1604681595
transform 1 0 16560 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 16744 0 1 5704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1604681595
transform 1 0 16836 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1604681595
transform 1 0 18032 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1604681595
transform 1 0 16928 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1604681595
transform 1 0 19136 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1604681595
transform 1 0 20240 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_220
timestamp 1604681595
transform 1 0 21344 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_232
timestamp 1604681595
transform 1 0 22448 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_227
timestamp 1604681595
transform 1 0 21988 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 -1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_245
timestamp 1604681595
transform 1 0 23644 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_239
timestamp 1604681595
transform 1 0 23092 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_251
timestamp 1604681595
transform 1 0 24196 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_257
timestamp 1604681595
transform 1 0 24748 0 -1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_269
timestamp 1604681595
transform 1 0 25852 0 -1 5704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_263
timestamp 1604681595
transform 1 0 25300 0 1 5704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1604681595
transform 1 0 5796 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1604681595
transform 1 0 7912 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_86
timestamp 1604681595
transform 1 0 9016 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_98
timestamp 1604681595
transform 1 0 10120 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_110
timestamp 1604681595
transform 1 0 11224 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_147
timestamp 1604681595
transform 1 0 14628 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_159
timestamp 1604681595
transform 1 0 15732 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_171
timestamp 1604681595
transform 1 0 16836 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1604681595
transform 1 0 20240 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_220
timestamp 1604681595
transform 1 0 21344 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_232
timestamp 1604681595
transform 1 0 22448 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 -1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_245
timestamp 1604681595
transform 1 0 23644 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1604681595
transform 1 0 24748 0 -1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_269
timestamp 1604681595
transform 1 0 25852 0 -1 6792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1604681595
transform 1 0 4048 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1604681595
transform 1 0 5152 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1604681595
transform 1 0 6256 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1604681595
transform 1 0 8464 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1604681595
transform 1 0 9660 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_105
timestamp 1604681595
transform 1 0 10764 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_117
timestamp 1604681595
transform 1 0 11868 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_129
timestamp 1604681595
transform 1 0 12972 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1604681595
transform 1 0 14076 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 17572 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 18124 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_183
timestamp 1604681595
transform 1 0 17940 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_187
timestamp 1604681595
transform 1 0 18308 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_199
timestamp 1604681595
transform 1 0 19412 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp 1604681595
transform 1 0 20516 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_227
timestamp 1604681595
transform 1 0 21988 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_239
timestamp 1604681595
transform 1 0 23092 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_251
timestamp 1604681595
transform 1 0 24196 0 1 6792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 24564 0 1 6792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 6792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 6792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 6792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 6792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1604681595
transform 1 0 4692 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1604681595
transform 1 0 5796 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1604681595
transform 1 0 6532 0 -1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_98
timestamp 1604681595
transform 1 0 10120 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1604681595
transform 1 0 12420 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1604681595
transform 1 0 13524 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_159
timestamp 1604681595
transform 1 0 15732 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_171
timestamp 1604681595
transform 1 0 16836 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1604681595
transform 1 0 19136 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_208
timestamp 1604681595
transform 1 0 20240 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1604681595
transform 1 0 21344 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_232
timestamp 1604681595
transform 1 0 22448 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 -1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_245
timestamp 1604681595
transform 1 0 23644 0 -1 7880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 24564 0 -1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1604681595
transform 1 0 24380 0 -1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_259
timestamp 1604681595
transform 1 0 24932 0 -1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_271
timestamp 1604681595
transform 1 0 26036 0 -1 7880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1604681595
transform 1 0 5152 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1604681595
transform 1 0 7360 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1604681595
transform 1 0 8464 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1604681595
transform 1 0 10764 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_129
timestamp 1604681595
transform 1 0 12972 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_141
timestamp 1604681595
transform 1 0 14076 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1604681595
transform 1 0 16376 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_190
timestamp 1604681595
transform 1 0 18584 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_239
timestamp 1604681595
transform 1 0 23092 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1604681595
transform 1 0 24196 0 1 7880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 24564 0 1 7880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 7880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 7880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 7880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 7880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1604681595
transform 1 0 4692 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1604681595
transform 1 0 5796 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1604681595
transform 1 0 6808 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1604681595
transform 1 0 7912 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1604681595
transform 1 0 9016 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1604681595
transform 1 0 10120 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1604681595
transform 1 0 12420 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_147
timestamp 1604681595
transform 1 0 14628 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_159
timestamp 1604681595
transform 1 0 15732 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1604681595
transform 1 0 16836 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1604681595
transform 1 0 19136 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_208
timestamp 1604681595
transform 1 0 20240 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_220
timestamp 1604681595
transform 1 0 21344 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_232
timestamp 1604681595
transform 1 0 22448 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 -1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_245
timestamp 1604681595
transform 1 0 23644 0 -1 8968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 24564 0 -1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1604681595
transform 1 0 24380 0 -1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1604681595
transform 1 0 24932 0 -1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 8968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1604681595
transform 1 0 4048 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1604681595
transform 1 0 5152 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1604681595
transform 1 0 4692 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1604681595
transform 1 0 5796 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1604681595
transform 1 0 6532 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1604681595
transform 1 0 8464 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1604681595
transform 1 0 9660 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_98
timestamp 1604681595
transform 1 0 10120 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_117
timestamp 1604681595
transform 1 0 11868 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_110
timestamp 1604681595
transform 1 0 11224 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1604681595
transform 1 0 12420 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_141
timestamp 1604681595
transform 1 0 14076 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_147
timestamp 1604681595
transform 1 0 14628 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1604681595
transform 1 0 15272 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1604681595
transform 1 0 16376 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_159
timestamp 1604681595
transform 1 0 15732 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_178
timestamp 1604681595
transform 1 0 17480 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_171
timestamp 1604681595
transform 1 0 16836 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1604681595
transform 1 0 18584 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_196
timestamp 1604681595
transform 1 0 19136 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_208
timestamp 1604681595
transform 1 0 20240 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1604681595
transform 1 0 21988 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_220
timestamp 1604681595
transform 1 0 21344 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 -1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_239
timestamp 1604681595
transform 1 0 23092 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_251
timestamp 1604681595
transform 1 0 24196 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_245
timestamp 1604681595
transform 1 0 23644 0 -1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 24564 0 -1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 24564 0 1 8968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 25116 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 24380 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604681595
transform 1 0 24932 0 1 8968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_263
timestamp 1604681595
transform 1 0 25300 0 1 8968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1604681595
transform 1 0 24380 0 -1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 8968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604681595
transform 1 0 26496 0 1 8968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_68
timestamp 1604681595
transform 1 0 7360 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_80
timestamp 1604681595
transform 1 0 8464 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1604681595
transform 1 0 10764 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1604681595
transform 1 0 15088 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_154
timestamp 1604681595
transform 1 0 15272 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_191
timestamp 1604681595
transform 1 0 18676 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_203
timestamp 1604681595
transform 1 0 19780 0 1 10056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_227
timestamp 1604681595
transform 1 0 21988 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_239
timestamp 1604681595
transform 1 0 23092 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_251
timestamp 1604681595
transform 1 0 24196 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 24564 0 1 10056
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 25116 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 24380 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_263
timestamp 1604681595
transform 1 0 25300 0 1 10056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1604681595
transform 1 0 4692 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1604681595
transform 1 0 6532 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_74
timestamp 1604681595
transform 1 0 7912 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10304 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_98
timestamp 1604681595
transform 1 0 10120 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1604681595
transform 1 0 10488 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_114
timestamp 1604681595
transform 1 0 11592 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13064 0 -1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1604681595
transform 1 0 12420 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_127
timestamp 1604681595
transform 1 0 12788 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1604681595
transform 1 0 13892 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_151
timestamp 1604681595
transform 1 0 14996 0 -1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16652 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_171
timestamp 1604681595
transform 1 0 16836 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1604681595
transform 1 0 18032 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19228 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_188
timestamp 1604681595
transform 1 0 18400 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_195
timestamp 1604681595
transform 1 0 19044 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_199
timestamp 1604681595
transform 1 0 19412 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_211
timestamp 1604681595
transform 1 0 20516 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_223
timestamp 1604681595
transform 1 0 21620 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_235
timestamp 1604681595
transform 1 0 22724 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_243
timestamp 1604681595
transform 1 0 23460 0 -1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_245
timestamp 1604681595
transform 1 0 23644 0 -1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 24564 0 -1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1604681595
transform 1 0 24380 0 -1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1604681595
transform 1 0 4048 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1604681595
transform 1 0 5152 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1604681595
transform 1 0 6256 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_68
timestamp 1604681595
transform 1 0 7360 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_80
timestamp 1604681595
transform 1 0 8464 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10304 0 1 11144
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10120 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1604681595
transform 1 0 9660 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12512 0 1 11144
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12328 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604681595
transform 1 0 12144 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14168 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_150
timestamp 1604681595
transform 1 0 14904 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15364 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16468 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15824 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16652 0 1 11144
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1604681595
transform 1 0 18124 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 11144
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18308 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_189
timestamp 1604681595
transform 1 0 18492 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_202
timestamp 1604681595
transform 1 0 19688 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1604681595
transform 1 0 20424 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1604681595
transform 1 0 21252 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_223
timestamp 1604681595
transform 1 0 21620 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_235
timestamp 1604681595
transform 1 0 22724 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_247
timestamp 1604681595
transform 1 0 23828 0 1 11144
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 24564 0 1 11144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_276
timestamp 1604681595
transform 1 0 26496 0 1 11144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1604681595
transform 1 0 4692 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1604681595
transform 1 0 5796 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1604681595
transform 1 0 6532 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_62
timestamp 1604681595
transform 1 0 6808 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_86
timestamp 1604681595
transform 1 0 9016 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_98
timestamp 1604681595
transform 1 0 10120 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 12232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15180 0 -1 12232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18124 0 -1 12232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_169
timestamp 1604681595
transform 1 0 16652 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1604681595
transform 1 0 17756 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1604681595
transform 1 0 19596 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20792 0 -1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604681595
transform 1 0 20700 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_223
timestamp 1604681595
transform 1 0 21620 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_235
timestamp 1604681595
transform 1 0 22724 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_243
timestamp 1604681595
transform 1 0 23460 0 -1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 24564 0 -1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1604681595
transform 1 0 24380 0 -1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_259
timestamp 1604681595
transform 1 0 24932 0 -1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_271
timestamp 1604681595
transform 1 0 26036 0 -1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1604681595
transform 1 0 6256 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_51
timestamp 1604681595
transform 1 0 5796 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1604681595
transform 1 0 6808 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_68
timestamp 1604681595
transform 1 0 7360 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1604681595
transform 1 0 8464 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1604681595
transform 1 0 9660 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_86
timestamp 1604681595
transform 1 0 9016 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_98
timestamp 1604681595
transform 1 0 10120 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 12696 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1604681595
transform 1 0 12788 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13156 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_133
timestamp 1604681595
transform 1 0 13340 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13156 0 1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_140
timestamp 1604681595
transform 1 0 13984 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_146
timestamp 1604681595
transform 1 0 14536 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1604681595
transform 1 0 15180 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1604681595
transform 1 0 15456 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16652 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16652 0 -1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1604681595
transform 1 0 18032 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1604681595
transform 1 0 17388 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17572 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 12232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 18216 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19596 0 -1 13320
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19596 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18676 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_200
timestamp 1604681595
transform 1 0 19504 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1604681595
transform 1 0 18492 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_193
timestamp 1604681595
transform 1 0 18860 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20884 0 1 12232
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1604681595
transform 1 0 19780 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1604681595
transform 1 0 20148 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_211
timestamp 1604681595
transform 1 0 20516 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_217
timestamp 1604681595
transform 1 0 21068 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 21804 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21252 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_231
timestamp 1604681595
transform 1 0 22356 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1604681595
transform 1 0 21436 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_228
timestamp 1604681595
transform 1 0 22080 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 24012 0 1 12232
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 -1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_243
timestamp 1604681595
transform 1 0 23460 0 1 12232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_240
timestamp 1604681595
transform 1 0 23184 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_245
timestamp 1604681595
transform 1 0 23644 0 -1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 24564 0 -1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 24564 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 24932 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_253
timestamp 1604681595
transform 1 0 24380 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1604681595
transform 1 0 24380 0 -1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1604681595
transform 1 0 24932 0 -1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_273
timestamp 1604681595
transform 1 0 26220 0 1 12232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_271
timestamp 1604681595
transform 1 0 26036 0 -1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1604681595
transform 1 0 5152 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_56
timestamp 1604681595
transform 1 0 6256 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_68
timestamp 1604681595
transform 1 0 7360 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_80
timestamp 1604681595
transform 1 0 8464 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_105
timestamp 1604681595
transform 1 0 10764 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_117
timestamp 1604681595
transform 1 0 11868 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12696 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 13432 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12512 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_148
timestamp 1604681595
transform 1 0 14720 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16008 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16376 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_164
timestamp 1604681595
transform 1 0 16192 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_168
timestamp 1604681595
transform 1 0 16560 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 16652 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17940 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17572 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 17204 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1604681595
transform 1 0 17020 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1604681595
transform 1 0 17388 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1604681595
transform 1 0 17756 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1604681595
transform 1 0 18124 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18492 0 1 13320
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 18308 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19504 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1604681595
transform 1 0 19320 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1604681595
transform 1 0 19688 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 13320
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1604681595
transform 1 0 20056 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1604681595
transform 1 0 20424 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_224
timestamp 1604681595
transform 1 0 21712 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_228
timestamp 1604681595
transform 1 0 22080 0 1 13320
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_246
timestamp 1604681595
transform 1 0 23736 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 24564 0 1 13320
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 25116 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 25484 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_259
timestamp 1604681595
transform 1 0 24932 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_263
timestamp 1604681595
transform 1 0 25300 0 1 13320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_267
timestamp 1604681595
transform 1 0 25668 0 1 13320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1604681595
transform 1 0 4692 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1604681595
transform 1 0 5796 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1604681595
transform 1 0 6532 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1604681595
transform 1 0 6808 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1604681595
transform 1 0 7912 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1604681595
transform 1 0 10120 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_110
timestamp 1604681595
transform 1 0 11224 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 13432 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_131
timestamp 1604681595
transform 1 0 13156 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_138
timestamp 1604681595
transform 1 0 13800 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1604681595
transform 1 0 14904 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 -1 14408
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 15272 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_156
timestamp 1604681595
transform 1 0 15456 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1604681595
transform 1 0 17020 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1604681595
transform 1 0 17756 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_184
timestamp 1604681595
transform 1 0 18032 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 14408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20792 0 -1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_203
timestamp 1604681595
transform 1 0 19780 0 -1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1604681595
transform 1 0 20516 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22448 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_220
timestamp 1604681595
transform 1 0 21344 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1604681595
transform 1 0 22632 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 -1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 -1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22816 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1604681595
transform 1 0 23644 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 25116 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24564 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1604681595
transform 1 0 24380 0 -1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_257
timestamp 1604681595
transform 1 0 24748 0 -1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1604681595
transform 1 0 25484 0 -1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1604681595
transform 1 0 4048 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1604681595
transform 1 0 5152 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_56
timestamp 1604681595
transform 1 0 6256 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_68
timestamp 1604681595
transform 1 0 7360 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_80
timestamp 1604681595
transform 1 0 8464 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1604681595
transform 1 0 9660 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_117
timestamp 1604681595
transform 1 0 11868 0 1 14408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_129
timestamp 1604681595
transform 1 0 12972 0 1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13616 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13984 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1604681595
transform 1 0 13800 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_142
timestamp 1604681595
transform 1 0 14168 0 1 14408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_150
timestamp 1604681595
transform 1 0 14904 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 15272 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16468 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_158
timestamp 1604681595
transform 1 0 15640 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16652 0 1 14408
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1604681595
transform 1 0 18124 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 14408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18676 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_189
timestamp 1604681595
transform 1 0 18492 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1604681595
transform 1 0 19688 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 20884 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19872 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_206
timestamp 1604681595
transform 1 0 20056 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1604681595
transform 1 0 20424 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1604681595
transform 1 0 21160 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 22448 0 1 14408
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 21344 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21712 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_226
timestamp 1604681595
transform 1 0 21896 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 1 14408
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23644 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_241
timestamp 1604681595
transform 1 0 23276 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_247
timestamp 1604681595
transform 1 0 23828 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 25300 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 25852 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 25116 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1604681595
transform 1 0 24564 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1604681595
transform 1 0 24932 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1604681595
transform 1 0 25668 0 1 14408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_271
timestamp 1604681595
transform 1 0 26036 0 1 14408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1604681595
transform 1 0 5796 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604681595
transform 1 0 6532 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1604681595
transform 1 0 6808 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1604681595
transform 1 0 7912 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13616 0 -1 15496
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_135
timestamp 1604681595
transform 1 0 13524 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 -1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15732 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_156
timestamp 1604681595
transform 1 0 15456 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16928 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1604681595
transform 1 0 16744 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_174
timestamp 1604681595
transform 1 0 17112 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18952 0 -1 15496
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21160 0 -1 15496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_234
timestamp 1604681595
transform 1 0 22632 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 -1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 22816 0 -1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_238
timestamp 1604681595
transform 1 0 23000 0 -1 15496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 25208 0 -1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_254
timestamp 1604681595
transform 1 0 24472 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_266
timestamp 1604681595
transform 1 0 25576 0 -1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1604681595
transform 1 0 4048 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1604681595
transform 1 0 5152 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_56
timestamp 1604681595
transform 1 0 6256 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_68
timestamp 1604681595
transform 1 0 7360 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_80
timestamp 1604681595
transform 1 0 8464 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_105
timestamp 1604681595
transform 1 0 10764 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_117
timestamp 1604681595
transform 1 0 11868 0 1 15496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14260 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1604681595
transform 1 0 13708 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_141
timestamp 1604681595
transform 1 0 14076 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1604681595
transform 1 0 14444 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1604681595
transform 1 0 16100 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_167
timestamp 1604681595
transform 1 0 16468 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16836 0 1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16652 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18584 0 1 15496
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18400 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_186
timestamp 1604681595
transform 1 0 18216 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_199
timestamp 1604681595
transform 1 0 19412 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1604681595
transform 1 0 20148 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1604681595
transform 1 0 20516 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 22172 0 1 15496
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 21988 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_219
timestamp 1604681595
transform 1 0 21252 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_223
timestamp 1604681595
transform 1 0 21620 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23920 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1604681595
transform 1 0 24104 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 24564 0 1 15496
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 25116 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 25484 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1604681595
transform 1 0 24932 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_263
timestamp 1604681595
transform 1 0 25300 0 1 15496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_267
timestamp 1604681595
transform 1 0 25668 0 1 15496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1604681595
transform 1 0 4048 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1604681595
transform 1 0 4692 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1604681595
transform 1 0 5796 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1604681595
transform 1 0 6532 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_74
timestamp 1604681595
transform 1 0 7912 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_68
timestamp 1604681595
transform 1 0 7360 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_80
timestamp 1604681595
transform 1 0 8464 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_98
timestamp 1604681595
transform 1 0 10120 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1604681595
transform 1 0 9660 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_110
timestamp 1604681595
transform 1 0 11224 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1604681595
transform 1 0 12972 0 1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_140
timestamp 1604681595
transform 1 0 13984 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_148
timestamp 1604681595
transform 1 0 14720 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1604681595
transform 1 0 14352 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14996 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14260 0 -1 16584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 16468 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 1 16584
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15916 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16284 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_159
timestamp 1604681595
transform 1 0 15732 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_176
timestamp 1604681595
transform 1 0 17296 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1604681595
transform 1 0 16744 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16928 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_182
timestamp 1604681595
transform 1 0 17848 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 17572 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_174
timestamp 1604681595
transform 1 0 17112 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18584 0 1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18676 0 -1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19596 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_188
timestamp 1604681595
transform 1 0 18400 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1604681595
transform 1 0 19504 0 -1 16584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_186
timestamp 1604681595
transform 1 0 18216 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1604681595
transform 1 0 19412 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20700 0 -1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_212
timestamp 1604681595
transform 1 0 20608 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_207
timestamp 1604681595
transform 1 0 20148 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1604681595
transform 1 0 20700 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1604681595
transform 1 0 20884 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1604681595
transform 1 0 21528 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1604681595
transform 1 0 21252 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_222
timestamp 1604681595
transform 1 0 21528 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21804 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21344 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21712 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_235
timestamp 1604681595
transform 1 0 22724 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1604681595
transform 1 0 22356 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22172 0 -1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 22540 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21896 0 1 16584
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_243
timestamp 1604681595
transform 1 0 23460 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_239
timestamp 1604681595
transform 1 0 23092 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22908 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 -1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1604681595
transform 1 0 23828 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_245
timestamp 1604681595
transform 1 0 23644 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23920 0 1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23920 0 -1 16584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_236
timestamp 1604681595
transform 1 0 22816 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 25024 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24656 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_266
timestamp 1604681595
transform 1 0 25576 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 25760 0 1 16584
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 25208 0 -1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 25208 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1604681595
transform 1 0 25576 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_254
timestamp 1604681595
transform 1 0 24472 0 -1 16584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1604681595
transform 1 0 25944 0 1 16584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_274
timestamp 1604681595
transform 1 0 26312 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_39
timestamp 1604681595
transform 1 0 4692 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1604681595
transform 1 0 6808 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1604681595
transform 1 0 9016 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1604681595
transform 1 0 10120 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1604681595
transform 1 0 12420 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14168 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_28_135
timestamp 1604681595
transform 1 0 13524 0 -1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_151
timestamp 1604681595
transform 1 0 14996 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 17672
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_156
timestamp 1604681595
transform 1 0 15456 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_175
timestamp 1604681595
transform 1 0 17204 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19596 0 -1 17672
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19412 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1604681595
transform 1 0 18860 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1604681595
transform 1 0 19228 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_217
timestamp 1604681595
transform 1 0 21068 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21804 0 -1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_222
timestamp 1604681595
transform 1 0 21528 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 -1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_242
timestamp 1604681595
transform 1 0 23368 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_245
timestamp 1604681595
transform 1 0 23644 0 -1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 24564 0 -1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1604681595
transform 1 0 24380 0 -1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1604681595
transform 1 0 4048 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1604681595
transform 1 0 5152 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_56
timestamp 1604681595
transform 1 0 6256 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1604681595
transform 1 0 7360 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_80
timestamp 1604681595
transform 1 0 8464 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1604681595
transform 1 0 9660 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_105
timestamp 1604681595
transform 1 0 10764 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_117
timestamp 1604681595
transform 1 0 11868 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_129
timestamp 1604681595
transform 1 0 12972 0 1 17672
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1604681595
transform 1 0 14812 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15364 0 1 17672
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_154
timestamp 1604681595
transform 1 0 15272 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17848 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16744 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17112 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17480 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1604681595
transform 1 0 17296 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18400 0 1 17672
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 18216 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20884 0 1 17672
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 20056 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_204
timestamp 1604681595
transform 1 0 19872 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 22540 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1604681595
transform 1 0 22356 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_235
timestamp 1604681595
transform 1 0 22724 0 1 17672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23644 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_243
timestamp 1604681595
transform 1 0 23460 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 25116 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 25668 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24564 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_253
timestamp 1604681595
transform 1 0 24380 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_265
timestamp 1604681595
transform 1 0 25484 0 1 17672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_39
timestamp 1604681595
transform 1 0 4692 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1604681595
transform 1 0 5796 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_74
timestamp 1604681595
transform 1 0 7912 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_86
timestamp 1604681595
transform 1 0 9016 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_98
timestamp 1604681595
transform 1 0 10120 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_110
timestamp 1604681595
transform 1 0 11224 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1604681595
transform 1 0 12236 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13984 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_135
timestamp 1604681595
transform 1 0 13524 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1604681595
transform 1 0 13800 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_142
timestamp 1604681595
transform 1 0 14168 0 -1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15640 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_156
timestamp 1604681595
transform 1 0 15456 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1604681595
transform 1 0 15824 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_164
timestamp 1604681595
transform 1 0 16192 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 -1 18760
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1604681595
transform 1 0 17204 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_200
timestamp 1604681595
transform 1 0 19504 0 -1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 20332 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20148 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_217
timestamp 1604681595
transform 1 0 21068 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21344 0 -1 18760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 -1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_236
timestamp 1604681595
transform 1 0 22816 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1604681595
transform 1 0 23184 0 -1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_245
timestamp 1604681595
transform 1 0 23644 0 -1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 25300 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_255
timestamp 1604681595
transform 1 0 24564 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_32
timestamp 1604681595
transform 1 0 4048 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_44
timestamp 1604681595
transform 1 0 5152 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_56
timestamp 1604681595
transform 1 0 6256 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_68
timestamp 1604681595
transform 1 0 7360 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_80
timestamp 1604681595
transform 1 0 8464 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_105
timestamp 1604681595
transform 1 0 10764 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_128
timestamp 1604681595
transform 1 0 12880 0 1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1604681595
transform 1 0 14444 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 18760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_183
timestamp 1604681595
transform 1 0 17940 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 18216 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18676 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1604681595
transform 1 0 18492 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 18760
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 18760
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1604681595
transform 1 0 19964 0 1 18760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1604681595
transform 1 0 20516 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22724 0 1 18760
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22540 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_224
timestamp 1604681595
transform 1 0 21712 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_229
timestamp 1604681595
transform 1 0 22172 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_251
timestamp 1604681595
transform 1 0 24196 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 24932 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24748 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 25484 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 25852 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_255
timestamp 1604681595
transform 1 0 24564 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_267
timestamp 1604681595
transform 1 0 25668 0 1 18760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 18760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_271
timestamp 1604681595
transform 1 0 26036 0 1 18760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604681595
transform 1 0 26496 0 1 18760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1604681595
transform 1 0 4692 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_62
timestamp 1604681595
transform 1 0 6808 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_74
timestamp 1604681595
transform 1 0 7912 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_98
timestamp 1604681595
transform 1 0 10120 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10488 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_104
timestamp 1604681595
transform 1 0 10672 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_116
timestamp 1604681595
transform 1 0 11776 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 12420 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13248 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12052 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1604681595
transform 1 0 13064 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1604681595
transform 1 0 13432 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13892 0 -1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_138
timestamp 1604681595
transform 1 0 13800 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 16100 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15640 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_155
timestamp 1604681595
transform 1 0 15364 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_160
timestamp 1604681595
transform 1 0 15824 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 17940 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18676 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_188
timestamp 1604681595
transform 1 0 18400 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1604681595
transform 1 0 19228 0 -1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20884 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_209
timestamp 1604681595
transform 1 0 20332 0 -1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_217
timestamp 1604681595
transform 1 0 21068 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 -1 19848
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 -1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 19848
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 23552 0 -1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_236
timestamp 1604681595
transform 1 0 22816 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 25208 0 -1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_254
timestamp 1604681595
transform 1 0 24472 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_266
timestamp 1604681595
transform 1 0 25576 0 -1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_274
timestamp 1604681595
transform 1 0 26312 0 -1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 3956 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_39
timestamp 1604681595
transform 1 0 4692 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 6716 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1604681595
transform 1 0 5796 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1604681595
transform 1 0 6532 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_62
timestamp 1604681595
transform 1 0 6808 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_68
timestamp 1604681595
transform 1 0 7360 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_80
timestamp 1604681595
transform 1 0 8464 0 1 19848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_74
timestamp 1604681595
transform 1 0 7912 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 9568 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 10304 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_93
timestamp 1604681595
transform 1 0 9660 0 1 19848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_86
timestamp 1604681595
transform 1 0 9016 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_98
timestamp 1604681595
transform 1 0 10120 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10488 0 1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1604681595
transform 1 0 11224 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_114
timestamp 1604681595
transform 1 0 11592 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 -1 20936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12696 0 1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 12328 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12512 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1604681595
transform 1 0 12328 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_121
timestamp 1604681595
transform 1 0 12236 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1604681595
transform 1 0 14168 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14260 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1604681595
transform 1 0 14812 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_146
timestamp 1604681595
transform 1 0 14536 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 14628 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_150
timestamp 1604681595
transform 1 0 14904 0 -1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15640 0 -1 20936
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 15180 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_156
timestamp 1604681595
transform 1 0 15456 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1604681595
transform 1 0 17296 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_170
timestamp 1604681595
transform 1 0 16744 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17112 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_182
timestamp 1604681595
transform 1 0 17848 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17480 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17848 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 17940 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_174
timestamp 1604681595
transform 1 0 17112 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 -1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19688 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1604681595
transform 1 0 19504 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_193
timestamp 1604681595
transform 1 0 18860 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_205
timestamp 1604681595
transform 1 0 19964 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_213
timestamp 1604681595
transform 1 0 20700 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20516 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 20792 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 20884 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20148 0 -1 20936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22724 0 1 19848
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 22540 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 22724 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21988 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_226
timestamp 1604681595
transform 1 0 21896 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1604681595
transform 1 0 22172 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_223
timestamp 1604681595
transform 1 0 21620 0 -1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 -1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 23552 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_251
timestamp 1604681595
transform 1 0 24196 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_237
timestamp 1604681595
transform 1 0 22908 0 -1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_243
timestamp 1604681595
transform 1 0 23460 0 -1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1604681595
transform 1 0 23644 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_255
timestamp 1604681595
transform 1 0 24564 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 24748 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 24932 0 1 19848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1604681595
transform 1 0 25300 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25484 0 1 19848
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25116 0 -1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_267
timestamp 1604681595
transform 1 0 25668 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1604681595
transform 1 0 24380 0 -1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_267
timestamp 1604681595
transform 1 0 25668 0 1 19848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 19848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26404 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 19848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_275
timestamp 1604681595
transform 1 0 26404 0 -1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 3956 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_68
timestamp 1604681595
transform 1 0 7360 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 9568 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1604681595
transform 1 0 9660 0 1 20936
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11684 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_105
timestamp 1604681595
transform 1 0 10764 0 1 20936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13248 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13064 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_124
timestamp 1604681595
transform 1 0 12512 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp 1604681595
transform 1 0 14168 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1604681595
transform 1 0 14444 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 15180 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_154
timestamp 1604681595
transform 1 0 15272 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_158
timestamp 1604681595
transform 1 0 15640 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17572 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1604681595
transform 1 0 17756 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1604681595
transform 1 0 18952 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_198
timestamp 1604681595
transform 1 0 19320 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 20936
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 20792 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 19872 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_206
timestamp 1604681595
transform 1 0 20056 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1604681595
transform 1 0 20424 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 22724 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_224
timestamp 1604681595
transform 1 0 21712 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_228
timestamp 1604681595
transform 1 0 22080 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23828 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 23276 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23644 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_239
timestamp 1604681595
transform 1 0 23092 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_243
timestamp 1604681595
transform 1 0 23460 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 25116 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 24564 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 25668 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_253
timestamp 1604681595
transform 1 0 24380 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 20936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_265
timestamp 1604681595
transform 1 0 25484 0 1 20936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 20936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 20936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 26404 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 20936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_39
timestamp 1604681595
transform 1 0 4692 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 6716 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_51
timestamp 1604681595
transform 1 0 5796 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_59
timestamp 1604681595
transform 1 0 6532 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_62
timestamp 1604681595
transform 1 0 6808 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_74
timestamp 1604681595
transform 1 0 7912 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_86
timestamp 1604681595
transform 1 0 9016 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_98
timestamp 1604681595
transform 1 0 10120 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11684 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_104
timestamp 1604681595
transform 1 0 10672 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1604681595
transform 1 0 10948 0 -1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_113
timestamp 1604681595
transform 1 0 11500 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 12328 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1604681595
transform 1 0 12236 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1604681595
transform 1 0 12420 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14260 0 -1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1604681595
transform 1 0 13524 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16192 0 -1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15640 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_152
timestamp 1604681595
transform 1 0 15088 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_160
timestamp 1604681595
transform 1 0 15824 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 17940 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17204 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_173
timestamp 1604681595
transform 1 0 17020 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_177
timestamp 1604681595
transform 1 0 17388 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 20240 0 -1 22024
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 22540 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_224
timestamp 1604681595
transform 1 0 21712 0 -1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_232
timestamp 1604681595
transform 1 0 22448 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 23552 0 -1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_236
timestamp 1604681595
transform 1 0 22816 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1604681595
transform 1 0 23184 0 -1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_245
timestamp 1604681595
transform 1 0 23644 0 -1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_249
timestamp 1604681595
transform 1 0 24012 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 24564 0 -1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_259
timestamp 1604681595
transform 1 0 24932 0 -1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_271
timestamp 1604681595
transform 1 0 26036 0 -1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_32
timestamp 1604681595
transform 1 0 4048 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_44
timestamp 1604681595
transform 1 0 5152 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_56
timestamp 1604681595
transform 1 0 6256 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_68
timestamp 1604681595
transform 1 0 7360 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_80
timestamp 1604681595
transform 1 0 8464 0 1 22024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_93
timestamp 1604681595
transform 1 0 9660 0 1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11316 0 1 22024
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_103
timestamp 1604681595
transform 1 0 10580 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_107
timestamp 1604681595
transform 1 0 10948 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12972 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_131
timestamp 1604681595
transform 1 0 13156 0 1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13892 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 14260 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_141
timestamp 1604681595
transform 1 0 14076 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_145
timestamp 1604681595
transform 1 0 14444 0 1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15916 0 1 22024
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 15180 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15732 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_154
timestamp 1604681595
transform 1 0 15272 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_158
timestamp 1604681595
transform 1 0 15640 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18032 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17572 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1604681595
transform 1 0 17388 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_181
timestamp 1604681595
transform 1 0 17756 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 19504 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18400 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_186
timestamp 1604681595
transform 1 0 18216 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_190
timestamp 1604681595
transform 1 0 18584 0 1 22024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_198
timestamp 1604681595
transform 1 0 19320 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 22024
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 20792 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1604681595
transform 1 0 19780 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_207
timestamp 1604681595
transform 1 0 20148 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 22540 0 1 22024
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22356 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_224
timestamp 1604681595
transform 1 0 21712 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_228
timestamp 1604681595
transform 1 0 22080 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_249
timestamp 1604681595
transform 1 0 24012 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 24748 0 1 22024
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 25300 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24564 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 25668 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1604681595
transform 1 0 24380 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1604681595
transform 1 0 25116 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_265
timestamp 1604681595
transform 1 0 25484 0 1 22024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 26404 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_39
timestamp 1604681595
transform 1 0 4692 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6716 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_51
timestamp 1604681595
transform 1 0 5796 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_59
timestamp 1604681595
transform 1 0 6532 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_62
timestamp 1604681595
transform 1 0 6808 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_74
timestamp 1604681595
transform 1 0 7912 0 -1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 9752 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_86
timestamp 1604681595
transform 1 0 9016 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_38_114
timestamp 1604681595
transform 1 0 11592 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 12328 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13892 0 -1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13616 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_135
timestamp 1604681595
transform 1 0 13524 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_138
timestamp 1604681595
transform 1 0 13800 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 15916 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_155
timestamp 1604681595
transform 1 0 15364 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_159
timestamp 1604681595
transform 1 0 15732 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_163
timestamp 1604681595
transform 1 0 16100 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 -1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 17940 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_175
timestamp 1604681595
transform 1 0 17204 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_200
timestamp 1604681595
transform 1 0 19504 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 21068 0 -1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20516 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_204
timestamp 1604681595
transform 1 0 19872 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_213
timestamp 1604681595
transform 1 0 20700 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22724 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_233
timestamp 1604681595
transform 1 0 22540 0 -1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 23552 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_237
timestamp 1604681595
transform 1 0 22908 0 -1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_243
timestamp 1604681595
transform 1 0 23460 0 -1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 25208 0 -1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_254
timestamp 1604681595
transform 1 0 24472 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1604681595
transform 1 0 25576 0 -1 23112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_274
timestamp 1604681595
transform 1 0 26312 0 -1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 3956 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_32
timestamp 1604681595
transform 1 0 4048 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_44
timestamp 1604681595
transform 1 0 5152 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_39
timestamp 1604681595
transform 1 0 4692 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 6716 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_56
timestamp 1604681595
transform 1 0 6256 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_51
timestamp 1604681595
transform 1 0 5796 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_59
timestamp 1604681595
transform 1 0 6532 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_62
timestamp 1604681595
transform 1 0 6808 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_68
timestamp 1604681595
transform 1 0 7360 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_80
timestamp 1604681595
transform 1 0 8464 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_74
timestamp 1604681595
transform 1 0 7912 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 9568 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1604681595
transform 1 0 9660 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_86
timestamp 1604681595
transform 1 0 9016 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_98
timestamp 1604681595
transform 1 0 10120 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11408 0 1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10856 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_105
timestamp 1604681595
transform 1 0 10764 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_108
timestamp 1604681595
transform 1 0 11040 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_114
timestamp 1604681595
transform 1 0 11592 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 12328 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13064 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_128
timestamp 1604681595
transform 1 0 12880 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1604681595
transform 1 0 12420 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13892 0 -1 24200
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_145
timestamp 1604681595
transform 1 0 14444 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1604681595
transform 1 0 14812 0 1 23112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_135
timestamp 1604681595
transform 1 0 13524 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_138
timestamp 1604681595
transform 1 0 13800 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_157
timestamp 1604681595
transform 1 0 15548 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 15180 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 15272 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_162
timestamp 1604681595
transform 1 0 16008 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16100 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 15824 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_155
timestamp 1604681595
transform 1 0 15364 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 24200
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16376 0 1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 17940 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_182
timestamp 1604681595
transform 1 0 17848 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_174
timestamp 1604681595
transform 1 0 17112 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_182
timestamp 1604681595
transform 1 0 17848 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_184
timestamp 1604681595
transform 1 0 18032 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 1 23112
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 24200
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18584 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_186
timestamp 1604681595
transform 1 0 18216 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_188
timestamp 1604681595
transform 1 0 18400 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_192
timestamp 1604681595
transform 1 0 18768 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_210
timestamp 1604681595
transform 1 0 20424 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1604681595
transform 1 0 20424 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_206
timestamp 1604681595
transform 1 0 20056 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_217
timestamp 1604681595
transform 1 0 21068 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_213
timestamp 1604681595
transform 1 0 20700 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20884 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 20792 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1604681595
transform 1 0 21712 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 21896 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 21344 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1604681595
transform 1 0 22080 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_229
timestamp 1604681595
transform 1 0 22172 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 22448 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22540 0 1 23112
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1604681595
transform 1 0 23184 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_236
timestamp 1604681595
transform 1 0 22816 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_242
timestamp 1604681595
transform 1 0 23368 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 23000 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_247
timestamp 1604681595
transform 1 0 23828 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23644 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 23552 0 -1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24104 0 1 23112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 24932 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 24932 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_256
timestamp 1604681595
transform 1 0 24656 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1604681595
transform 1 0 25116 0 1 23112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 26404 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_273
timestamp 1604681595
transform 1 0 26220 0 1 23112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_275
timestamp 1604681595
transform 1 0 26404 0 -1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 3956 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_32
timestamp 1604681595
transform 1 0 4048 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_44
timestamp 1604681595
transform 1 0 5152 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_56
timestamp 1604681595
transform 1 0 6256 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_68
timestamp 1604681595
transform 1 0 7360 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_80
timestamp 1604681595
transform 1 0 8464 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 9568 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1604681595
transform 1 0 9660 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11408 0 1 24200
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11224 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_105
timestamp 1604681595
transform 1 0 10764 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_109
timestamp 1604681595
transform 1 0 11132 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_121
timestamp 1604681595
transform 1 0 12236 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_133
timestamp 1604681595
transform 1 0 13340 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_145
timestamp 1604681595
transform 1 0 14444 0 1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 15180 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16376 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_154
timestamp 1604681595
transform 1 0 15272 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 17388 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_176
timestamp 1604681595
transform 1 0 17296 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_180
timestamp 1604681595
transform 1 0 17664 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 20792 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_204
timestamp 1604681595
transform 1 0 19872 0 1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_212
timestamp 1604681595
transform 1 0 20608 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_215
timestamp 1604681595
transform 1 0 20884 0 1 24200
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 22540 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_227
timestamp 1604681595
transform 1 0 21988 0 1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 24200
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 23092 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 23460 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1604681595
transform 1 0 22908 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_241
timestamp 1604681595
transform 1 0 23276 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_251
timestamp 1604681595
transform 1 0 24196 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 24932 0 1 24200
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 25484 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 24748 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_255
timestamp 1604681595
transform 1 0 24564 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_267
timestamp 1604681595
transform 1 0 25668 0 1 24200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 26404 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604681595
transform 1 0 26496 0 1 24200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 3956 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 6808 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 9660 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 -1 25288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1604681595
transform 1 0 11592 0 -1 25288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 12512 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 15364 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 18216 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 21068 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 22816 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1604681595
transform 1 0 23920 0 -1 25288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 24564 0 -1 25288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25288
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 6664 480 6784 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 20672 480 20792 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 27520 3536 28000 3656 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 27520 9520 28000 9640 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 27520 10064 28000 10184 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 27520 10608 28000 10728 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 27520 11288 28000 11408 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 27520 11832 28000 11952 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 27520 12512 28000 12632 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 27520 13056 28000 13176 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 27520 13600 28000 13720 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 27520 14280 28000 14400 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 27520 14824 28000 14944 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 27520 4080 28000 4200 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 27520 4760 28000 4880 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 27520 5304 28000 5424 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 27520 5848 28000 5968 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 27520 6528 28000 6648 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 27520 7072 28000 7192 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 27520 7616 28000 7736 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 27520 8296 28000 8416 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 27520 8840 28000 8960 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 27520 15368 28000 15488 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 27520 21352 28000 21472 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 27520 22032 28000 22152 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 27520 22576 28000 22696 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 27520 23120 28000 23240 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 27520 23800 28000 23920 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 27520 24344 28000 24464 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 27520 25024 28000 25144 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 27520 25568 28000 25688 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 27520 26112 28000 26232 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 27520 26792 28000 26912 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 27520 16048 28000 16168 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 27520 16592 28000 16712 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 27520 17272 28000 17392 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 27520 17816 28000 17936 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 27520 18360 28000 18480 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 27520 19040 28000 19160 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 27520 19584 28000 19704 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 27520 20264 28000 20384 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 27520 20808 28000 20928 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 938 27240 994 27720 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 7746 27240 7802 27720 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8390 27240 8446 27720 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9126 27240 9182 27720 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9770 27240 9826 27720 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10506 27240 10562 27720 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 11150 27240 11206 27720 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11886 27240 11942 27720 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 12530 27240 12586 27720 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 13174 27240 13230 27720 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 13910 27240 13966 27720 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1582 27240 1638 27720 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 2318 27240 2374 27720 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2962 27240 3018 27720 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3698 27240 3754 27720 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 4342 27240 4398 27720 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4986 27240 5042 27720 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 5722 27240 5778 27720 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 6366 27240 6422 27720 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 7102 27240 7158 27720 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 14554 27240 14610 27720 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21362 27240 21418 27720 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22098 27240 22154 27720 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 22742 27240 22798 27720 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23478 27240 23534 27720 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24122 27240 24178 27720 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27240 24822 27720 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25502 27240 25558 27720 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 26146 27240 26202 27720 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26882 27240 26938 27720 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27526 27240 27582 27720 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 15290 27240 15346 27720 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 15934 27240 15990 27720 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 16578 27240 16634 27720 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 17314 27240 17370 27720 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 17958 27240 18014 27720 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 18694 27240 18750 27720 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 19338 27240 19394 27720 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20074 27240 20130 27720 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 20718 27240 20774 27720 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 27520 27336 28000 27456 6 prog_clk
port 82 nsew default input
rlabel metal3 s 27520 2856 28000 2976 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 27520 0 28000 120 6 right_bottom_grid_pin_1_
port 84 nsew default input
rlabel metal3 s 27520 544 28000 664 6 right_bottom_grid_pin_3_
port 85 nsew default input
rlabel metal3 s 27520 1088 28000 1208 6 right_bottom_grid_pin_5_
port 86 nsew default input
rlabel metal3 s 27520 1768 28000 1888 6 right_bottom_grid_pin_7_
port 87 nsew default input
rlabel metal3 s 27520 2312 28000 2432 6 right_bottom_grid_pin_9_
port 88 nsew default input
rlabel metal2 s 294 27240 350 27720 6 top_left_grid_pin_1_
port 89 nsew default input
rlabel metal4 s 5611 1848 5931 25336 6 VPWR
port 90 nsew default input
rlabel metal4 s 10277 1848 10597 25336 6 VGND
port 91 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27720
<< end >>
