magic
tech sky130A
magscale 1 2
timestamp 1608763155
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 6561 18139 6595 18309
rect 4445 16983 4479 17085
rect 2731 16949 2789 16983
rect 9413 16643 9447 16745
rect 13001 16439 13035 16745
rect 8033 14807 8067 14977
rect 11253 13175 11287 13277
rect 12173 13175 12207 13413
rect 4813 12767 4847 12937
rect 6653 12835 6687 12937
rect 7757 12631 7791 12869
rect 12173 12087 12207 12189
rect 6561 10659 6595 10761
rect 10057 8959 10091 9061
rect 10149 8823 10183 9061
rect 8217 8347 8251 8449
rect 11345 6647 11379 6749
rect 18797 5559 18831 5729
rect 10425 3927 10459 4097
rect 8493 3519 8527 3689
rect 10701 2907 10735 3077
rect 12265 2907 12299 3145
rect 2823 2465 2915 2499
rect 2881 2431 2915 2465
rect 15853 2363 15887 2465
<< viali >>
rect 2513 20009 2547 20043
rect 3065 20009 3099 20043
rect 3617 20009 3651 20043
rect 12817 20009 12851 20043
rect 18705 20009 18739 20043
rect 19533 20009 19567 20043
rect 10241 19941 10275 19975
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 2881 19873 2915 19907
rect 3433 19873 3467 19907
rect 5917 19873 5951 19907
rect 7757 19873 7791 19907
rect 10149 19873 10183 19907
rect 12633 19873 12667 19907
rect 13185 19873 13219 19907
rect 18521 19873 18555 19907
rect 19349 19873 19383 19907
rect 4077 19805 4111 19839
rect 6009 19805 6043 19839
rect 6193 19805 6227 19839
rect 7849 19805 7883 19839
rect 8033 19805 8067 19839
rect 10333 19805 10367 19839
rect 1961 19669 1995 19703
rect 5549 19669 5583 19703
rect 7389 19669 7423 19703
rect 9781 19669 9815 19703
rect 13369 19669 13403 19703
rect 3341 19465 3375 19499
rect 7849 19465 7883 19499
rect 10977 19397 11011 19431
rect 2697 19329 2731 19363
rect 4353 19329 4387 19363
rect 8493 19329 8527 19363
rect 9045 19329 9079 19363
rect 1685 19261 1719 19295
rect 1961 19261 1995 19295
rect 2421 19261 2455 19295
rect 3157 19261 3191 19295
rect 4077 19261 4111 19295
rect 4905 19261 4939 19295
rect 6837 19261 6871 19295
rect 8861 19261 8895 19295
rect 9597 19261 9631 19295
rect 11529 19261 11563 19295
rect 11805 19261 11839 19295
rect 12725 19261 12759 19295
rect 13001 19261 13035 19295
rect 13461 19261 13495 19295
rect 14013 19261 14047 19295
rect 14565 19261 14599 19295
rect 15117 19261 15151 19295
rect 15669 19261 15703 19295
rect 16221 19261 16255 19295
rect 16773 19261 16807 19295
rect 17325 19261 17359 19295
rect 18061 19261 18095 19295
rect 19257 19261 19291 19295
rect 20361 19261 20395 19295
rect 5172 19193 5206 19227
rect 7113 19193 7147 19227
rect 9864 19193 9898 19227
rect 19901 19193 19935 19227
rect 3709 19125 3743 19159
rect 4169 19125 4203 19159
rect 6285 19125 6319 19159
rect 8217 19125 8251 19159
rect 8309 19125 8343 19159
rect 13645 19125 13679 19159
rect 14197 19125 14231 19159
rect 14749 19125 14783 19159
rect 15301 19125 15335 19159
rect 15853 19125 15887 19159
rect 16405 19125 16439 19159
rect 16957 19125 16991 19159
rect 17509 19125 17543 19159
rect 18245 19125 18279 19159
rect 20545 19125 20579 19159
rect 3433 18921 3467 18955
rect 6469 18921 6503 18955
rect 6929 18921 6963 18955
rect 11069 18921 11103 18955
rect 13277 18921 13311 18955
rect 14749 18921 14783 18955
rect 16221 18921 16255 18955
rect 18245 18921 18279 18955
rect 19165 18921 19199 18955
rect 2329 18853 2363 18887
rect 7656 18853 7690 18887
rect 11888 18853 11922 18887
rect 1501 18785 1535 18819
rect 2053 18785 2087 18819
rect 3341 18785 3375 18819
rect 4077 18785 4111 18819
rect 5080 18785 5114 18819
rect 9956 18785 9990 18819
rect 11621 18785 11655 18819
rect 13645 18785 13679 18819
rect 13737 18785 13771 18819
rect 14565 18785 14599 18819
rect 15301 18785 15335 18819
rect 16037 18785 16071 18819
rect 18061 18785 18095 18819
rect 18981 18785 19015 18819
rect 3617 18717 3651 18751
rect 4813 18717 4847 18751
rect 7389 18717 7423 18751
rect 9137 18717 9171 18751
rect 9696 18717 9730 18751
rect 13829 18717 13863 18751
rect 15485 18717 15519 18751
rect 1685 18649 1719 18683
rect 4261 18649 4295 18683
rect 13001 18649 13035 18683
rect 2973 18581 3007 18615
rect 6193 18581 6227 18615
rect 8769 18581 8803 18615
rect 4905 18377 4939 18411
rect 5733 18377 5767 18411
rect 9689 18377 9723 18411
rect 14197 18377 14231 18411
rect 6561 18309 6595 18343
rect 12909 18309 12943 18343
rect 6193 18241 6227 18275
rect 6377 18241 6411 18275
rect 1869 18173 1903 18207
rect 3525 18173 3559 18207
rect 7389 18241 7423 18275
rect 10333 18241 10367 18275
rect 11437 18241 11471 18275
rect 15301 18241 15335 18275
rect 16865 18241 16899 18275
rect 18705 18241 18739 18275
rect 7656 18173 7690 18207
rect 10057 18173 10091 18207
rect 12725 18173 12759 18207
rect 13277 18173 13311 18207
rect 13553 18173 13587 18207
rect 14013 18173 14047 18207
rect 15025 18173 15059 18207
rect 16589 18173 16623 18207
rect 18429 18173 18463 18207
rect 2136 18105 2170 18139
rect 3792 18105 3826 18139
rect 6561 18105 6595 18139
rect 1409 18037 1443 18071
rect 3249 18037 3283 18071
rect 6101 18037 6135 18071
rect 8769 18037 8803 18071
rect 10149 18037 10183 18071
rect 10793 18037 10827 18071
rect 11161 18037 11195 18071
rect 11253 18037 11287 18071
rect 1685 17833 1719 17867
rect 2881 17833 2915 17867
rect 3341 17833 3375 17867
rect 4997 17833 5031 17867
rect 7941 17833 7975 17867
rect 8585 17833 8619 17867
rect 12541 17833 12575 17867
rect 12817 17833 12851 17867
rect 13829 17833 13863 17867
rect 2329 17765 2363 17799
rect 3249 17765 3283 17799
rect 6828 17765 6862 17799
rect 10057 17765 10091 17799
rect 13277 17765 13311 17799
rect 1501 17697 1535 17731
rect 2053 17697 2087 17731
rect 4077 17697 4111 17731
rect 5365 17697 5399 17731
rect 8677 17697 8711 17731
rect 9781 17697 9815 17731
rect 11428 17697 11462 17731
rect 13185 17697 13219 17731
rect 14197 17697 14231 17731
rect 3433 17629 3467 17663
rect 5457 17629 5491 17663
rect 5549 17629 5583 17663
rect 6561 17629 6595 17663
rect 8769 17629 8803 17663
rect 11161 17629 11195 17663
rect 13369 17629 13403 17663
rect 14289 17629 14323 17663
rect 14381 17629 14415 17663
rect 4261 17561 4295 17595
rect 8217 17493 8251 17527
rect 1869 17289 1903 17323
rect 11345 17289 11379 17323
rect 12449 17289 12483 17323
rect 5917 17221 5951 17255
rect 2329 17153 2363 17187
rect 2513 17153 2547 17187
rect 4537 17153 4571 17187
rect 8217 17153 8251 17187
rect 9597 17153 9631 17187
rect 13001 17153 13035 17187
rect 2881 17085 2915 17119
rect 4445 17085 4479 17119
rect 6193 17085 6227 17119
rect 9965 17085 9999 17119
rect 14105 17085 14139 17119
rect 14372 17085 14406 17119
rect 3148 17017 3182 17051
rect 4782 17017 4816 17051
rect 10232 17017 10266 17051
rect 12817 17017 12851 17051
rect 2237 16949 2271 16983
rect 2697 16949 2731 16983
rect 2789 16949 2823 16983
rect 4261 16949 4295 16983
rect 4445 16949 4479 16983
rect 7573 16949 7607 16983
rect 7941 16949 7975 16983
rect 8033 16949 8067 16983
rect 8953 16949 8987 16983
rect 9321 16949 9355 16983
rect 9413 16949 9447 16983
rect 11621 16949 11655 16983
rect 12909 16949 12943 16983
rect 15485 16949 15519 16983
rect 1685 16745 1719 16779
rect 5457 16745 5491 16779
rect 7297 16745 7331 16779
rect 7573 16745 7607 16779
rect 8033 16745 8067 16779
rect 8585 16745 8619 16779
rect 9413 16745 9447 16779
rect 11069 16745 11103 16779
rect 11345 16745 11379 16779
rect 11805 16745 11839 16779
rect 13001 16745 13035 16779
rect 14473 16745 14507 16779
rect 2329 16677 2363 16711
rect 4322 16677 4356 16711
rect 6184 16677 6218 16711
rect 8953 16677 8987 16711
rect 1501 16609 1535 16643
rect 2053 16609 2087 16643
rect 3341 16609 3375 16643
rect 7941 16609 7975 16643
rect 9413 16609 9447 16643
rect 9956 16609 9990 16643
rect 11713 16609 11747 16643
rect 3433 16541 3467 16575
rect 3617 16541 3651 16575
rect 4077 16541 4111 16575
rect 5917 16541 5951 16575
rect 8217 16541 8251 16575
rect 9045 16541 9079 16575
rect 9229 16541 9263 16575
rect 9689 16541 9723 16575
rect 11897 16541 11931 16575
rect 13360 16609 13394 16643
rect 13093 16541 13127 16575
rect 2973 16405 3007 16439
rect 13001 16405 13035 16439
rect 1685 16201 1719 16235
rect 3985 16201 4019 16235
rect 8585 16201 8619 16235
rect 10517 16201 10551 16235
rect 13829 16201 13863 16235
rect 15117 16201 15151 16235
rect 16129 16201 16163 16235
rect 5273 16133 5307 16167
rect 10241 16133 10275 16167
rect 2237 16065 2271 16099
rect 3065 16065 3099 16099
rect 3525 16065 3559 16099
rect 4537 16065 4571 16099
rect 5825 16065 5859 16099
rect 11069 16065 11103 16099
rect 14657 16065 14691 16099
rect 15669 16065 15703 16099
rect 16681 16065 16715 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2789 15997 2823 16031
rect 4445 15997 4479 16031
rect 7205 15997 7239 16031
rect 8861 15997 8895 16031
rect 9117 15997 9151 16031
rect 12449 15997 12483 16031
rect 12716 15997 12750 16031
rect 14565 15997 14599 16031
rect 15485 15997 15519 16031
rect 4353 15929 4387 15963
rect 5733 15929 5767 15963
rect 7472 15929 7506 15963
rect 10885 15929 10919 15963
rect 15577 15929 15611 15963
rect 16589 15929 16623 15963
rect 5641 15861 5675 15895
rect 10977 15861 11011 15895
rect 14105 15861 14139 15895
rect 14473 15861 14507 15895
rect 16497 15861 16531 15895
rect 1777 15657 1811 15691
rect 3065 15657 3099 15691
rect 8493 15657 8527 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 11253 15657 11287 15691
rect 11713 15657 11747 15691
rect 12265 15657 12299 15691
rect 14933 15657 14967 15691
rect 15301 15657 15335 15691
rect 2421 15589 2455 15623
rect 5448 15589 5482 15623
rect 1593 15521 1627 15555
rect 2134 15521 2168 15555
rect 2881 15521 2915 15555
rect 5181 15521 5215 15555
rect 7093 15521 7127 15555
rect 10057 15521 10091 15555
rect 11621 15521 11655 15555
rect 12633 15521 12667 15555
rect 13809 15521 13843 15555
rect 15669 15521 15703 15555
rect 6837 15453 6871 15487
rect 10241 15453 10275 15487
rect 11897 15453 11931 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 15761 15453 15795 15487
rect 15853 15453 15887 15487
rect 8217 15385 8251 15419
rect 6561 15317 6595 15351
rect 1777 15113 1811 15147
rect 12449 15113 12483 15147
rect 15209 15113 15243 15147
rect 2329 14977 2363 15011
rect 3065 14977 3099 15011
rect 5825 14977 5859 15011
rect 7481 14977 7515 15011
rect 8033 14977 8067 15011
rect 9689 14977 9723 15011
rect 10977 14977 11011 15011
rect 13093 14977 13127 15011
rect 13737 14977 13771 15011
rect 14749 14977 14783 15011
rect 15853 14977 15887 15011
rect 1593 14909 1627 14943
rect 2145 14909 2179 14943
rect 2881 14909 2915 14943
rect 4169 14909 4203 14943
rect 4436 14841 4470 14875
rect 7205 14841 7239 14875
rect 8309 14909 8343 14943
rect 12909 14909 12943 14943
rect 10793 14841 10827 14875
rect 12817 14841 12851 14875
rect 15669 14841 15703 14875
rect 5549 14773 5583 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 8033 14773 8067 14807
rect 8125 14773 8159 14807
rect 10425 14773 10459 14807
rect 10885 14773 10919 14807
rect 14197 14773 14231 14807
rect 14565 14773 14599 14807
rect 14657 14773 14691 14807
rect 15577 14773 15611 14807
rect 1869 14569 1903 14603
rect 2973 14569 3007 14603
rect 5457 14569 5491 14603
rect 10149 14569 10183 14603
rect 12357 14569 12391 14603
rect 12725 14569 12759 14603
rect 14013 14569 14047 14603
rect 6653 14501 6687 14535
rect 8208 14501 8242 14535
rect 11713 14501 11747 14535
rect 11805 14501 11839 14535
rect 15669 14501 15703 14535
rect 1685 14433 1719 14467
rect 2237 14433 2271 14467
rect 3341 14433 3375 14467
rect 4344 14433 4378 14467
rect 6009 14433 6043 14467
rect 6745 14433 6779 14467
rect 7941 14433 7975 14467
rect 10057 14433 10091 14467
rect 12817 14433 12851 14467
rect 14381 14433 14415 14467
rect 14473 14433 14507 14467
rect 15761 14433 15795 14467
rect 2421 14365 2455 14399
rect 3433 14365 3467 14399
rect 3617 14365 3651 14399
rect 4077 14365 4111 14399
rect 6837 14365 6871 14399
rect 10241 14365 10275 14399
rect 11989 14365 12023 14399
rect 13001 14365 13035 14399
rect 14657 14365 14691 14399
rect 15853 14365 15887 14399
rect 6285 14297 6319 14331
rect 9321 14297 9355 14331
rect 5825 14229 5859 14263
rect 9689 14229 9723 14263
rect 11345 14229 11379 14263
rect 15301 14229 15335 14263
rect 2789 14025 2823 14059
rect 4077 14025 4111 14059
rect 5365 14025 5399 14059
rect 8401 14025 8435 14059
rect 10057 14025 10091 14059
rect 12633 13957 12667 13991
rect 13185 13957 13219 13991
rect 14197 13957 14231 13991
rect 4721 13889 4755 13923
rect 6009 13889 6043 13923
rect 10885 13889 10919 13923
rect 11989 13889 12023 13923
rect 13737 13889 13771 13923
rect 15025 13889 15059 13923
rect 1869 13821 1903 13855
rect 2605 13821 2639 13855
rect 3145 13821 3179 13855
rect 4537 13821 4571 13855
rect 5825 13821 5859 13855
rect 7021 13821 7055 13855
rect 7277 13821 7311 13855
rect 8677 13821 8711 13855
rect 11805 13821 11839 13855
rect 12817 13821 12851 13855
rect 14381 13821 14415 13855
rect 15292 13821 15326 13855
rect 2145 13753 2179 13787
rect 5733 13753 5767 13787
rect 8944 13753 8978 13787
rect 10701 13753 10735 13787
rect 13553 13753 13587 13787
rect 3341 13685 3375 13719
rect 4445 13685 4479 13719
rect 10333 13685 10367 13719
rect 10793 13685 10827 13719
rect 11345 13685 11379 13719
rect 11713 13685 11747 13719
rect 13645 13685 13679 13719
rect 16405 13685 16439 13719
rect 4445 13481 4479 13515
rect 7389 13481 7423 13515
rect 7665 13481 7699 13515
rect 11713 13481 11747 13515
rect 12357 13481 12391 13515
rect 12817 13481 12851 13515
rect 15761 13481 15795 13515
rect 3433 13413 3467 13447
rect 11805 13413 11839 13447
rect 12173 13413 12207 13447
rect 15669 13413 15703 13447
rect 1869 13345 1903 13379
rect 3341 13345 3375 13379
rect 6276 13345 6310 13379
rect 8033 13345 8067 13379
rect 8677 13345 8711 13379
rect 9956 13345 9990 13379
rect 2053 13277 2087 13311
rect 3617 13277 3651 13311
rect 6009 13277 6043 13311
rect 8125 13277 8159 13311
rect 8217 13277 8251 13311
rect 9689 13277 9723 13311
rect 11253 13277 11287 13311
rect 11897 13277 11931 13311
rect 11345 13209 11379 13243
rect 2973 13141 3007 13175
rect 11069 13141 11103 13175
rect 11253 13141 11287 13175
rect 12725 13345 12759 13379
rect 13461 13345 13495 13379
rect 13728 13345 13762 13379
rect 12909 13277 12943 13311
rect 15945 13277 15979 13311
rect 14841 13209 14875 13243
rect 12173 13141 12207 13175
rect 15301 13141 15335 13175
rect 1593 12937 1627 12971
rect 1961 12937 1995 12971
rect 4813 12937 4847 12971
rect 2605 12801 2639 12835
rect 3617 12801 3651 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 6653 12937 6687 12971
rect 6929 12937 6963 12971
rect 12081 12937 12115 12971
rect 14197 12937 14231 12971
rect 14473 12937 14507 12971
rect 15485 12937 15519 12971
rect 7757 12869 7791 12903
rect 7941 12869 7975 12903
rect 5549 12801 5583 12835
rect 6653 12801 6687 12835
rect 7481 12801 7515 12835
rect 1409 12733 1443 12767
rect 2329 12733 2363 12767
rect 4353 12733 4387 12767
rect 4813 12733 4847 12767
rect 3341 12665 3375 12699
rect 5457 12665 5491 12699
rect 7297 12665 7331 12699
rect 9873 12801 9907 12835
rect 15025 12801 15059 12835
rect 16037 12801 16071 12835
rect 8125 12733 8159 12767
rect 10140 12733 10174 12767
rect 12265 12733 12299 12767
rect 12817 12733 12851 12767
rect 15853 12733 15887 12767
rect 13084 12665 13118 12699
rect 14933 12665 14967 12699
rect 15945 12665 15979 12699
rect 2421 12597 2455 12631
rect 2973 12597 3007 12631
rect 3433 12597 3467 12631
rect 3985 12597 4019 12631
rect 4997 12597 5031 12631
rect 5365 12597 5399 12631
rect 7389 12597 7423 12631
rect 7757 12597 7791 12631
rect 11253 12597 11287 12631
rect 14841 12597 14875 12631
rect 5457 12393 5491 12427
rect 7113 12393 7147 12427
rect 7481 12393 7515 12427
rect 8493 12393 8527 12427
rect 10057 12393 10091 12427
rect 10149 12393 10183 12427
rect 12725 12393 12759 12427
rect 12817 12393 12851 12427
rect 13369 12393 13403 12427
rect 1746 12325 1780 12359
rect 7941 12325 7975 12359
rect 10968 12325 11002 12359
rect 1501 12257 1535 12291
rect 4344 12257 4378 12291
rect 6000 12257 6034 12291
rect 7849 12257 7883 12291
rect 8861 12257 8895 12291
rect 10701 12257 10735 12291
rect 13737 12257 13771 12291
rect 15301 12257 15335 12291
rect 15568 12257 15602 12291
rect 4077 12189 4111 12223
rect 5733 12189 5767 12223
rect 8033 12189 8067 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 10241 12189 10275 12223
rect 12173 12189 12207 12223
rect 12909 12189 12943 12223
rect 13829 12189 13863 12223
rect 13921 12189 13955 12223
rect 2881 12053 2915 12087
rect 9689 12053 9723 12087
rect 12081 12053 12115 12087
rect 12173 12053 12207 12087
rect 12357 12053 12391 12087
rect 16681 12053 16715 12087
rect 2605 11849 2639 11883
rect 3617 11849 3651 11883
rect 6469 11849 6503 11883
rect 8309 11849 8343 11883
rect 13829 11849 13863 11883
rect 14105 11849 14139 11883
rect 10333 11781 10367 11815
rect 3249 11713 3283 11747
rect 4169 11713 4203 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10793 11713 10827 11747
rect 10977 11713 11011 11747
rect 11989 11713 12023 11747
rect 12449 11713 12483 11747
rect 14657 11713 14691 11747
rect 15117 11713 15151 11747
rect 17325 11713 17359 11747
rect 1685 11645 1719 11679
rect 3985 11645 4019 11679
rect 4077 11645 4111 11679
rect 5089 11645 5123 11679
rect 8033 11645 8067 11679
rect 9689 11645 9723 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 17141 11645 17175 11679
rect 17233 11645 17267 11679
rect 1961 11577 1995 11611
rect 2973 11577 3007 11611
rect 4629 11577 4663 11611
rect 5356 11577 5390 11611
rect 10701 11577 10735 11611
rect 12716 11577 12750 11611
rect 14565 11577 14599 11611
rect 15384 11577 15418 11611
rect 3065 11509 3099 11543
rect 6837 11509 6871 11543
rect 7849 11509 7883 11543
rect 8677 11509 8711 11543
rect 9321 11509 9355 11543
rect 11345 11509 11379 11543
rect 14473 11509 14507 11543
rect 16497 11509 16531 11543
rect 16773 11509 16807 11543
rect 1685 11305 1719 11339
rect 6469 11305 6503 11339
rect 9229 11305 9263 11339
rect 11437 11305 11471 11339
rect 11989 11305 12023 11339
rect 12449 11305 12483 11339
rect 12817 11305 12851 11339
rect 13277 11305 13311 11339
rect 13645 11305 13679 11339
rect 15301 11305 15335 11339
rect 16313 11305 16347 11339
rect 16773 11305 16807 11339
rect 2320 11237 2354 11271
rect 4344 11237 4378 11271
rect 9689 11237 9723 11271
rect 10149 11237 10183 11271
rect 13185 11237 13219 11271
rect 1501 11169 1535 11203
rect 4077 11169 4111 11203
rect 7113 11169 7147 11203
rect 7380 11169 7414 11203
rect 9137 11169 9171 11203
rect 12357 11169 12391 11203
rect 14013 11169 14047 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 16681 11169 16715 11203
rect 2053 11101 2087 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 9321 11101 9355 11135
rect 12633 11101 12667 11135
rect 13369 11101 13403 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 15945 11101 15979 11135
rect 16865 11101 16899 11135
rect 5457 11033 5491 11067
rect 3433 10965 3467 10999
rect 6101 10965 6135 10999
rect 8493 10965 8527 10999
rect 8769 10965 8803 10999
rect 1593 10761 1627 10795
rect 3801 10761 3835 10795
rect 4721 10761 4755 10795
rect 6561 10761 6595 10795
rect 8217 10761 8251 10795
rect 10149 10761 10183 10795
rect 13461 10761 13495 10795
rect 15853 10761 15887 10795
rect 9873 10693 9907 10727
rect 12449 10693 12483 10727
rect 2237 10625 2271 10659
rect 3249 10625 3283 10659
rect 5365 10625 5399 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 10793 10625 10827 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 14013 10625 14047 10659
rect 15485 10625 15519 10659
rect 16497 10625 16531 10659
rect 3617 10557 3651 10591
rect 6101 10557 6135 10591
rect 6837 10557 6871 10591
rect 8493 10557 8527 10591
rect 8749 10557 8783 10591
rect 13829 10557 13863 10591
rect 2053 10489 2087 10523
rect 2973 10489 3007 10523
rect 7104 10489 7138 10523
rect 10517 10489 10551 10523
rect 16221 10489 16255 10523
rect 1961 10421 1995 10455
rect 2605 10421 2639 10455
rect 3065 10421 3099 10455
rect 5089 10421 5123 10455
rect 5181 10421 5215 10455
rect 5733 10421 5767 10455
rect 6193 10421 6227 10455
rect 10609 10421 10643 10455
rect 12817 10421 12851 10455
rect 13921 10421 13955 10455
rect 14841 10421 14875 10455
rect 15209 10421 15243 10455
rect 15301 10421 15335 10455
rect 16313 10421 16347 10455
rect 1593 10217 1627 10251
rect 2053 10217 2087 10251
rect 2605 10217 2639 10251
rect 2973 10217 3007 10251
rect 5825 10217 5859 10251
rect 6101 10217 6135 10251
rect 8493 10217 8527 10251
rect 8585 10217 8619 10251
rect 12173 10217 12207 10251
rect 14289 10217 14323 10251
rect 14749 10217 14783 10251
rect 16681 10217 16715 10251
rect 1961 10149 1995 10183
rect 3065 10149 3099 10183
rect 15568 10149 15602 10183
rect 4712 10081 4746 10115
rect 6469 10081 6503 10115
rect 7481 10081 7515 10115
rect 10517 10081 10551 10115
rect 10784 10081 10818 10115
rect 12357 10081 12391 10115
rect 12633 10081 12667 10115
rect 12900 10081 12934 10115
rect 15301 10081 15335 10115
rect 2145 10013 2179 10047
rect 3249 10013 3283 10047
rect 4445 10013 4479 10047
rect 6561 10013 6595 10047
rect 6745 10013 6779 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8677 10013 8711 10047
rect 7113 9945 7147 9979
rect 11897 9945 11931 9979
rect 8125 9877 8159 9911
rect 14013 9877 14047 9911
rect 7481 9673 7515 9707
rect 4629 9605 4663 9639
rect 10057 9605 10091 9639
rect 13829 9605 13863 9639
rect 15117 9605 15151 9639
rect 3709 9537 3743 9571
rect 5273 9537 5307 9571
rect 6193 9537 6227 9571
rect 8033 9537 8067 9571
rect 11529 9537 11563 9571
rect 14565 9537 14599 9571
rect 14657 9537 14691 9571
rect 15761 9537 15795 9571
rect 2053 9469 2087 9503
rect 2320 9469 2354 9503
rect 7205 9469 7239 9503
rect 7941 9469 7975 9503
rect 8677 9469 8711 9503
rect 8944 9469 8978 9503
rect 11345 9469 11379 9503
rect 12449 9469 12483 9503
rect 15485 9469 15519 9503
rect 5089 9401 5123 9435
rect 6009 9401 6043 9435
rect 11253 9401 11287 9435
rect 11897 9401 11931 9435
rect 12694 9401 12728 9435
rect 3433 9333 3467 9367
rect 4997 9333 5031 9367
rect 5641 9333 5675 9367
rect 6101 9333 6135 9367
rect 7021 9333 7055 9367
rect 7849 9333 7883 9367
rect 10885 9333 10919 9367
rect 14105 9333 14139 9367
rect 14473 9333 14507 9367
rect 15577 9333 15611 9367
rect 2789 9129 2823 9163
rect 5089 9129 5123 9163
rect 5549 9129 5583 9163
rect 7205 9129 7239 9163
rect 8861 9129 8895 9163
rect 10241 9129 10275 9163
rect 11621 9129 11655 9163
rect 12541 9129 12575 9163
rect 14289 9129 14323 9163
rect 1676 9061 1710 9095
rect 7748 9061 7782 9095
rect 10057 9061 10091 9095
rect 1409 8993 1443 9027
rect 4445 8993 4479 9027
rect 4537 8993 4571 9027
rect 5733 8993 5767 9027
rect 5825 8993 5859 9027
rect 6092 8993 6126 9027
rect 4721 8925 4755 8959
rect 7481 8925 7515 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 10149 9061 10183 9095
rect 10701 9061 10735 9095
rect 11713 9061 11747 9095
rect 13001 9061 13035 9095
rect 10609 8993 10643 9027
rect 12909 8993 12943 9027
rect 14381 8993 14415 9027
rect 10885 8925 10919 8959
rect 11897 8925 11931 8959
rect 13093 8925 13127 8959
rect 14473 8925 14507 8959
rect 11253 8857 11287 8891
rect 4077 8789 4111 8823
rect 10149 8789 10183 8823
rect 13921 8789 13955 8823
rect 2881 8585 2915 8619
rect 5457 8585 5491 8619
rect 7297 8585 7331 8619
rect 10977 8585 11011 8619
rect 13277 8585 13311 8619
rect 8309 8517 8343 8551
rect 2145 8449 2179 8483
rect 3341 8449 3375 8483
rect 3433 8449 3467 8483
rect 4353 8449 4387 8483
rect 4537 8449 4571 8483
rect 6009 8449 6043 8483
rect 7757 8449 7791 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 8953 8449 8987 8483
rect 11437 8449 11471 8483
rect 11529 8449 11563 8483
rect 13737 8449 13771 8483
rect 13829 8449 13863 8483
rect 1961 8381 1995 8415
rect 5825 8381 5859 8415
rect 6653 8381 6687 8415
rect 7665 8381 7699 8415
rect 8677 8381 8711 8415
rect 9321 8381 9355 8415
rect 9588 8381 9622 8415
rect 12817 8381 12851 8415
rect 14289 8381 14323 8415
rect 3249 8313 3283 8347
rect 4261 8313 4295 8347
rect 4997 8313 5031 8347
rect 8217 8313 8251 8347
rect 13645 8313 13679 8347
rect 14556 8313 14590 8347
rect 3893 8245 3927 8279
rect 5917 8245 5951 8279
rect 6469 8245 6503 8279
rect 8769 8245 8803 8279
rect 10701 8245 10735 8279
rect 11345 8245 11379 8279
rect 12633 8245 12667 8279
rect 15669 8245 15703 8279
rect 6101 8041 6135 8075
rect 6377 8041 6411 8075
rect 6745 8041 6779 8075
rect 7941 8041 7975 8075
rect 8585 8041 8619 8075
rect 9689 8041 9723 8075
rect 14565 8041 14599 8075
rect 15669 8041 15703 8075
rect 15761 8041 15795 8075
rect 1777 7973 1811 8007
rect 2482 7973 2516 8007
rect 8033 7973 8067 8007
rect 1501 7905 1535 7939
rect 4988 7905 5022 7939
rect 8953 7905 8987 7939
rect 10057 7905 10091 7939
rect 10977 7905 11011 7939
rect 11428 7905 11462 7939
rect 13084 7905 13118 7939
rect 2237 7837 2271 7871
rect 4721 7837 4755 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 8217 7837 8251 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 11161 7837 11195 7871
rect 12817 7837 12851 7871
rect 15853 7837 15887 7871
rect 7573 7769 7607 7803
rect 10793 7769 10827 7803
rect 14197 7769 14231 7803
rect 3617 7701 3651 7735
rect 12541 7701 12575 7735
rect 15301 7701 15335 7735
rect 4445 7497 4479 7531
rect 5733 7497 5767 7531
rect 8217 7497 8251 7531
rect 8677 7497 8711 7531
rect 9689 7497 9723 7531
rect 1961 7361 1995 7395
rect 2973 7361 3007 7395
rect 3985 7361 4019 7395
rect 4997 7361 5031 7395
rect 6285 7361 6319 7395
rect 9321 7361 9355 7395
rect 10333 7361 10367 7395
rect 15025 7361 15059 7395
rect 6193 7293 6227 7327
rect 6844 7293 6878 7327
rect 9137 7293 9171 7327
rect 10701 7293 10735 7327
rect 10968 7293 11002 7327
rect 14013 7293 14047 7327
rect 14841 7293 14875 7327
rect 15485 7293 15519 7327
rect 15741 7293 15775 7327
rect 2881 7225 2915 7259
rect 3801 7225 3835 7259
rect 6101 7225 6135 7259
rect 7104 7225 7138 7259
rect 10149 7225 10183 7259
rect 1409 7157 1443 7191
rect 1777 7157 1811 7191
rect 1869 7157 1903 7191
rect 2421 7157 2455 7191
rect 2789 7157 2823 7191
rect 3433 7157 3467 7191
rect 3893 7157 3927 7191
rect 4813 7157 4847 7191
rect 4905 7157 4939 7191
rect 9045 7157 9079 7191
rect 10057 7157 10091 7191
rect 12081 7157 12115 7191
rect 13829 7157 13863 7191
rect 14473 7157 14507 7191
rect 14933 7157 14967 7191
rect 16865 7157 16899 7191
rect 5549 6953 5583 6987
rect 6193 6953 6227 6987
rect 8493 6953 8527 6987
rect 10701 6953 10735 6987
rect 13461 6953 13495 6987
rect 14657 6953 14691 6987
rect 15669 6953 15703 6987
rect 11704 6885 11738 6919
rect 14565 6885 14599 6919
rect 2320 6817 2354 6851
rect 4169 6817 4203 6851
rect 4436 6817 4470 6851
rect 6837 6817 6871 6851
rect 7104 6817 7138 6851
rect 8861 6817 8895 6851
rect 8953 6817 8987 6851
rect 10057 6817 10091 6851
rect 13553 6817 13587 6851
rect 19156 6817 19190 6851
rect 2053 6749 2087 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 9045 6749 9079 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 11345 6749 11379 6783
rect 11437 6749 11471 6783
rect 13737 6749 13771 6783
rect 14749 6749 14783 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 18889 6749 18923 6783
rect 14197 6681 14231 6715
rect 3433 6613 3467 6647
rect 5825 6613 5859 6647
rect 8217 6613 8251 6647
rect 9689 6613 9723 6647
rect 11345 6613 11379 6647
rect 12817 6613 12851 6647
rect 13093 6613 13127 6647
rect 15301 6613 15335 6647
rect 20269 6613 20303 6647
rect 1409 6409 1443 6443
rect 2421 6409 2455 6443
rect 3893 6409 3927 6443
rect 14197 6409 14231 6443
rect 4997 6341 5031 6375
rect 12449 6341 12483 6375
rect 2053 6273 2087 6307
rect 2973 6273 3007 6307
rect 4537 6273 4571 6307
rect 5549 6273 5583 6307
rect 8125 6273 8159 6307
rect 8493 6273 8527 6307
rect 11253 6273 11287 6307
rect 11345 6273 11379 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 17141 6273 17175 6307
rect 1777 6205 1811 6239
rect 1869 6205 1903 6239
rect 7941 6205 7975 6239
rect 9137 6205 9171 6239
rect 11161 6205 11195 6239
rect 17049 6205 17083 6239
rect 18981 6205 19015 6239
rect 2789 6137 2823 6171
rect 3433 6137 3467 6171
rect 5365 6137 5399 6171
rect 9404 6137 9438 6171
rect 19257 6137 19291 6171
rect 2881 6069 2915 6103
rect 4261 6069 4295 6103
rect 4353 6069 4387 6103
rect 5457 6069 5491 6103
rect 7481 6069 7515 6103
rect 7849 6069 7883 6103
rect 10517 6069 10551 6103
rect 10793 6069 10827 6103
rect 12817 6069 12851 6103
rect 14565 6069 14599 6103
rect 15209 6069 15243 6103
rect 15577 6069 15611 6103
rect 16589 6069 16623 6103
rect 16957 6069 16991 6103
rect 2789 5865 2823 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 6101 5865 6135 5899
rect 6561 5865 6595 5899
rect 6929 5865 6963 5899
rect 11069 5865 11103 5899
rect 14749 5865 14783 5899
rect 20269 5865 20303 5899
rect 1676 5797 1710 5831
rect 4537 5797 4571 5831
rect 5457 5729 5491 5763
rect 7941 5729 7975 5763
rect 9956 5729 9990 5763
rect 11713 5729 11747 5763
rect 13084 5729 13118 5763
rect 15844 5729 15878 5763
rect 17489 5729 17523 5763
rect 18797 5729 18831 5763
rect 19145 5729 19179 5763
rect 1409 5661 1443 5695
rect 4629 5661 4663 5695
rect 5549 5661 5583 5695
rect 5733 5661 5767 5695
rect 7021 5661 7055 5695
rect 7205 5661 7239 5695
rect 8033 5661 8067 5695
rect 8217 5661 8251 5695
rect 9689 5661 9723 5695
rect 11805 5661 11839 5695
rect 11989 5661 12023 5695
rect 12817 5661 12851 5695
rect 15577 5661 15611 5695
rect 17233 5661 17267 5695
rect 7573 5593 7607 5627
rect 18889 5661 18923 5695
rect 5089 5525 5123 5559
rect 11345 5525 11379 5559
rect 14197 5525 14231 5559
rect 16957 5525 16991 5559
rect 18613 5525 18647 5559
rect 18797 5525 18831 5559
rect 1777 5321 1811 5355
rect 4169 5321 4203 5355
rect 2329 5185 2363 5219
rect 9873 5185 9907 5219
rect 10977 5185 11011 5219
rect 11989 5185 12023 5219
rect 13001 5185 13035 5219
rect 17049 5185 17083 5219
rect 2789 5117 2823 5151
rect 3056 5117 3090 5151
rect 5089 5117 5123 5151
rect 7113 5117 7147 5151
rect 7380 5117 7414 5151
rect 9689 5117 9723 5151
rect 10701 5117 10735 5151
rect 14381 5117 14415 5151
rect 16865 5117 16899 5151
rect 19809 5117 19843 5151
rect 5356 5049 5390 5083
rect 12909 5049 12943 5083
rect 14648 5049 14682 5083
rect 17417 5049 17451 5083
rect 2145 4981 2179 5015
rect 2237 4981 2271 5015
rect 6469 4981 6503 5015
rect 8493 4981 8527 5015
rect 9321 4981 9355 5015
rect 9781 4981 9815 5015
rect 10333 4981 10367 5015
rect 10793 4981 10827 5015
rect 11345 4981 11379 5015
rect 11713 4981 11747 5015
rect 11805 4981 11839 5015
rect 12449 4981 12483 5015
rect 12817 4981 12851 5015
rect 15761 4981 15795 5015
rect 16405 4981 16439 5015
rect 16773 4981 16807 5015
rect 19993 4981 20027 5015
rect 7849 4777 7883 4811
rect 10241 4777 10275 4811
rect 10793 4777 10827 4811
rect 11805 4777 11839 4811
rect 15669 4777 15703 4811
rect 15761 4777 15795 4811
rect 16773 4777 16807 4811
rect 17325 4777 17359 4811
rect 2114 4709 2148 4743
rect 7757 4709 7791 4743
rect 13820 4709 13854 4743
rect 16681 4709 16715 4743
rect 1869 4641 1903 4675
rect 4344 4641 4378 4675
rect 6745 4641 6779 4675
rect 8769 4641 8803 4675
rect 10149 4641 10183 4675
rect 11161 4641 11195 4675
rect 12173 4641 12207 4675
rect 12265 4641 12299 4675
rect 17693 4641 17727 4675
rect 18337 4641 18371 4675
rect 4077 4573 4111 4607
rect 6837 4573 6871 4607
rect 6929 4573 6963 4607
rect 7941 4573 7975 4607
rect 8861 4573 8895 4607
rect 9045 4573 9079 4607
rect 10333 4573 10367 4607
rect 11253 4573 11287 4607
rect 11437 4573 11471 4607
rect 12357 4573 12391 4607
rect 13553 4573 13587 4607
rect 15853 4573 15887 4607
rect 16957 4573 16991 4607
rect 17785 4573 17819 4607
rect 17969 4573 18003 4607
rect 18521 4573 18555 4607
rect 5457 4505 5491 4539
rect 8401 4505 8435 4539
rect 16313 4505 16347 4539
rect 3249 4437 3283 4471
rect 6377 4437 6411 4471
rect 7389 4437 7423 4471
rect 9781 4437 9815 4471
rect 14933 4437 14967 4471
rect 15301 4437 15335 4471
rect 2513 4233 2547 4267
rect 8585 4233 8619 4267
rect 1501 4165 1535 4199
rect 15301 4165 15335 4199
rect 2053 4097 2087 4131
rect 3157 4097 3191 4131
rect 4261 4097 4295 4131
rect 5365 4097 5399 4131
rect 6377 4097 6411 4131
rect 7389 4097 7423 4131
rect 9045 4097 9079 4131
rect 9229 4097 9263 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 10425 4097 10459 4131
rect 11069 4097 11103 4131
rect 11253 4097 11287 4131
rect 13093 4097 13127 4131
rect 14933 4097 14967 4131
rect 15945 4097 15979 4131
rect 16865 4097 16899 4131
rect 2881 4029 2915 4063
rect 6101 4029 6135 4063
rect 7297 4029 7331 4063
rect 1869 3961 1903 3995
rect 8953 3961 8987 3995
rect 11621 4029 11655 4063
rect 12909 4029 12943 4063
rect 13461 4029 13495 4063
rect 16773 4029 16807 4063
rect 18061 4029 18095 4063
rect 10977 3961 11011 3995
rect 11897 3961 11931 3995
rect 15761 3961 15795 3995
rect 16681 3961 16715 3995
rect 1961 3893 1995 3927
rect 2973 3893 3007 3927
rect 3709 3893 3743 3927
rect 4077 3893 4111 3927
rect 4169 3893 4203 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 5181 3893 5215 3927
rect 5733 3893 5767 3927
rect 6193 3893 6227 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 9597 3893 9631 3927
rect 9965 3893 9999 3927
rect 10425 3893 10459 3927
rect 10609 3893 10643 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 13645 3893 13679 3927
rect 14289 3893 14323 3927
rect 14657 3893 14691 3927
rect 14749 3893 14783 3927
rect 15669 3893 15703 3927
rect 16313 3893 16347 3927
rect 18245 3893 18279 3927
rect 3065 3689 3099 3723
rect 4721 3689 4755 3723
rect 8493 3689 8527 3723
rect 8585 3689 8619 3723
rect 13001 3689 13035 3723
rect 14013 3689 14047 3723
rect 15301 3689 15335 3723
rect 7941 3621 7975 3655
rect 1685 3553 1719 3587
rect 1952 3553 1986 3587
rect 5089 3553 5123 3587
rect 5733 3553 5767 3587
rect 6000 3553 6034 3587
rect 11244 3621 11278 3655
rect 14105 3621 14139 3655
rect 15669 3621 15703 3655
rect 8953 3553 8987 3587
rect 10149 3553 10183 3587
rect 10977 3553 11011 3587
rect 15761 3553 15795 3587
rect 16313 3553 16347 3587
rect 16865 3553 16899 3587
rect 17417 3553 17451 3587
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 8493 3485 8527 3519
rect 9045 3485 9079 3519
rect 9229 3485 9263 3519
rect 10241 3485 10275 3519
rect 10333 3485 10367 3519
rect 13093 3485 13127 3519
rect 13185 3485 13219 3519
rect 14289 3485 14323 3519
rect 15853 3485 15887 3519
rect 12357 3417 12391 3451
rect 13645 3417 13679 3451
rect 17049 3417 17083 3451
rect 7113 3349 7147 3383
rect 7573 3349 7607 3383
rect 9781 3349 9815 3383
rect 12633 3349 12667 3383
rect 16497 3349 16531 3383
rect 17601 3349 17635 3383
rect 3433 3145 3467 3179
rect 5917 3145 5951 3179
rect 10885 3145 10919 3179
rect 12265 3145 12299 3179
rect 10609 3077 10643 3111
rect 10701 3077 10735 3111
rect 4537 3009 4571 3043
rect 7113 3009 7147 3043
rect 2053 2941 2087 2975
rect 4804 2941 4838 2975
rect 7380 2941 7414 2975
rect 9229 2941 9263 2975
rect 11437 3009 11471 3043
rect 16773 3077 16807 3111
rect 12541 2941 12575 2975
rect 12808 2941 12842 2975
rect 14197 2941 14231 2975
rect 15853 2941 15887 2975
rect 16589 2941 16623 2975
rect 17141 2941 17175 2975
rect 18061 2941 18095 2975
rect 18889 2941 18923 2975
rect 2320 2873 2354 2907
rect 9474 2873 9508 2907
rect 10701 2873 10735 2907
rect 11253 2873 11287 2907
rect 12265 2873 12299 2907
rect 14464 2873 14498 2907
rect 16129 2873 16163 2907
rect 3709 2805 3743 2839
rect 8493 2805 8527 2839
rect 11345 2805 11379 2839
rect 13921 2805 13955 2839
rect 15577 2805 15611 2839
rect 17325 2805 17359 2839
rect 18245 2805 18279 2839
rect 19073 2805 19107 2839
rect 1961 2601 1995 2635
rect 2329 2601 2363 2635
rect 3433 2601 3467 2635
rect 5457 2601 5491 2635
rect 7389 2601 7423 2635
rect 7941 2601 7975 2635
rect 8309 2601 8343 2635
rect 9873 2601 9907 2635
rect 10425 2601 10459 2635
rect 10885 2601 10919 2635
rect 11897 2601 11931 2635
rect 16221 2601 16255 2635
rect 16773 2601 16807 2635
rect 2421 2533 2455 2567
rect 5365 2533 5399 2567
rect 7297 2533 7331 2567
rect 10793 2533 10827 2567
rect 12909 2533 12943 2567
rect 2789 2465 2823 2499
rect 3341 2465 3375 2499
rect 6009 2465 6043 2499
rect 6285 2465 6319 2499
rect 8401 2465 8435 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 14289 2465 14323 2499
rect 15485 2465 15519 2499
rect 15853 2465 15887 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19441 2465 19475 2499
rect 20269 2465 20303 2499
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 3525 2397 3559 2431
rect 5641 2397 5675 2431
rect 7573 2397 7607 2431
rect 8585 2397 8619 2431
rect 10977 2397 11011 2431
rect 11989 2397 12023 2431
rect 14565 2397 14599 2431
rect 2973 2329 3007 2363
rect 4997 2329 5031 2363
rect 11437 2329 11471 2363
rect 15853 2329 15887 2363
rect 17325 2329 17359 2363
rect 6929 2261 6963 2295
rect 13553 2261 13587 2295
rect 15669 2261 15703 2295
rect 17877 2261 17911 2295
rect 18521 2261 18555 2295
rect 19073 2261 19107 2295
rect 19625 2261 19659 2295
rect 20453 2261 20487 2295
<< metal1 >>
rect 4246 21904 4252 21956
rect 4304 21944 4310 21956
rect 4614 21944 4620 21956
rect 4304 21916 4620 21944
rect 4304 21904 4310 21916
rect 4614 21904 4620 21916
rect 4672 21904 4678 21956
rect 6086 21904 6092 21956
rect 6144 21944 6150 21956
rect 6270 21944 6276 21956
rect 6144 21916 6276 21944
rect 6144 21904 6150 21916
rect 6270 21904 6276 21916
rect 6328 21904 6334 21956
rect 7098 20272 7104 20324
rect 7156 20312 7162 20324
rect 7926 20312 7932 20324
rect 7156 20284 7932 20312
rect 7156 20272 7162 20284
rect 7926 20272 7932 20284
rect 7984 20272 7990 20324
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 2774 20040 2780 20052
rect 2547 20012 2780 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3050 20040 3056 20052
rect 3011 20012 3056 20040
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3602 20040 3608 20052
rect 3563 20012 3608 20040
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 12894 20040 12900 20052
rect 12851 20012 12900 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19334 20040 19340 20052
rect 18739 20012 19340 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19521 20043 19579 20049
rect 19521 20009 19533 20043
rect 19567 20040 19579 20043
rect 20254 20040 20260 20052
rect 19567 20012 20260 20040
rect 19567 20009 19579 20012
rect 19521 20003 19579 20009
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 4982 19972 4988 19984
rect 2332 19944 4988 19972
rect 2332 19913 2360 19944
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 10229 19975 10287 19981
rect 10229 19941 10241 19975
rect 10275 19972 10287 19975
rect 13262 19972 13268 19984
rect 10275 19944 13268 19972
rect 10275 19941 10287 19944
rect 10229 19935 10287 19941
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 1780 19768 1808 19867
rect 2682 19864 2688 19916
rect 2740 19904 2746 19916
rect 2869 19907 2927 19913
rect 2869 19904 2881 19907
rect 2740 19876 2881 19904
rect 2740 19864 2746 19876
rect 2869 19873 2881 19876
rect 2915 19873 2927 19907
rect 2869 19867 2927 19873
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19873 3479 19907
rect 5902 19904 5908 19916
rect 5863 19876 5908 19904
rect 3421 19867 3479 19873
rect 2038 19796 2044 19848
rect 2096 19836 2102 19848
rect 3436 19836 3464 19867
rect 5902 19864 5908 19876
rect 5960 19864 5966 19916
rect 7742 19904 7748 19916
rect 7703 19876 7748 19904
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13630 19904 13636 19916
rect 13219 19876 13636 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 18598 19904 18604 19916
rect 18555 19876 18604 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 19334 19904 19340 19916
rect 19295 19876 19340 19904
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 4062 19836 4068 19848
rect 2096 19808 3464 19836
rect 4023 19808 4068 19836
rect 2096 19796 2102 19808
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 5994 19836 6000 19848
rect 5955 19808 6000 19836
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 6914 19836 6920 19848
rect 6227 19808 6920 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19836 8079 19839
rect 8202 19836 8208 19848
rect 8067 19808 8208 19836
rect 8067 19805 8079 19808
rect 8021 19799 8079 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 10321 19839 10379 19845
rect 10321 19836 10333 19839
rect 9916 19808 10333 19836
rect 9916 19796 9922 19808
rect 10321 19805 10333 19808
rect 10367 19805 10379 19839
rect 10321 19799 10379 19805
rect 9030 19768 9036 19780
rect 1780 19740 9036 19768
rect 9030 19728 9036 19740
rect 9088 19728 9094 19780
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 5534 19700 5540 19712
rect 5495 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 6362 19700 6368 19712
rect 5684 19672 6368 19700
rect 5684 19660 5690 19672
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 6822 19660 6828 19712
rect 6880 19700 6886 19712
rect 7377 19703 7435 19709
rect 7377 19700 7389 19703
rect 6880 19672 7389 19700
rect 6880 19660 6886 19672
rect 7377 19669 7389 19672
rect 7423 19669 7435 19703
rect 7377 19663 7435 19669
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 9769 19703 9827 19709
rect 9769 19700 9781 19703
rect 8904 19672 9781 19700
rect 8904 19660 8910 19672
rect 9769 19669 9781 19672
rect 9815 19669 9827 19703
rect 9769 19663 9827 19669
rect 13357 19703 13415 19709
rect 13357 19669 13369 19703
rect 13403 19700 13415 19703
rect 16666 19700 16672 19712
rect 13403 19672 16672 19700
rect 13403 19669 13415 19672
rect 13357 19663 13415 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3326 19496 3332 19508
rect 3287 19468 3332 19496
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 7834 19496 7840 19508
rect 4908 19468 5948 19496
rect 7795 19468 7840 19496
rect 2866 19388 2872 19440
rect 2924 19428 2930 19440
rect 4908 19428 4936 19468
rect 2924 19400 4936 19428
rect 2924 19388 2930 19400
rect 2682 19360 2688 19372
rect 2643 19332 2688 19360
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19261 1731 19295
rect 1673 19255 1731 19261
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19292 2007 19295
rect 2038 19292 2044 19304
rect 1995 19264 2044 19292
rect 1995 19261 2007 19264
rect 1949 19255 2007 19261
rect 1688 19156 1716 19255
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19261 2467 19295
rect 3142 19292 3148 19304
rect 3103 19264 3148 19292
rect 2409 19255 2467 19261
rect 2424 19224 2452 19255
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 2424 19196 3740 19224
rect 2866 19156 2872 19168
rect 1688 19128 2872 19156
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 3712 19165 3740 19196
rect 3786 19184 3792 19236
rect 3844 19224 3850 19236
rect 4356 19224 4384 19323
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4856 19264 4905 19292
rect 4856 19252 4862 19264
rect 4893 19261 4905 19264
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5920 19292 5948 19468
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 6086 19388 6092 19440
rect 6144 19428 6150 19440
rect 6270 19428 6276 19440
rect 6144 19400 6276 19428
rect 6144 19388 6150 19400
rect 6270 19388 6276 19400
rect 6328 19388 6334 19440
rect 10965 19431 11023 19437
rect 10965 19397 10977 19431
rect 11011 19397 11023 19431
rect 10965 19391 11023 19397
rect 8481 19363 8539 19369
rect 6656 19332 6960 19360
rect 6656 19292 6684 19332
rect 6822 19292 6828 19304
rect 5040 19264 5580 19292
rect 5920 19264 6684 19292
rect 6783 19264 6828 19292
rect 5040 19252 5046 19264
rect 3844 19196 4384 19224
rect 3844 19184 3850 19196
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19125 3755 19159
rect 4154 19156 4160 19168
rect 4115 19128 4160 19156
rect 3697 19119 3755 19125
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4356 19156 4384 19196
rect 5160 19227 5218 19233
rect 5160 19193 5172 19227
rect 5206 19224 5218 19227
rect 5442 19224 5448 19236
rect 5206 19196 5448 19224
rect 5206 19193 5218 19196
rect 5160 19187 5218 19193
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 5552 19224 5580 19264
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 6932 19292 6960 19332
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 9030 19360 9036 19372
rect 8991 19332 9036 19360
rect 8481 19323 8539 19329
rect 6932 19264 7604 19292
rect 7101 19227 7159 19233
rect 7101 19224 7113 19227
rect 5552 19196 7113 19224
rect 7101 19193 7113 19196
rect 7147 19193 7159 19227
rect 7576 19224 7604 19264
rect 7650 19252 7656 19304
rect 7708 19292 7714 19304
rect 8496 19292 8524 19323
rect 9030 19320 9036 19332
rect 9088 19320 9094 19372
rect 8846 19292 8852 19304
rect 7708 19264 8616 19292
rect 8807 19264 8852 19292
rect 7708 19252 7714 19264
rect 8478 19224 8484 19236
rect 7576 19196 8484 19224
rect 7101 19187 7159 19193
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 8588 19224 8616 19264
rect 8846 19252 8852 19264
rect 8904 19252 8910 19304
rect 8956 19264 9260 19292
rect 8956 19224 8984 19264
rect 8588 19196 8984 19224
rect 9232 19224 9260 19264
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 9548 19264 9597 19292
rect 9548 19252 9554 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 10980 19292 11008 19391
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12216 19332 12940 19360
rect 12216 19320 12222 19332
rect 9585 19255 9643 19261
rect 9692 19264 11008 19292
rect 11517 19295 11575 19301
rect 9692 19224 9720 19264
rect 11517 19261 11529 19295
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12618 19292 12624 19304
rect 11839 19264 12624 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 9858 19233 9864 19236
rect 9852 19224 9864 19233
rect 9232 19196 9720 19224
rect 9819 19196 9864 19224
rect 9852 19187 9864 19196
rect 9858 19184 9864 19187
rect 9916 19184 9922 19236
rect 11532 19224 11560 19255
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 12768 19264 12813 19292
rect 12768 19252 12774 19264
rect 11882 19224 11888 19236
rect 10888 19196 11100 19224
rect 11532 19196 11888 19224
rect 6273 19159 6331 19165
rect 6273 19156 6285 19159
rect 4356 19128 6285 19156
rect 6273 19125 6285 19128
rect 6319 19125 6331 19159
rect 6273 19119 6331 19125
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 7616 19128 8217 19156
rect 7616 19116 7622 19128
rect 8205 19125 8217 19128
rect 8251 19125 8263 19159
rect 8205 19119 8263 19125
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 10888 19156 10916 19196
rect 8343 19128 10916 19156
rect 11072 19156 11100 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 11974 19184 11980 19236
rect 12032 19224 12038 19236
rect 12802 19224 12808 19236
rect 12032 19196 12808 19224
rect 12032 19184 12038 19196
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 12912 19224 12940 19332
rect 16684 19332 17080 19360
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 13035 19264 13461 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 14090 19292 14096 19304
rect 14047 19264 14096 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14516 19264 14565 19292
rect 14516 19252 14522 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 15102 19292 15108 19304
rect 15063 19264 15108 19292
rect 14553 19255 14611 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15470 19252 15476 19304
rect 15528 19292 15534 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15528 19264 15669 19292
rect 15528 19252 15534 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 16206 19292 16212 19304
rect 16167 19264 16212 19292
rect 15657 19255 15715 19261
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16684 19292 16712 19332
rect 16316 19264 16712 19292
rect 16761 19295 16819 19301
rect 16316 19224 16344 19264
rect 16761 19261 16773 19295
rect 16807 19292 16819 19295
rect 16942 19292 16948 19304
rect 16807 19264 16948 19292
rect 16807 19261 16819 19264
rect 16761 19255 16819 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17052 19292 17080 19332
rect 17052 19264 17172 19292
rect 17034 19224 17040 19236
rect 12912 19196 16344 19224
rect 16408 19196 17040 19224
rect 12434 19156 12440 19168
rect 11072 19128 12440 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13412 19128 13645 19156
rect 13412 19116 13418 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 14185 19159 14243 19165
rect 14185 19125 14197 19159
rect 14231 19156 14243 19159
rect 14274 19156 14280 19168
rect 14231 19128 14280 19156
rect 14231 19125 14243 19128
rect 14185 19119 14243 19125
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 14737 19159 14795 19165
rect 14737 19125 14749 19159
rect 14783 19156 14795 19159
rect 15194 19156 15200 19168
rect 14783 19128 15200 19156
rect 14783 19125 14795 19128
rect 14737 19119 14795 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15654 19156 15660 19168
rect 15335 19128 15660 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 15841 19159 15899 19165
rect 15841 19125 15853 19159
rect 15887 19156 15899 19159
rect 16114 19156 16120 19168
rect 15887 19128 16120 19156
rect 15887 19125 15899 19128
rect 15841 19119 15899 19125
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16408 19165 16436 19196
rect 17034 19184 17040 19196
rect 17092 19184 17098 19236
rect 17144 19224 17172 19264
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 17276 19264 17325 19292
rect 17276 19252 17282 19264
rect 17313 19261 17325 19264
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17552 19264 18061 19292
rect 17552 19252 17558 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19292 19303 19295
rect 19291 19264 20300 19292
rect 19291 19261 19303 19264
rect 19245 19255 19303 19261
rect 19889 19227 19947 19233
rect 19889 19224 19901 19227
rect 17144 19196 19901 19224
rect 19889 19193 19901 19196
rect 19935 19193 19947 19227
rect 20272 19224 20300 19264
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 20404 19264 20449 19292
rect 20404 19252 20410 19264
rect 22094 19224 22100 19236
rect 20272 19196 22100 19224
rect 19889 19187 19947 19193
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 16393 19159 16451 19165
rect 16393 19125 16405 19159
rect 16439 19125 16451 19159
rect 16393 19119 16451 19125
rect 16945 19159 17003 19165
rect 16945 19125 16957 19159
rect 16991 19156 17003 19159
rect 17402 19156 17408 19168
rect 16991 19128 17408 19156
rect 16991 19125 17003 19128
rect 16945 19119 17003 19125
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17497 19159 17555 19165
rect 17497 19125 17509 19159
rect 17543 19156 17555 19159
rect 17954 19156 17960 19168
rect 17543 19128 17960 19156
rect 17543 19125 17555 19128
rect 17497 19119 17555 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 20533 19159 20591 19165
rect 20533 19125 20545 19159
rect 20579 19156 20591 19159
rect 20714 19156 20720 19168
rect 20579 19128 20720 19156
rect 20579 19125 20591 19128
rect 20533 19119 20591 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 3467 18924 5672 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 2317 18887 2375 18893
rect 2317 18853 2329 18887
rect 2363 18884 2375 18887
rect 3142 18884 3148 18896
rect 2363 18856 3148 18884
rect 2363 18853 2375 18856
rect 2317 18847 2375 18853
rect 3142 18844 3148 18856
rect 3200 18844 3206 18896
rect 5534 18884 5540 18896
rect 3252 18856 4108 18884
rect 1489 18819 1547 18825
rect 1489 18785 1501 18819
rect 1535 18816 1547 18819
rect 1946 18816 1952 18828
rect 1535 18788 1952 18816
rect 1535 18785 1547 18788
rect 1489 18779 1547 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 1670 18680 1676 18692
rect 1631 18652 1676 18680
rect 1670 18640 1676 18652
rect 1728 18640 1734 18692
rect 2056 18680 2084 18779
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 3252 18816 3280 18856
rect 2832 18788 3280 18816
rect 3329 18819 3387 18825
rect 2832 18776 2838 18788
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 3878 18816 3884 18828
rect 3375 18788 3884 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 3878 18776 3884 18788
rect 3936 18776 3942 18828
rect 4080 18825 4108 18856
rect 4172 18856 5540 18884
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 3694 18748 3700 18760
rect 3651 18720 3700 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 4172 18748 4200 18856
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 5644 18884 5672 18924
rect 5902 18912 5908 18964
rect 5960 18952 5966 18964
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 5960 18924 6469 18952
rect 5960 18912 5966 18924
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6457 18915 6515 18921
rect 6917 18955 6975 18961
rect 6917 18921 6929 18955
rect 6963 18952 6975 18955
rect 7742 18952 7748 18964
rect 6963 18924 7748 18952
rect 6963 18921 6975 18924
rect 6917 18915 6975 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 9674 18952 9680 18964
rect 8536 18924 9680 18952
rect 8536 18912 8542 18924
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 9916 18924 11069 18952
rect 9916 18912 9922 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 12618 18952 12624 18964
rect 11057 18915 11115 18921
rect 11624 18924 12624 18952
rect 7006 18884 7012 18896
rect 5644 18856 7012 18884
rect 7006 18844 7012 18856
rect 7064 18844 7070 18896
rect 7650 18893 7656 18896
rect 7644 18884 7656 18893
rect 7611 18856 7656 18884
rect 7644 18847 7656 18856
rect 7650 18844 7656 18847
rect 7708 18844 7714 18896
rect 8018 18844 8024 18896
rect 8076 18884 8082 18896
rect 9490 18884 9496 18896
rect 8076 18856 9496 18884
rect 8076 18844 8082 18856
rect 9490 18844 9496 18856
rect 9548 18844 9554 18896
rect 11624 18884 11652 18924
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14608 18924 14749 18952
rect 14608 18912 14614 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 14737 18915 14795 18921
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16574 18952 16580 18964
rect 16255 18924 16580 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 18233 18955 18291 18961
rect 18233 18921 18245 18955
rect 18279 18952 18291 18955
rect 18874 18952 18880 18964
rect 18279 18924 18880 18952
rect 18279 18921 18291 18924
rect 18233 18915 18291 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19153 18955 19211 18961
rect 19153 18921 19165 18955
rect 19199 18952 19211 18955
rect 19794 18952 19800 18964
rect 19199 18924 19800 18952
rect 19199 18921 19211 18924
rect 19153 18915 19211 18921
rect 19794 18912 19800 18924
rect 19852 18912 19858 18964
rect 9876 18856 11652 18884
rect 11876 18887 11934 18893
rect 5068 18819 5126 18825
rect 5068 18785 5080 18819
rect 5114 18816 5126 18819
rect 6914 18816 6920 18828
rect 5114 18788 6920 18816
rect 5114 18785 5126 18788
rect 5068 18779 5126 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 9876 18816 9904 18856
rect 11876 18853 11888 18887
rect 11922 18884 11934 18887
rect 12526 18884 12532 18896
rect 11922 18856 12532 18884
rect 11922 18853 11934 18856
rect 11876 18847 11934 18853
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 12710 18844 12716 18896
rect 12768 18884 12774 18896
rect 13998 18884 14004 18896
rect 12768 18856 14004 18884
rect 12768 18844 12774 18856
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 15102 18884 15108 18896
rect 14240 18856 15108 18884
rect 14240 18844 14246 18856
rect 15102 18844 15108 18856
rect 15160 18844 15166 18896
rect 16666 18844 16672 18896
rect 16724 18884 16730 18896
rect 21634 18884 21640 18896
rect 16724 18856 21640 18884
rect 16724 18844 16730 18856
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 7300 18788 9904 18816
rect 9944 18819 10002 18825
rect 4080 18720 4200 18748
rect 4080 18680 4108 18720
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 4798 18748 4804 18760
rect 4396 18720 4804 18748
rect 4396 18708 4402 18720
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 4246 18680 4252 18692
rect 2056 18652 4108 18680
rect 4207 18652 4252 18680
rect 4246 18640 4252 18652
rect 4304 18640 4310 18692
rect 7300 18680 7328 18788
rect 9944 18785 9956 18819
rect 9990 18816 10002 18819
rect 10318 18816 10324 18828
rect 9990 18788 10324 18816
rect 9990 18785 10002 18788
rect 9944 18779 10002 18785
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 12342 18816 12348 18828
rect 11655 18788 12348 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 13446 18776 13452 18828
rect 13504 18816 13510 18828
rect 13630 18816 13636 18828
rect 13504 18788 13636 18816
rect 13504 18776 13510 18788
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18816 13783 18819
rect 14553 18819 14611 18825
rect 13771 18788 14228 18816
rect 13771 18785 13783 18788
rect 13725 18779 13783 18785
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18717 7435 18751
rect 9122 18748 9128 18760
rect 9083 18720 9128 18748
rect 7377 18711 7435 18717
rect 5736 18652 7328 18680
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 5736 18612 5764 18652
rect 3292 18584 5764 18612
rect 3292 18572 3298 18584
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 6181 18615 6239 18621
rect 6181 18612 6193 18615
rect 5868 18584 6193 18612
rect 5868 18572 5874 18584
rect 6181 18581 6193 18584
rect 6227 18581 6239 18615
rect 6181 18575 6239 18581
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 7392 18612 7420 18711
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9684 18751 9742 18757
rect 9684 18748 9696 18751
rect 9548 18720 9696 18748
rect 9548 18708 9554 18720
rect 9684 18717 9696 18720
rect 9730 18717 9742 18751
rect 9684 18711 9742 18717
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 13740 18748 13768 18779
rect 12860 18720 13768 18748
rect 13817 18751 13875 18757
rect 12860 18708 12866 18720
rect 13817 18717 13829 18751
rect 13863 18717 13875 18751
rect 13817 18711 13875 18717
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13832 18680 13860 18711
rect 13035 18652 13860 18680
rect 14200 18680 14228 18788
rect 14553 18785 14565 18819
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 15289 18819 15347 18825
rect 15289 18785 15301 18819
rect 15335 18816 15347 18819
rect 16022 18816 16028 18828
rect 15335 18788 15884 18816
rect 15983 18788 16028 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 14568 18748 14596 18779
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 14568 18720 15485 18748
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15856 18748 15884 18788
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16390 18776 16396 18828
rect 16448 18816 16454 18828
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 16448 18788 18061 18816
rect 16448 18776 16454 18788
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18966 18816 18972 18828
rect 18927 18788 18972 18816
rect 18049 18779 18107 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 16298 18748 16304 18760
rect 15856 18720 16304 18748
rect 15473 18711 15531 18717
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 15930 18680 15936 18692
rect 14200 18652 15936 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 8018 18612 8024 18624
rect 7340 18584 8024 18612
rect 7340 18572 7346 18584
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 8757 18615 8815 18621
rect 8757 18612 8769 18615
rect 8168 18584 8769 18612
rect 8168 18572 8174 18584
rect 8757 18581 8769 18584
rect 8803 18581 8815 18615
rect 8757 18575 8815 18581
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 13004 18612 13032 18643
rect 15930 18640 15936 18652
rect 15988 18640 15994 18692
rect 10376 18584 13032 18612
rect 10376 18572 10382 18584
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1486 18368 1492 18420
rect 1544 18408 1550 18420
rect 2498 18408 2504 18420
rect 1544 18380 2504 18408
rect 1544 18368 1550 18380
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 3694 18408 3700 18420
rect 3436 18380 3700 18408
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 1946 18204 1952 18216
rect 1903 18176 1952 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 3436 18204 3464 18380
rect 3694 18368 3700 18380
rect 3752 18408 3758 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 3752 18380 4905 18408
rect 3752 18368 3758 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5721 18411 5779 18417
rect 5721 18377 5733 18411
rect 5767 18408 5779 18411
rect 5994 18408 6000 18420
rect 5767 18380 6000 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18408 9735 18411
rect 10134 18408 10140 18420
rect 9723 18380 10140 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14185 18411 14243 18417
rect 14185 18408 14197 18411
rect 13872 18380 14197 18408
rect 13872 18368 13878 18380
rect 14185 18377 14197 18380
rect 14231 18377 14243 18411
rect 14185 18371 14243 18377
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 22554 18408 22560 18420
rect 15344 18380 22560 18408
rect 15344 18368 15350 18380
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 6549 18343 6607 18349
rect 6549 18340 6561 18343
rect 6196 18312 6561 18340
rect 6196 18281 6224 18312
rect 6549 18309 6561 18312
rect 6595 18309 6607 18343
rect 6549 18303 6607 18309
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 7340 18312 7420 18340
rect 7340 18300 7346 18312
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 6365 18275 6423 18281
rect 6365 18241 6377 18275
rect 6411 18272 6423 18275
rect 6822 18272 6828 18284
rect 6411 18244 6828 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 7392 18281 7420 18312
rect 8570 18300 8576 18352
rect 8628 18340 8634 18352
rect 10042 18340 10048 18352
rect 8628 18312 10048 18340
rect 8628 18300 8634 18312
rect 10042 18300 10048 18312
rect 10100 18300 10106 18352
rect 10594 18300 10600 18352
rect 10652 18340 10658 18352
rect 12158 18340 12164 18352
rect 10652 18312 12164 18340
rect 10652 18300 10658 18312
rect 12158 18300 12164 18312
rect 12216 18300 12222 18352
rect 12897 18343 12955 18349
rect 12897 18309 12909 18343
rect 12943 18340 12955 18343
rect 21174 18340 21180 18352
rect 12943 18312 21180 18340
rect 12943 18309 12955 18312
rect 12897 18303 12955 18309
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 10318 18272 10324 18284
rect 8536 18244 10180 18272
rect 10279 18244 10324 18272
rect 8536 18232 8542 18244
rect 2608 18176 3464 18204
rect 3513 18207 3571 18213
rect 2124 18139 2182 18145
rect 2124 18105 2136 18139
rect 2170 18136 2182 18139
rect 2608 18136 2636 18176
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 4246 18204 4252 18216
rect 3559 18176 4252 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 7282 18204 7288 18216
rect 4764 18176 7288 18204
rect 4764 18164 4770 18176
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 7644 18207 7702 18213
rect 7644 18173 7656 18207
rect 7690 18204 7702 18207
rect 8110 18204 8116 18216
rect 7690 18176 8116 18204
rect 7690 18173 7702 18176
rect 7644 18167 7702 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 9180 18176 10057 18204
rect 9180 18164 9186 18176
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10152 18204 10180 18244
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 12526 18272 12532 18284
rect 11471 18244 12532 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18272 15347 18275
rect 16022 18272 16028 18284
rect 15335 18244 16028 18272
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18272 16911 18275
rect 17494 18272 17500 18284
rect 16899 18244 17500 18272
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 19334 18272 19340 18284
rect 18739 18244 19340 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 12250 18204 12256 18216
rect 10152 18176 12256 18204
rect 10045 18167 10103 18173
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12713 18207 12771 18213
rect 12713 18173 12725 18207
rect 12759 18204 12771 18207
rect 12894 18204 12900 18216
rect 12759 18176 12900 18204
rect 12759 18173 12771 18176
rect 12713 18167 12771 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13587 18176 14013 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 15010 18204 15016 18216
rect 14971 18176 15016 18204
rect 14001 18167 14059 18173
rect 3786 18145 3792 18148
rect 2170 18108 2636 18136
rect 2170 18105 2182 18108
rect 2124 18099 2182 18105
rect 3780 18099 3792 18145
rect 3844 18136 3850 18148
rect 6549 18139 6607 18145
rect 3844 18108 3880 18136
rect 3786 18096 3792 18099
rect 3844 18096 3850 18108
rect 6549 18105 6561 18139
rect 6595 18136 6607 18139
rect 10686 18136 10692 18148
rect 6595 18108 10692 18136
rect 6595 18105 6607 18108
rect 6549 18099 6607 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 11606 18096 11612 18148
rect 11664 18136 11670 18148
rect 13078 18136 13084 18148
rect 11664 18108 13084 18136
rect 11664 18096 11670 18108
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 13280 18136 13308 18167
rect 15010 18164 15016 18176
rect 15068 18164 15074 18216
rect 16577 18207 16635 18213
rect 16577 18173 16589 18207
rect 16623 18173 16635 18207
rect 18414 18204 18420 18216
rect 18375 18176 18420 18204
rect 16577 18167 16635 18173
rect 13814 18136 13820 18148
rect 13280 18108 13820 18136
rect 13814 18096 13820 18108
rect 13872 18096 13878 18148
rect 16592 18136 16620 18167
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 16850 18136 16856 18148
rect 16592 18108 16856 18136
rect 16850 18096 16856 18108
rect 16908 18096 16914 18148
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 3050 18068 3056 18080
rect 1443 18040 3056 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 4856 18040 6101 18068
rect 4856 18028 4862 18040
rect 6089 18037 6101 18040
rect 6135 18037 6147 18071
rect 6089 18031 6147 18037
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 8757 18071 8815 18077
rect 8757 18068 8769 18071
rect 6880 18040 8769 18068
rect 6880 18028 6886 18040
rect 8757 18037 8769 18040
rect 8803 18037 8815 18071
rect 8757 18031 8815 18037
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 9950 18068 9956 18080
rect 9364 18040 9956 18068
rect 9364 18028 9370 18040
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10137 18071 10195 18077
rect 10137 18037 10149 18071
rect 10183 18068 10195 18071
rect 10318 18068 10324 18080
rect 10183 18040 10324 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11146 18068 11152 18080
rect 11107 18040 11152 18068
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11241 18071 11299 18077
rect 11241 18037 11253 18071
rect 11287 18068 11299 18071
rect 12802 18068 12808 18080
rect 11287 18040 12808 18068
rect 11287 18037 11299 18040
rect 11241 18031 11299 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 2866 17864 2872 17876
rect 2827 17836 2872 17864
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3016 17836 3341 17864
rect 3016 17824 3022 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4212 17836 4997 17864
rect 4212 17824 4218 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 4985 17827 5043 17833
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7929 17867 7987 17873
rect 7929 17864 7941 17867
rect 6972 17836 7941 17864
rect 6972 17824 6978 17836
rect 7929 17833 7941 17836
rect 7975 17833 7987 17867
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 7929 17827 7987 17833
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 12526 17864 12532 17876
rect 12487 17836 12532 17864
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12802 17864 12808 17876
rect 12763 17836 12808 17864
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13814 17864 13820 17876
rect 13775 17836 13820 17864
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 2317 17799 2375 17805
rect 2317 17765 2329 17799
rect 2363 17796 2375 17799
rect 2774 17796 2780 17808
rect 2363 17768 2780 17796
rect 2363 17765 2375 17768
rect 2317 17759 2375 17765
rect 2774 17756 2780 17768
rect 2832 17756 2838 17808
rect 3050 17756 3056 17808
rect 3108 17796 3114 17808
rect 3237 17799 3295 17805
rect 3237 17796 3249 17799
rect 3108 17768 3249 17796
rect 3108 17756 3114 17768
rect 3237 17765 3249 17768
rect 3283 17765 3295 17799
rect 3237 17759 3295 17765
rect 5442 17756 5448 17808
rect 5500 17756 5506 17808
rect 6822 17805 6828 17808
rect 6816 17796 6828 17805
rect 6783 17768 6828 17796
rect 6816 17759 6828 17768
rect 6822 17756 6828 17759
rect 6880 17756 6886 17808
rect 8754 17796 8760 17808
rect 7116 17768 8760 17796
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17728 1547 17731
rect 1762 17728 1768 17740
rect 1535 17700 1768 17728
rect 1535 17697 1547 17700
rect 1489 17691 1547 17697
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 1854 17688 1860 17740
rect 1912 17728 1918 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1912 17700 2053 17728
rect 1912 17688 1918 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 3142 17688 3148 17740
rect 3200 17728 3206 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3200 17700 4077 17728
rect 3200 17688 3206 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 5350 17728 5356 17740
rect 5311 17700 5356 17728
rect 4065 17691 4123 17697
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 5460 17728 5488 17756
rect 7116 17728 7144 17768
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 10042 17796 10048 17808
rect 10003 17768 10048 17796
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 11790 17756 11796 17808
rect 11848 17756 11854 17808
rect 13078 17756 13084 17808
rect 13136 17796 13142 17808
rect 13265 17799 13323 17805
rect 13265 17796 13277 17799
rect 13136 17768 13277 17796
rect 13136 17756 13142 17768
rect 13265 17765 13277 17768
rect 13311 17796 13323 17799
rect 13630 17796 13636 17808
rect 13311 17768 13636 17796
rect 13311 17765 13323 17768
rect 13265 17759 13323 17765
rect 13630 17756 13636 17768
rect 13688 17756 13694 17808
rect 5460 17700 5580 17728
rect 3234 17620 3240 17672
rect 3292 17660 3298 17672
rect 3421 17663 3479 17669
rect 3421 17660 3433 17663
rect 3292 17632 3433 17660
rect 3292 17620 3298 17632
rect 3421 17629 3433 17632
rect 3467 17629 3479 17663
rect 5258 17660 5264 17672
rect 3421 17623 3479 17629
rect 3528 17632 5264 17660
rect 1026 17552 1032 17604
rect 1084 17592 1090 17604
rect 3528 17592 3556 17632
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5552 17669 5580 17700
rect 5644 17700 7144 17728
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 1084 17564 3556 17592
rect 1084 17552 1090 17564
rect 3602 17552 3608 17604
rect 3660 17592 3666 17604
rect 4249 17595 4307 17601
rect 4249 17592 4261 17595
rect 3660 17564 4261 17592
rect 3660 17552 3666 17564
rect 4249 17561 4261 17564
rect 4295 17561 4307 17595
rect 5460 17592 5488 17623
rect 5644 17592 5672 17700
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 8665 17731 8723 17737
rect 8665 17728 8677 17731
rect 7340 17700 8677 17728
rect 7340 17688 7346 17700
rect 8665 17697 8677 17700
rect 8711 17697 8723 17731
rect 8665 17691 8723 17697
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 10778 17728 10784 17740
rect 9815 17700 10784 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 11416 17731 11474 17737
rect 11416 17697 11428 17731
rect 11462 17728 11474 17731
rect 11808 17728 11836 17756
rect 11462 17700 12204 17728
rect 11462 17697 11474 17700
rect 11416 17691 11474 17697
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 5868 17632 6561 17660
rect 5868 17620 5874 17632
rect 6549 17629 6561 17632
rect 6595 17629 6607 17663
rect 6549 17623 6607 17629
rect 8754 17620 8760 17672
rect 8812 17660 8818 17672
rect 11149 17663 11207 17669
rect 8812 17632 8857 17660
rect 8812 17620 8818 17632
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 12176 17660 12204 17700
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 13173 17731 13231 17737
rect 13173 17728 13185 17731
rect 12952 17700 13185 17728
rect 12952 17688 12958 17700
rect 13173 17697 13185 17700
rect 13219 17697 13231 17731
rect 13173 17691 13231 17697
rect 14185 17731 14243 17737
rect 14185 17697 14197 17731
rect 14231 17728 14243 17731
rect 16114 17728 16120 17740
rect 14231 17700 16120 17728
rect 14231 17697 14243 17700
rect 14185 17691 14243 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12176 17632 13369 17660
rect 11149 17623 11207 17629
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 13357 17623 13415 17629
rect 5460 17564 5672 17592
rect 4249 17555 4307 17561
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 7742 17524 7748 17536
rect 3936 17496 7748 17524
rect 3936 17484 3942 17496
rect 7742 17484 7748 17496
rect 7800 17484 7806 17536
rect 8202 17524 8208 17536
rect 8163 17496 8208 17524
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10778 17524 10784 17536
rect 9732 17496 10784 17524
rect 9732 17484 9738 17496
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 11164 17524 11192 17623
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 14424 17632 14469 17660
rect 14424 17620 14430 17632
rect 12342 17524 12348 17536
rect 11164 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 16390 17524 16396 17536
rect 12768 17496 16396 17524
rect 12768 17484 12774 17496
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1854 17320 1860 17332
rect 1815 17292 1860 17320
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 8202 17320 8208 17332
rect 2332 17292 8208 17320
rect 2332 17193 2360 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 11333 17323 11391 17329
rect 8628 17292 11284 17320
rect 8628 17280 8634 17292
rect 5905 17255 5963 17261
rect 5905 17221 5917 17255
rect 5951 17252 5963 17255
rect 6178 17252 6184 17264
rect 5951 17224 6184 17252
rect 5951 17221 5963 17224
rect 5905 17215 5963 17221
rect 6178 17212 6184 17224
rect 6236 17252 6242 17264
rect 8754 17252 8760 17264
rect 6236 17224 8760 17252
rect 6236 17212 6242 17224
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2317 17147 2375 17153
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 3970 17144 3976 17196
rect 4028 17184 4034 17196
rect 4246 17184 4252 17196
rect 4028 17156 4252 17184
rect 4028 17144 4034 17156
rect 4246 17144 4252 17156
rect 4304 17184 4310 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4304 17156 4537 17184
rect 4304 17144 4310 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4525 17147 4583 17153
rect 7098 17144 7104 17196
rect 7156 17184 7162 17196
rect 7374 17184 7380 17196
rect 7156 17156 7380 17184
rect 7156 17144 7162 17156
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8570 17184 8576 17196
rect 8251 17156 8576 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 11256 17184 11284 17292
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11790 17320 11796 17332
rect 11379 17292 11796 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 15102 17320 15108 17332
rect 12483 17292 15108 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 12986 17184 12992 17196
rect 9631 17156 10088 17184
rect 11256 17156 11836 17184
rect 12947 17156 12992 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2866 17116 2872 17128
rect 2004 17088 2872 17116
rect 2004 17076 2010 17088
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 2958 17076 2964 17128
rect 3016 17116 3022 17128
rect 4433 17119 4491 17125
rect 4433 17116 4445 17119
rect 3016 17088 4445 17116
rect 3016 17076 3022 17088
rect 4433 17085 4445 17088
rect 4479 17085 4491 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 4433 17079 4491 17085
rect 4540 17088 6193 17116
rect 3136 17051 3194 17057
rect 3136 17017 3148 17051
rect 3182 17048 3194 17051
rect 3234 17048 3240 17060
rect 3182 17020 3240 17048
rect 3182 17017 3194 17020
rect 3136 17011 3194 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 4540 17048 4568 17088
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9548 17088 9965 17116
rect 9548 17076 9554 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 4080 17020 4568 17048
rect 2225 16983 2283 16989
rect 2225 16949 2237 16983
rect 2271 16980 2283 16983
rect 2685 16983 2743 16989
rect 2685 16980 2697 16983
rect 2271 16952 2697 16980
rect 2271 16949 2283 16952
rect 2225 16943 2283 16949
rect 2685 16949 2697 16952
rect 2731 16949 2743 16983
rect 2685 16943 2743 16949
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 4080 16980 4108 17020
rect 4706 17008 4712 17060
rect 4764 17057 4770 17060
rect 4764 17051 4828 17057
rect 4764 17017 4782 17051
rect 4816 17017 4828 17051
rect 4764 17011 4828 17017
rect 4764 17008 4770 17011
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 10060 17048 10088 17156
rect 11808 17128 11836 17156
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 13906 17076 13912 17128
rect 13964 17116 13970 17128
rect 14366 17125 14372 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13964 17088 14105 17116
rect 13964 17076 13970 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14360 17116 14372 17125
rect 14327 17088 14372 17116
rect 14093 17079 14151 17085
rect 14360 17079 14372 17088
rect 14366 17076 14372 17079
rect 14424 17076 14430 17128
rect 10220 17051 10278 17057
rect 10220 17048 10232 17051
rect 6972 17020 8984 17048
rect 10060 17020 10232 17048
rect 6972 17008 6978 17020
rect 4246 16980 4252 16992
rect 2823 16952 4108 16980
rect 4207 16952 4252 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 4433 16983 4491 16989
rect 4433 16949 4445 16983
rect 4479 16980 4491 16983
rect 5902 16980 5908 16992
rect 4479 16952 5908 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 7561 16983 7619 16989
rect 7561 16980 7573 16983
rect 6052 16952 7573 16980
rect 6052 16940 6058 16952
rect 7561 16949 7573 16952
rect 7607 16949 7619 16983
rect 7561 16943 7619 16949
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 7929 16983 7987 16989
rect 7929 16980 7941 16983
rect 7708 16952 7941 16980
rect 7708 16940 7714 16952
rect 7929 16949 7941 16952
rect 7975 16949 7987 16983
rect 7929 16943 7987 16949
rect 8021 16983 8079 16989
rect 8021 16949 8033 16983
rect 8067 16980 8079 16983
rect 8846 16980 8852 16992
rect 8067 16952 8852 16980
rect 8067 16949 8079 16952
rect 8021 16943 8079 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 8956 16989 8984 17020
rect 10220 17017 10232 17020
rect 10266 17048 10278 17051
rect 11054 17048 11060 17060
rect 10266 17020 11060 17048
rect 10266 17017 10278 17020
rect 10220 17011 10278 17017
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 12342 17008 12348 17060
rect 12400 17048 12406 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12400 17020 12817 17048
rect 12400 17008 12406 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 17954 17048 17960 17060
rect 13780 17020 17960 17048
rect 13780 17008 13786 17020
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 8941 16983 8999 16989
rect 8941 16949 8953 16983
rect 8987 16949 8999 16983
rect 9306 16980 9312 16992
rect 9267 16952 9312 16980
rect 8941 16943 8999 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16980 9459 16983
rect 10502 16980 10508 16992
rect 9447 16952 10508 16980
rect 9447 16949 9459 16952
rect 9401 16943 9459 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11698 16980 11704 16992
rect 11655 16952 11704 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 15473 16983 15531 16989
rect 15473 16949 15485 16983
rect 15519 16980 15531 16983
rect 15838 16980 15844 16992
rect 15519 16952 15844 16980
rect 15519 16949 15531 16952
rect 15473 16943 15531 16949
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1486 16736 1492 16788
rect 1544 16776 1550 16788
rect 1673 16779 1731 16785
rect 1673 16776 1685 16779
rect 1544 16748 1685 16776
rect 1544 16736 1550 16748
rect 1673 16745 1685 16748
rect 1719 16745 1731 16779
rect 1673 16739 1731 16745
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 2958 16776 2964 16788
rect 2556 16748 2964 16776
rect 2556 16736 2562 16748
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3160 16748 4476 16776
rect 1762 16668 1768 16720
rect 1820 16708 1826 16720
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 1820 16680 2329 16708
rect 1820 16668 1826 16680
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16609 1547 16643
rect 1489 16603 1547 16609
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 3160 16640 3188 16748
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 3878 16708 3884 16720
rect 3292 16680 3884 16708
rect 3292 16668 3298 16680
rect 3878 16668 3884 16680
rect 3936 16668 3942 16720
rect 4246 16668 4252 16720
rect 4304 16717 4310 16720
rect 4304 16711 4368 16717
rect 4304 16677 4322 16711
rect 4356 16677 4368 16711
rect 4448 16708 4476 16748
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 4764 16748 5457 16776
rect 4764 16736 4770 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 5445 16739 5503 16745
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 7285 16779 7343 16785
rect 7285 16776 7297 16779
rect 5960 16748 7297 16776
rect 5960 16736 5966 16748
rect 7285 16745 7297 16748
rect 7331 16745 7343 16779
rect 7285 16739 7343 16745
rect 7561 16779 7619 16785
rect 7561 16745 7573 16779
rect 7607 16776 7619 16779
rect 7650 16776 7656 16788
rect 7607 16748 7656 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 5994 16708 6000 16720
rect 4448 16680 6000 16708
rect 4304 16671 4368 16677
rect 4304 16668 4310 16671
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6178 16717 6184 16720
rect 6172 16708 6184 16717
rect 6139 16680 6184 16708
rect 6172 16671 6184 16680
rect 6178 16668 6184 16671
rect 6236 16668 6242 16720
rect 7300 16708 7328 16739
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 7800 16748 8033 16776
rect 7800 16736 7806 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 9306 16776 9312 16788
rect 8619 16748 9312 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9401 16779 9459 16785
rect 9401 16745 9413 16779
rect 9447 16776 9459 16779
rect 11054 16776 11060 16788
rect 9447 16748 9812 16776
rect 11015 16748 11060 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 8941 16711 8999 16717
rect 7300 16680 8616 16708
rect 3326 16640 3332 16652
rect 2087 16612 3188 16640
rect 3287 16612 3332 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 1504 16572 1532 16603
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 4706 16640 4712 16652
rect 3988 16612 4712 16640
rect 2130 16572 2136 16584
rect 1504 16544 2136 16572
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 3418 16572 3424 16584
rect 3379 16544 3424 16572
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3988 16572 4016 16612
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 7929 16643 7987 16649
rect 4948 16612 7880 16640
rect 4948 16600 4954 16612
rect 3651 16544 4016 16572
rect 4065 16575 4123 16581
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 5810 16572 5816 16584
rect 4065 16535 4123 16541
rect 5083 16544 5816 16572
rect 2866 16464 2872 16516
rect 2924 16504 2930 16516
rect 3970 16504 3976 16516
rect 2924 16476 3976 16504
rect 2924 16464 2930 16476
rect 3970 16464 3976 16476
rect 4028 16504 4034 16516
rect 4080 16504 4108 16535
rect 4028 16476 4108 16504
rect 4028 16464 4034 16476
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 2961 16439 3019 16445
rect 2961 16436 2973 16439
rect 2832 16408 2973 16436
rect 2832 16396 2838 16408
rect 2961 16405 2973 16408
rect 3007 16405 3019 16439
rect 4080 16436 4108 16476
rect 5083 16436 5111 16544
rect 5810 16532 5816 16544
rect 5868 16572 5874 16584
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 5868 16544 5917 16572
rect 5868 16532 5874 16544
rect 5905 16541 5917 16544
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 7852 16504 7880 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8478 16640 8484 16652
rect 7975 16612 8484 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8588 16640 8616 16680
rect 8941 16677 8953 16711
rect 8987 16708 8999 16711
rect 9674 16708 9680 16720
rect 8987 16680 9680 16708
rect 8987 16677 8999 16680
rect 8941 16671 8999 16677
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 9784 16708 9812 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 11204 16748 11345 16776
rect 11204 16736 11210 16748
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 11790 16776 11796 16788
rect 11751 16748 11796 16776
rect 11333 16739 11391 16745
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 12989 16779 13047 16785
rect 12989 16745 13001 16779
rect 13035 16776 13047 16779
rect 13035 16748 14136 16776
rect 13035 16745 13047 16748
rect 12989 16739 13047 16745
rect 13722 16708 13728 16720
rect 9784 16680 13728 16708
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 9401 16643 9459 16649
rect 9401 16640 9413 16643
rect 8588 16612 9413 16640
rect 9401 16609 9413 16612
rect 9447 16609 9459 16643
rect 9944 16643 10002 16649
rect 9944 16640 9956 16643
rect 9401 16603 9459 16609
rect 9600 16612 9956 16640
rect 8202 16572 8208 16584
rect 8163 16544 8208 16572
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9033 16575 9091 16581
rect 9033 16572 9045 16575
rect 8312 16544 9045 16572
rect 8312 16504 8340 16544
rect 9033 16541 9045 16544
rect 9079 16541 9091 16575
rect 9033 16535 9091 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16572 9275 16575
rect 9600 16572 9628 16612
rect 9944 16609 9956 16612
rect 9990 16640 10002 16643
rect 10226 16640 10232 16652
rect 9990 16612 10232 16640
rect 9990 16609 10002 16612
rect 9944 16603 10002 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 11698 16640 11704 16652
rect 11659 16612 11704 16640
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 13348 16643 13406 16649
rect 13348 16609 13360 16643
rect 13394 16640 13406 16643
rect 13814 16640 13820 16652
rect 13394 16612 13820 16640
rect 13394 16609 13406 16612
rect 13348 16603 13406 16609
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 9263 16544 9628 16572
rect 9677 16575 9735 16581
rect 9263 16541 9275 16544
rect 9217 16535 9275 16541
rect 9677 16541 9689 16575
rect 9723 16541 9735 16575
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 9677 16535 9735 16541
rect 7852 16476 8340 16504
rect 8754 16464 8760 16516
rect 8812 16504 8818 16516
rect 9490 16504 9496 16516
rect 8812 16476 9496 16504
rect 8812 16464 8818 16476
rect 9490 16464 9496 16476
rect 9548 16504 9554 16516
rect 9692 16504 9720 16535
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 14108 16572 14136 16748
rect 14366 16736 14372 16788
rect 14424 16776 14430 16788
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 14424 16748 14473 16776
rect 14424 16736 14430 16748
rect 14461 16745 14473 16748
rect 14507 16745 14519 16779
rect 14461 16739 14519 16745
rect 15562 16572 15568 16584
rect 14108 16544 15568 16572
rect 13081 16535 13139 16541
rect 11698 16504 11704 16516
rect 9548 16476 9720 16504
rect 10980 16476 11704 16504
rect 9548 16464 9554 16476
rect 4080 16408 5111 16436
rect 2961 16399 3019 16405
rect 5258 16396 5264 16448
rect 5316 16436 5322 16448
rect 10980 16436 11008 16476
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 5316 16408 11008 16436
rect 5316 16396 5322 16408
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 11112 16408 13001 16436
rect 11112 16396 11118 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 13096 16436 13124 16535
rect 15562 16532 15568 16544
rect 15620 16532 15626 16584
rect 13722 16436 13728 16448
rect 13096 16408 13728 16436
rect 12989 16399 13047 16405
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 20346 16436 20352 16448
rect 17460 16408 20352 16436
rect 17460 16396 17466 16408
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1673 16235 1731 16241
rect 1673 16232 1685 16235
rect 1636 16204 1685 16232
rect 1636 16192 1642 16204
rect 1673 16201 1685 16204
rect 1719 16201 1731 16235
rect 1673 16195 1731 16201
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3973 16235 4031 16241
rect 3973 16232 3985 16235
rect 3476 16204 3985 16232
rect 3476 16192 3482 16204
rect 3973 16201 3985 16204
rect 4019 16201 4031 16235
rect 6914 16232 6920 16244
rect 3973 16195 4031 16201
rect 5184 16204 6920 16232
rect 5184 16164 5212 16204
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 8570 16232 8576 16244
rect 8531 16204 8576 16232
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 10502 16232 10508 16244
rect 10463 16204 10508 16232
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 14332 16204 15117 16232
rect 14332 16192 14338 16204
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 16114 16232 16120 16244
rect 16075 16204 16120 16232
rect 15105 16195 15163 16201
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 2056 16136 5212 16164
rect 5261 16167 5319 16173
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 2056 16037 2084 16136
rect 5261 16133 5273 16167
rect 5307 16164 5319 16167
rect 5718 16164 5724 16176
rect 5307 16136 5724 16164
rect 5307 16133 5319 16136
rect 5261 16127 5319 16133
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 2188 16068 2237 16096
rect 2188 16056 2194 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3142 16096 3148 16108
rect 3099 16068 3148 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 3326 16056 3332 16108
rect 3384 16096 3390 16108
rect 3513 16099 3571 16105
rect 3513 16096 3525 16099
rect 3384 16068 3525 16096
rect 3384 16056 3390 16068
rect 3513 16065 3525 16068
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 4304 16068 4537 16096
rect 4304 16056 4310 16068
rect 4525 16065 4537 16068
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 5534 16056 5540 16108
rect 5592 16096 5598 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5592 16068 5825 16096
rect 5592 16056 5598 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 8588 16096 8616 16192
rect 10226 16164 10232 16176
rect 10139 16136 10232 16164
rect 10226 16124 10232 16136
rect 10284 16124 10290 16176
rect 13832 16164 13860 16192
rect 13832 16136 15700 16164
rect 10244 16096 10272 16124
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 8588 16068 8984 16096
rect 10244 16068 11069 16096
rect 5813 16059 5871 16065
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 4433 16031 4491 16037
rect 2832 16000 2877 16028
rect 2832 15988 2838 16000
rect 4433 15997 4445 16031
rect 4479 16028 4491 16031
rect 5166 16028 5172 16040
rect 4479 16000 5172 16028
rect 4479 15997 4491 16000
rect 4433 15991 4491 15997
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 16028 7251 16031
rect 8294 16028 8300 16040
rect 7239 16000 8300 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 8294 15988 8300 16000
rect 8352 16028 8358 16040
rect 8754 16028 8760 16040
rect 8352 16000 8760 16028
rect 8352 15988 8358 16000
rect 8754 15988 8760 16000
rect 8812 16028 8818 16040
rect 8849 16031 8907 16037
rect 8849 16028 8861 16031
rect 8812 16000 8861 16028
rect 8812 15988 8818 16000
rect 8849 15997 8861 16000
rect 8895 15997 8907 16031
rect 8956 16028 8984 16068
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 11057 16059 11115 16065
rect 13740 16068 14657 16096
rect 9105 16031 9163 16037
rect 9105 16028 9117 16031
rect 8956 16000 9117 16028
rect 8849 15991 8907 15997
rect 9105 15997 9117 16000
rect 9151 15997 9163 16031
rect 9105 15991 9163 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12704 16031 12762 16037
rect 12704 15997 12716 16031
rect 12750 16028 12762 16031
rect 12986 16028 12992 16040
rect 12750 16000 12992 16028
rect 12750 15997 12762 16000
rect 12704 15991 12762 15997
rect 4341 15963 4399 15969
rect 4341 15929 4353 15963
rect 4387 15960 4399 15963
rect 4890 15960 4896 15972
rect 4387 15932 4896 15960
rect 4387 15929 4399 15932
rect 4341 15923 4399 15929
rect 4890 15920 4896 15932
rect 4948 15920 4954 15972
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 5350 15960 5356 15972
rect 5040 15932 5356 15960
rect 5040 15920 5046 15932
rect 5350 15920 5356 15932
rect 5408 15960 5414 15972
rect 5721 15963 5779 15969
rect 5721 15960 5733 15963
rect 5408 15932 5733 15960
rect 5408 15920 5414 15932
rect 5721 15929 5733 15932
rect 5767 15929 5779 15963
rect 5721 15923 5779 15929
rect 7460 15963 7518 15969
rect 7460 15929 7472 15963
rect 7506 15960 7518 15963
rect 8202 15960 8208 15972
rect 7506 15932 8208 15960
rect 7506 15929 7518 15932
rect 7460 15923 7518 15929
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 10870 15960 10876 15972
rect 10831 15932 10876 15960
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 12452 15960 12480 15991
rect 12986 15988 12992 16000
rect 13044 16028 13050 16040
rect 13740 16028 13768 16068
rect 14645 16065 14657 16068
rect 14691 16096 14703 16099
rect 15194 16096 15200 16108
rect 14691 16068 15200 16096
rect 14691 16065 14703 16068
rect 14645 16059 14703 16065
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15672 16105 15700 16136
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 15703 16068 16681 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 13044 16000 13768 16028
rect 13044 15988 13050 16000
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 13872 16000 14565 16028
rect 13872 15988 13878 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15160 16000 15485 16028
rect 15160 15988 15166 16000
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 13906 15960 13912 15972
rect 12452 15932 13912 15960
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 15565 15963 15623 15969
rect 15565 15960 15577 15963
rect 14108 15932 15577 15960
rect 4908 15892 4936 15920
rect 5258 15892 5264 15904
rect 4908 15864 5264 15892
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 5626 15892 5632 15904
rect 5587 15864 5632 15892
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 10965 15895 11023 15901
rect 10965 15861 10977 15895
rect 11011 15892 11023 15895
rect 11054 15892 11060 15904
rect 11011 15864 11060 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 14108 15901 14136 15932
rect 15565 15929 15577 15932
rect 15611 15929 15623 15963
rect 15565 15923 15623 15929
rect 15654 15920 15660 15972
rect 15712 15960 15718 15972
rect 16577 15963 16635 15969
rect 16577 15960 16589 15963
rect 15712 15932 16589 15960
rect 15712 15920 15718 15932
rect 16577 15929 16589 15932
rect 16623 15929 16635 15963
rect 16577 15923 16635 15929
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15861 14151 15895
rect 14458 15892 14464 15904
rect 14419 15864 14464 15892
rect 14093 15855 14151 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 16482 15892 16488 15904
rect 16443 15864 16488 15892
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1728 15660 1777 15688
rect 1728 15648 1734 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 3050 15688 3056 15700
rect 3011 15660 3056 15688
rect 1765 15651 1823 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 8478 15688 8484 15700
rect 8439 15660 8484 15688
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8904 15660 9689 15688
rect 8904 15648 8910 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 10134 15688 10140 15700
rect 10095 15660 10140 15688
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 11241 15691 11299 15697
rect 11241 15657 11253 15691
rect 11287 15657 11299 15691
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 11241 15651 11299 15657
rect 1486 15580 1492 15632
rect 1544 15620 1550 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 1544 15592 2421 15620
rect 1544 15580 1550 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 5436 15623 5494 15629
rect 5436 15589 5448 15623
rect 5482 15620 5494 15623
rect 5534 15620 5540 15632
rect 5482 15592 5540 15620
rect 5482 15589 5494 15592
rect 5436 15583 5494 15589
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 9876 15620 9904 15648
rect 11256 15620 11284 15651
rect 11698 15648 11704 15660
rect 11756 15688 11762 15700
rect 11882 15688 11888 15700
rect 11756 15660 11888 15688
rect 11756 15648 11762 15660
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15688 12311 15691
rect 12894 15688 12900 15700
rect 12299 15660 12900 15688
rect 12299 15657 12311 15660
rect 12253 15651 12311 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14366 15688 14372 15700
rect 14148 15660 14372 15688
rect 14148 15648 14154 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 14921 15691 14979 15697
rect 14921 15657 14933 15691
rect 14967 15688 14979 15691
rect 15194 15688 15200 15700
rect 14967 15660 15200 15688
rect 14967 15657 14979 15660
rect 14921 15651 14979 15657
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15688 15347 15691
rect 16482 15688 16488 15700
rect 15335 15660 16488 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 14458 15620 14464 15632
rect 9876 15592 10180 15620
rect 11256 15592 14464 15620
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 1854 15552 1860 15564
rect 1627 15524 1860 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2122 15555 2180 15561
rect 2122 15521 2134 15555
rect 2168 15521 2180 15555
rect 2122 15515 2180 15521
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 3050 15552 3056 15564
rect 2915 15524 3056 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 2139 15416 2167 15515
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 5169 15555 5227 15561
rect 5169 15552 5181 15555
rect 4028 15524 5181 15552
rect 4028 15512 4034 15524
rect 5169 15521 5181 15524
rect 5215 15521 5227 15555
rect 7081 15555 7139 15561
rect 7081 15552 7093 15555
rect 5169 15515 5227 15521
rect 6564 15524 7093 15552
rect 4706 15416 4712 15428
rect 2139 15388 4712 15416
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 6454 15308 6460 15360
rect 6512 15348 6518 15360
rect 6564 15357 6592 15524
rect 7081 15521 7093 15524
rect 7127 15521 7139 15555
rect 7081 15515 7139 15521
rect 9858 15512 9864 15564
rect 9916 15552 9922 15564
rect 10042 15552 10048 15564
rect 9916 15524 10048 15552
rect 9916 15512 9922 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10152 15552 10180 15592
rect 14458 15580 14464 15592
rect 14516 15580 14522 15632
rect 15212 15620 15240 15648
rect 15212 15592 15792 15620
rect 10686 15552 10692 15564
rect 10152 15524 10692 15552
rect 10686 15512 10692 15524
rect 10744 15552 10750 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 10744 15524 11621 15552
rect 10744 15512 10750 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 12066 15552 12072 15564
rect 11848 15524 12072 15552
rect 11848 15512 11854 15524
rect 12066 15512 12072 15524
rect 12124 15552 12130 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12124 15524 12633 15552
rect 12124 15512 12130 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 13630 15512 13636 15564
rect 13688 15552 13694 15564
rect 13797 15555 13855 15561
rect 13797 15552 13809 15555
rect 13688 15524 13809 15552
rect 13688 15512 13694 15524
rect 13797 15521 13809 15524
rect 13843 15521 13855 15555
rect 13797 15515 13855 15521
rect 14090 15512 14096 15564
rect 14148 15552 14154 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 14148 15524 15669 15552
rect 14148 15512 14154 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15764 15552 15792 15592
rect 15764 15524 15884 15552
rect 15657 15515 15715 15521
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 6512 15320 6561 15348
rect 6512 15308 6518 15320
rect 6549 15317 6561 15320
rect 6595 15317 6607 15351
rect 6840 15348 6868 15447
rect 8202 15416 8208 15428
rect 8115 15388 8208 15416
rect 8202 15376 8208 15388
rect 8260 15416 8266 15428
rect 10244 15416 10272 15447
rect 8260 15388 10272 15416
rect 11900 15416 11928 15447
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 12308 15456 12725 15484
rect 12308 15444 12314 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 12713 15447 12771 15453
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15484 12955 15487
rect 12986 15484 12992 15496
rect 12943 15456 12992 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 12912 15416 12940 15447
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15453 13599 15487
rect 15746 15484 15752 15496
rect 15707 15456 15752 15484
rect 13541 15447 13599 15453
rect 11900 15388 12940 15416
rect 8260 15376 8266 15388
rect 8294 15348 8300 15360
rect 6840 15320 8300 15348
rect 6549 15311 6607 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 12066 15348 12072 15360
rect 10192 15320 12072 15348
rect 10192 15308 10198 15320
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 13556 15348 13584 15447
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 15856 15493 15884 15524
rect 15841 15487 15899 15493
rect 15841 15453 15853 15487
rect 15887 15484 15899 15487
rect 15930 15484 15936 15496
rect 15887 15456 15936 15484
rect 15887 15453 15899 15456
rect 15841 15447 15899 15453
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 13906 15348 13912 15360
rect 13556 15320 13912 15348
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 12437 15147 12495 15153
rect 1872 15116 5111 15144
rect 566 15036 572 15088
rect 624 15076 630 15088
rect 1872 15076 1900 15116
rect 624 15048 1900 15076
rect 5083 15076 5111 15116
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 13814 15144 13820 15156
rect 12483 15116 13820 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 15197 15147 15255 15153
rect 15197 15113 15209 15147
rect 15243 15144 15255 15147
rect 15654 15144 15660 15156
rect 15243 15116 15660 15144
rect 15243 15113 15255 15116
rect 15197 15107 15255 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 12802 15076 12808 15088
rect 5083 15048 12808 15076
rect 624 15036 630 15048
rect 12802 15036 12808 15048
rect 12860 15036 12866 15088
rect 13630 15076 13636 15088
rect 13096 15048 13636 15076
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 2317 15011 2375 15017
rect 2317 15008 2329 15011
rect 1912 14980 2329 15008
rect 1912 14968 1918 14980
rect 2317 14977 2329 14980
rect 2363 14977 2375 15011
rect 3050 15008 3056 15020
rect 3011 14980 3056 15008
rect 2317 14971 2375 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5684 14980 5825 15008
rect 5684 14968 5690 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 9398 15008 9404 15020
rect 8067 14980 9404 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 1578 14940 1584 14952
rect 1539 14912 1584 14940
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14909 2191 14943
rect 2133 14903 2191 14909
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 2958 14940 2964 14952
rect 2915 14912 2964 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 2148 14804 2176 14903
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 4028 14912 4169 14940
rect 4028 14900 4034 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 5534 14940 5540 14952
rect 5447 14912 5540 14940
rect 4157 14903 4215 14909
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 7484 14940 7512 14971
rect 9398 14968 9404 14980
rect 9456 14968 9462 15020
rect 9674 15008 9680 15020
rect 9635 14980 9680 15008
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 10962 15008 10968 15020
rect 10923 14980 10968 15008
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13096 15017 13124 15048
rect 13630 15036 13636 15048
rect 13688 15076 13694 15088
rect 13688 15048 14596 15076
rect 13688 15036 13694 15048
rect 14568 15020 14596 15048
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 13044 14980 13093 15008
rect 13044 14968 13050 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 14090 15008 14096 15020
rect 13771 14980 14096 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 14608 14980 14749 15008
rect 14608 14968 14614 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 15930 15008 15936 15020
rect 15887 14980 15936 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 5592 14912 7512 14940
rect 5592 14900 5598 14912
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 8260 14912 8309 14940
rect 8260 14900 8266 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 8938 14900 8944 14952
rect 8996 14940 9002 14952
rect 11606 14940 11612 14952
rect 8996 14912 11612 14940
rect 8996 14900 9002 14912
rect 11606 14900 11612 14912
rect 11664 14940 11670 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 11664 14912 12909 14940
rect 11664 14900 11670 14912
rect 12897 14909 12909 14912
rect 12943 14940 12955 14943
rect 15378 14940 15384 14952
rect 12943 14912 15384 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 4424 14875 4482 14881
rect 4424 14841 4436 14875
rect 4470 14872 4482 14875
rect 5442 14872 5448 14884
rect 4470 14844 5448 14872
rect 4470 14841 4482 14844
rect 4424 14835 4482 14841
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 5074 14804 5080 14816
rect 2148 14776 5080 14804
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5552 14813 5580 14900
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 10134 14872 10140 14884
rect 7239 14844 10140 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 10781 14875 10839 14881
rect 10781 14841 10793 14875
rect 10827 14872 10839 14875
rect 12250 14872 12256 14884
rect 10827 14844 12256 14872
rect 10827 14841 10839 14844
rect 10781 14835 10839 14841
rect 12250 14832 12256 14844
rect 12308 14832 12314 14884
rect 12802 14872 12808 14884
rect 12763 14844 12808 14872
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 15657 14875 15715 14881
rect 15657 14872 15669 14875
rect 14200 14844 15669 14872
rect 5537 14807 5595 14813
rect 5537 14773 5549 14807
rect 5583 14773 5595 14807
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 5537 14767 5595 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7331 14776 8033 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 8021 14773 8033 14776
rect 8067 14773 8079 14807
rect 8021 14767 8079 14773
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 8294 14804 8300 14816
rect 8159 14776 8300 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 8294 14764 8300 14776
rect 8352 14804 8358 14816
rect 8662 14804 8668 14816
rect 8352 14776 8668 14804
rect 8352 14764 8358 14776
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 10410 14804 10416 14816
rect 10371 14776 10416 14804
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10873 14807 10931 14813
rect 10873 14773 10885 14807
rect 10919 14804 10931 14807
rect 11146 14804 11152 14816
rect 10919 14776 11152 14804
rect 10919 14773 10931 14776
rect 10873 14767 10931 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 14200 14813 14228 14844
rect 15657 14841 15669 14844
rect 15703 14841 15715 14875
rect 15657 14835 15715 14841
rect 14185 14807 14243 14813
rect 14185 14773 14197 14807
rect 14231 14773 14243 14807
rect 14185 14767 14243 14773
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 14332 14776 14565 14804
rect 14332 14764 14338 14776
rect 14553 14773 14565 14776
rect 14599 14773 14611 14807
rect 14553 14767 14611 14773
rect 14645 14807 14703 14813
rect 14645 14773 14657 14807
rect 14691 14804 14703 14807
rect 15286 14804 15292 14816
rect 14691 14776 15292 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15562 14804 15568 14816
rect 15523 14776 15568 14804
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 1857 14603 1915 14609
rect 1857 14600 1869 14603
rect 1728 14572 1869 14600
rect 1728 14560 1734 14572
rect 1857 14569 1869 14572
rect 1903 14569 1915 14603
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 1857 14563 1915 14569
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 4890 14600 4896 14612
rect 3712 14572 4896 14600
rect 3712 14532 3740 14572
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5442 14600 5448 14612
rect 5403 14572 5448 14600
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 8294 14600 8300 14612
rect 6012 14572 8300 14600
rect 5460 14532 5488 14560
rect 2240 14504 3740 14532
rect 3988 14504 5488 14532
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 1854 14464 1860 14476
rect 1719 14436 1860 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 2240 14473 2268 14504
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14433 2283 14467
rect 3326 14464 3332 14476
rect 3287 14436 3332 14464
rect 2225 14427 2283 14433
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 1578 14356 1584 14408
rect 1636 14396 1642 14408
rect 2409 14399 2467 14405
rect 2409 14396 2421 14399
rect 1636 14368 2421 14396
rect 1636 14356 1642 14368
rect 2409 14365 2421 14368
rect 2455 14365 2467 14399
rect 2409 14359 2467 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14396 3663 14399
rect 3988 14396 4016 14504
rect 4332 14467 4390 14473
rect 4332 14433 4344 14467
rect 4378 14464 4390 14467
rect 5902 14464 5908 14476
rect 4378 14436 5908 14464
rect 4378 14433 4390 14436
rect 4332 14427 4390 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6012 14473 6040 14572
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 10008 14572 10149 14600
rect 10008 14560 10014 14572
rect 10137 14569 10149 14572
rect 10183 14600 10195 14603
rect 11054 14600 11060 14612
rect 10183 14572 11060 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 12342 14600 12348 14612
rect 12303 14572 12348 14600
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12676 14572 12725 14600
rect 12676 14560 12682 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 14001 14603 14059 14609
rect 14001 14569 14013 14603
rect 14047 14600 14059 14603
rect 15562 14600 15568 14612
rect 14047 14572 15568 14600
rect 14047 14569 14059 14572
rect 14001 14563 14059 14569
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 6641 14535 6699 14541
rect 6641 14501 6653 14535
rect 6687 14532 6699 14535
rect 7650 14532 7656 14544
rect 6687 14504 7656 14532
rect 6687 14501 6699 14504
rect 6641 14495 6699 14501
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 8196 14535 8254 14541
rect 8196 14501 8208 14535
rect 8242 14532 8254 14535
rect 8478 14532 8484 14544
rect 8242 14504 8484 14532
rect 8242 14501 8254 14504
rect 8196 14495 8254 14501
rect 8478 14492 8484 14504
rect 8536 14532 8542 14544
rect 8536 14504 10272 14532
rect 8536 14492 8542 14504
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 6914 14464 6920 14476
rect 6779 14436 6920 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8662 14464 8668 14476
rect 7975 14436 8668 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8662 14424 8668 14436
rect 8720 14424 8726 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 3651 14368 4016 14396
rect 4065 14399 4123 14405
rect 3651 14365 3663 14368
rect 3605 14359 3663 14365
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 6825 14399 6883 14405
rect 6825 14365 6837 14399
rect 6871 14396 6883 14399
rect 7098 14396 7104 14408
rect 6871 14368 7104 14396
rect 6871 14365 6883 14368
rect 6825 14359 6883 14365
rect 3436 14260 3464 14359
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4080 14328 4108 14359
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 10244 14405 10272 14504
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 10778 14532 10784 14544
rect 10652 14504 10784 14532
rect 10652 14492 10658 14504
rect 10778 14492 10784 14504
rect 10836 14532 10842 14544
rect 11701 14535 11759 14541
rect 11701 14532 11713 14535
rect 10836 14504 11713 14532
rect 10836 14492 10842 14504
rect 11701 14501 11713 14504
rect 11747 14501 11759 14535
rect 11701 14495 11759 14501
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 12158 14532 12164 14544
rect 11839 14504 12164 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 11716 14464 11744 14495
rect 12158 14492 12164 14504
rect 12216 14532 12222 14544
rect 15657 14535 15715 14541
rect 15657 14532 15669 14535
rect 12216 14504 15669 14532
rect 12216 14492 12222 14504
rect 15657 14501 15669 14504
rect 15703 14501 15715 14535
rect 15657 14495 15715 14501
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 11716 14436 12817 14464
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 14366 14464 14372 14476
rect 14327 14436 14372 14464
rect 12805 14427 12863 14433
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 14507 14436 15240 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12158 14396 12164 14408
rect 12023 14368 12164 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12986 14396 12992 14408
rect 12947 14368 12992 14396
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 14476 14396 14504 14427
rect 13136 14368 14504 14396
rect 13136 14356 13142 14368
rect 14550 14356 14556 14408
rect 14608 14396 14614 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14608 14368 14657 14396
rect 14608 14356 14614 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 4028 14300 4108 14328
rect 4028 14288 4034 14300
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 6273 14331 6331 14337
rect 6273 14328 6285 14331
rect 5132 14300 6285 14328
rect 5132 14288 5138 14300
rect 6273 14297 6285 14300
rect 6319 14297 6331 14331
rect 6273 14291 6331 14297
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 10870 14328 10876 14340
rect 9355 14300 10876 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 5626 14260 5632 14272
rect 3436 14232 5632 14260
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 5810 14260 5816 14272
rect 5771 14232 5816 14260
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 9324 14260 9352 14291
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 14660 14328 14688 14359
rect 15102 14328 15108 14340
rect 14660 14300 15108 14328
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15212 14328 15240 14436
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15749 14467 15807 14473
rect 15749 14464 15761 14467
rect 15436 14436 15761 14464
rect 15436 14424 15442 14436
rect 15749 14433 15761 14436
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 15896 14368 15941 14396
rect 15896 14356 15902 14368
rect 18966 14328 18972 14340
rect 15212 14300 18972 14328
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 5960 14232 9352 14260
rect 9677 14263 9735 14269
rect 5960 14220 5966 14232
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 10778 14260 10784 14272
rect 9723 14232 10784 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11333 14263 11391 14269
rect 11333 14229 11345 14263
rect 11379 14260 11391 14263
rect 11698 14260 11704 14272
rect 11379 14232 11704 14260
rect 11379 14229 11391 14232
rect 11333 14223 11391 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 15286 14260 15292 14272
rect 15247 14232 15292 14260
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 2832 14028 2877 14056
rect 2832 14016 2838 14028
rect 3326 14016 3332 14068
rect 3384 14056 3390 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 3384 14028 4077 14056
rect 3384 14016 3390 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 4065 14019 4123 14025
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 4764 14028 5365 14056
rect 4764 14016 4770 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 5353 14019 5411 14025
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 8389 14059 8447 14065
rect 5684 14028 7972 14056
rect 5684 14016 5690 14028
rect 4246 13988 4252 14000
rect 1872 13960 4252 13988
rect 1872 13861 1900 13960
rect 4246 13948 4252 13960
rect 4304 13948 4310 14000
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 4890 13988 4896 14000
rect 4672 13960 4896 13988
rect 4672 13948 4678 13960
rect 4890 13948 4896 13960
rect 4948 13948 4954 14000
rect 7944 13988 7972 14028
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 8478 14056 8484 14068
rect 8435 14028 8484 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 10008 14028 10057 14056
rect 10008 14016 10014 14028
rect 10045 14025 10057 14028
rect 10091 14056 10103 14059
rect 10962 14056 10968 14068
rect 10091 14028 10968 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 15194 14056 15200 14068
rect 11072 14028 15200 14056
rect 7944 13960 8064 13988
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 5902 13920 5908 13932
rect 4755 13892 5908 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 5902 13880 5908 13892
rect 5960 13880 5966 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6454 13920 6460 13932
rect 6043 13892 6460 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 8036 13920 8064 13960
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 11072 13988 11100 14028
rect 15194 14016 15200 14028
rect 15252 14056 15258 14068
rect 18598 14056 18604 14068
rect 15252 14028 18604 14056
rect 15252 14016 15258 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 10192 13960 11100 13988
rect 10192 13948 10198 13960
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 11664 13960 11836 13988
rect 11664 13948 11670 13960
rect 10870 13920 10876 13932
rect 8036 13892 8800 13920
rect 10831 13892 10876 13920
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2096 13824 2605 13852
rect 2096 13812 2102 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 3133 13855 3191 13861
rect 3133 13821 3145 13855
rect 3179 13821 3191 13855
rect 3133 13815 3191 13821
rect 2133 13787 2191 13793
rect 2133 13753 2145 13787
rect 2179 13784 2191 13787
rect 3151 13784 3179 13815
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 4525 13855 4583 13861
rect 3292 13824 3372 13852
rect 3292 13812 3298 13824
rect 2179 13756 3179 13784
rect 2179 13753 2191 13756
rect 2133 13747 2191 13753
rect 3344 13725 3372 13824
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4798 13852 4804 13864
rect 4571 13824 4804 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6822 13852 6828 13864
rect 5859 13824 6828 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 5718 13784 5724 13796
rect 5679 13756 5724 13784
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 7024 13784 7052 13815
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7265 13855 7323 13861
rect 7265 13852 7277 13855
rect 7156 13824 7277 13852
rect 7156 13812 7162 13824
rect 7265 13821 7277 13824
rect 7311 13821 7323 13855
rect 8662 13852 8668 13864
rect 7265 13815 7323 13821
rect 7392 13824 8668 13852
rect 7392 13784 7420 13824
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 8772 13852 8800 13892
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11808 13861 11836 13960
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12621 13991 12679 13997
rect 12621 13988 12633 13991
rect 12492 13960 12633 13988
rect 12492 13948 12498 13960
rect 12621 13957 12633 13960
rect 12667 13957 12679 13991
rect 13170 13988 13176 14000
rect 13131 13960 13176 13988
rect 12621 13951 12679 13957
rect 13170 13948 13176 13960
rect 13228 13948 13234 14000
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 14185 13991 14243 13997
rect 14185 13988 14197 13991
rect 13964 13960 14197 13988
rect 13964 13948 13970 13960
rect 14185 13957 14197 13960
rect 14231 13988 14243 13991
rect 14274 13988 14280 14000
rect 14231 13960 14280 13988
rect 14231 13957 14243 13960
rect 14185 13951 14243 13957
rect 14274 13948 14280 13960
rect 14332 13988 14338 14000
rect 14332 13960 15056 13988
rect 14332 13948 14338 13960
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12158 13920 12164 13932
rect 12023 13892 12164 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12158 13880 12164 13892
rect 12216 13920 12222 13932
rect 15028 13929 15056 13960
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 12216 13892 13737 13920
rect 12216 13880 12222 13892
rect 13725 13889 13737 13892
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 11793 13855 11851 13861
rect 8772 13824 10364 13852
rect 7024 13756 7420 13784
rect 3329 13719 3387 13725
rect 3329 13685 3341 13719
rect 3375 13685 3387 13719
rect 4430 13716 4436 13728
rect 4391 13688 4436 13716
rect 3329 13679 3387 13685
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 8680 13716 8708 13812
rect 8932 13787 8990 13793
rect 8932 13753 8944 13787
rect 8978 13784 8990 13787
rect 9122 13784 9128 13796
rect 8978 13756 9128 13784
rect 8978 13753 8990 13756
rect 8932 13747 8990 13753
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 9582 13716 9588 13728
rect 8680 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10226 13716 10232 13728
rect 9824 13688 10232 13716
rect 9824 13676 9830 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10336 13725 10364 13824
rect 11793 13821 11805 13855
rect 11839 13821 11851 13855
rect 12802 13852 12808 13864
rect 12715 13824 12808 13852
rect 11793 13815 11851 13821
rect 12802 13812 12808 13824
rect 12860 13852 12866 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 12860 13824 14381 13852
rect 12860 13812 12866 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 15280 13855 15338 13861
rect 15280 13821 15292 13855
rect 15326 13852 15338 13855
rect 15838 13852 15844 13864
rect 15326 13824 15844 13852
rect 15326 13821 15338 13824
rect 15280 13815 15338 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 10689 13787 10747 13793
rect 10689 13753 10701 13787
rect 10735 13784 10747 13787
rect 13354 13784 13360 13796
rect 10735 13756 13360 13784
rect 10735 13753 10747 13756
rect 10689 13747 10747 13753
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 13541 13787 13599 13793
rect 13541 13753 13553 13787
rect 13587 13784 13599 13787
rect 14182 13784 14188 13796
rect 13587 13756 14188 13784
rect 13587 13753 13599 13756
rect 13541 13747 13599 13753
rect 10321 13719 10379 13725
rect 10321 13685 10333 13719
rect 10367 13685 10379 13719
rect 10778 13716 10784 13728
rect 10739 13688 10784 13716
rect 10321 13679 10379 13685
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11422 13716 11428 13728
rect 11379 13688 11428 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 11882 13716 11888 13728
rect 11747 13688 11888 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 13556 13716 13584 13747
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 12584 13688 13584 13716
rect 13633 13719 13691 13725
rect 12584 13676 12590 13688
rect 13633 13685 13645 13719
rect 13679 13716 13691 13719
rect 15378 13716 15384 13728
rect 13679 13688 15384 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 16390 13716 16396 13728
rect 16351 13688 16396 13716
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 4430 13512 4436 13524
rect 4391 13484 4436 13512
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 7156 13484 7389 13512
rect 7156 13472 7162 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7650 13512 7656 13524
rect 7611 13484 7656 13512
rect 7377 13475 7435 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 11514 13512 11520 13524
rect 9180 13484 11520 13512
rect 9180 13472 9186 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 12308 13484 12357 13512
rect 12308 13472 12314 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12345 13475 12403 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12805 13515 12863 13521
rect 12492 13484 12756 13512
rect 12492 13472 12498 13484
rect 3421 13447 3479 13453
rect 3421 13413 3433 13447
rect 3467 13444 3479 13447
rect 3602 13444 3608 13456
rect 3467 13416 3608 13444
rect 3467 13413 3479 13416
rect 3421 13407 3479 13413
rect 3602 13404 3608 13416
rect 3660 13404 3666 13456
rect 3878 13404 3884 13456
rect 3936 13444 3942 13456
rect 3936 13416 10088 13444
rect 3936 13404 3942 13416
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 1946 13376 1952 13388
rect 1903 13348 1952 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 3326 13376 3332 13388
rect 3287 13348 3332 13376
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 6264 13379 6322 13385
rect 6264 13345 6276 13379
rect 6310 13376 6322 13379
rect 7098 13376 7104 13388
rect 6310 13348 7104 13376
rect 6310 13345 6322 13348
rect 6264 13339 6322 13345
rect 7098 13336 7104 13348
rect 7156 13376 7162 13388
rect 7466 13376 7472 13388
rect 7156 13348 7472 13376
rect 7156 13336 7162 13348
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 9950 13385 9956 13388
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8067 13348 8677 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 9944 13376 9956 13385
rect 9911 13348 9956 13376
rect 8665 13339 8723 13345
rect 9944 13339 9956 13348
rect 9950 13336 9956 13339
rect 10008 13336 10014 13388
rect 10060 13376 10088 13416
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 10594 13444 10600 13456
rect 10376 13416 10600 13444
rect 10376 13404 10382 13416
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 11422 13404 11428 13456
rect 11480 13444 11486 13456
rect 11793 13447 11851 13453
rect 11793 13444 11805 13447
rect 11480 13416 11805 13444
rect 11480 13404 11486 13416
rect 11793 13413 11805 13416
rect 11839 13413 11851 13447
rect 11793 13407 11851 13413
rect 12161 13447 12219 13453
rect 12161 13413 12173 13447
rect 12207 13444 12219 13447
rect 12526 13444 12532 13456
rect 12207 13416 12532 13444
rect 12207 13413 12219 13416
rect 12161 13407 12219 13413
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 12728 13444 12756 13484
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 13170 13512 13176 13524
rect 12851 13484 13176 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15344 13484 15761 13512
rect 15344 13472 15350 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 12728 13416 13492 13444
rect 12710 13376 12716 13388
rect 10060 13348 11376 13376
rect 12671 13348 12716 13376
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1452 13280 2053 13308
rect 1452 13268 1458 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2041 13271 2099 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 3694 13308 3700 13320
rect 3651 13280 3700 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 3694 13268 3700 13280
rect 3752 13308 3758 13320
rect 5534 13308 5540 13320
rect 3752 13280 5540 13308
rect 3752 13268 3758 13280
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5776 13280 6009 13308
rect 5776 13268 5782 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7616 13280 8125 13308
rect 7616 13268 7622 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 7466 13200 7472 13252
rect 7524 13240 7530 13252
rect 8220 13240 8248 13271
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9640 13280 9689 13308
rect 9640 13268 9646 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 9677 13271 9735 13277
rect 10704 13280 11253 13308
rect 7524 13212 8248 13240
rect 7524 13200 7530 13212
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 2961 13175 3019 13181
rect 2961 13172 2973 13175
rect 2372 13144 2973 13172
rect 2372 13132 2378 13144
rect 2961 13141 2973 13144
rect 3007 13141 3019 13175
rect 2961 13135 3019 13141
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 10704 13172 10732 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 11348 13308 11376 13348
rect 12710 13336 12716 13348
rect 12768 13336 12774 13388
rect 13464 13385 13492 13416
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14550 13444 14556 13456
rect 14056 13416 14556 13444
rect 14056 13404 14062 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 15436 13416 15669 13444
rect 15436 13404 15442 13416
rect 15657 13413 15669 13416
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13345 13507 13379
rect 13449 13339 13507 13345
rect 13716 13379 13774 13385
rect 13716 13345 13728 13379
rect 13762 13376 13774 13379
rect 14182 13376 14188 13388
rect 13762 13348 14188 13376
rect 13762 13345 13774 13348
rect 13716 13339 13774 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 11348 13280 11468 13308
rect 11241 13271 11299 13277
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11333 13243 11391 13249
rect 11333 13240 11345 13243
rect 11204 13212 11345 13240
rect 11204 13200 11210 13212
rect 11333 13209 11345 13212
rect 11379 13209 11391 13243
rect 11440 13240 11468 13280
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11572 13280 11897 13308
rect 11572 13268 11578 13280
rect 11885 13277 11897 13280
rect 11931 13308 11943 13311
rect 12897 13311 12955 13317
rect 12897 13308 12909 13311
rect 11931 13280 12909 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12897 13277 12909 13280
rect 12943 13277 12955 13311
rect 15930 13308 15936 13320
rect 15843 13280 15936 13308
rect 12897 13271 12955 13277
rect 15930 13268 15936 13280
rect 15988 13308 15994 13320
rect 16390 13308 16396 13320
rect 15988 13280 16396 13308
rect 15988 13268 15994 13280
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 12342 13240 12348 13252
rect 11440 13212 12348 13240
rect 11333 13203 11391 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 14829 13243 14887 13249
rect 14829 13209 14841 13243
rect 14875 13240 14887 13243
rect 15102 13240 15108 13252
rect 14875 13212 15108 13240
rect 14875 13209 14887 13212
rect 14829 13203 14887 13209
rect 15102 13200 15108 13212
rect 15160 13240 15166 13252
rect 16022 13240 16028 13252
rect 15160 13212 16028 13240
rect 15160 13200 15166 13212
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 5408 13144 10732 13172
rect 5408 13132 5414 13144
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 11020 13144 11069 13172
rect 11020 13132 11026 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 12161 13175 12219 13181
rect 12161 13172 12173 13175
rect 11287 13144 12173 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 12161 13141 12173 13144
rect 12207 13141 12219 13175
rect 12161 13135 12219 13141
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 17218 13172 17224 13184
rect 15335 13144 17224 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 5166 12968 5172 12980
rect 4847 12940 5172 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5166 12928 5172 12940
rect 5224 12968 5230 12980
rect 6641 12971 6699 12977
rect 6641 12968 6653 12971
rect 5224 12940 6653 12968
rect 5224 12928 5230 12940
rect 6641 12937 6653 12940
rect 6687 12937 6699 12971
rect 6914 12968 6920 12980
rect 6875 12940 6920 12968
rect 6641 12931 6699 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 10594 12968 10600 12980
rect 7024 12940 10600 12968
rect 1670 12860 1676 12912
rect 1728 12900 1734 12912
rect 1728 12872 3648 12900
rect 1728 12860 1734 12872
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12832 2651 12835
rect 2682 12832 2688 12844
rect 2639 12804 2688 12832
rect 2639 12801 2651 12804
rect 2593 12795 2651 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3620 12841 3648 12872
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 7024 12900 7052 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 11882 12968 11888 12980
rect 11664 12940 11888 12968
rect 11664 12928 11670 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12802 12968 12808 12980
rect 12115 12940 12808 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 14182 12968 14188 12980
rect 14143 12940 14188 12968
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 14550 12968 14556 12980
rect 14507 12940 14556 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15473 12971 15531 12977
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 15746 12968 15752 12980
rect 15519 12940 15752 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 7745 12903 7803 12909
rect 7745 12900 7757 12903
rect 4120 12872 7052 12900
rect 7116 12872 7757 12900
rect 4120 12860 4126 12872
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12832 3663 12835
rect 3694 12832 3700 12844
rect 3651 12804 3700 12832
rect 3651 12801 3663 12804
rect 3605 12795 3663 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4212 12804 4445 12832
rect 4212 12792 4218 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5442 12832 5448 12844
rect 4663 12804 5448 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5442 12792 5448 12804
rect 5500 12832 5506 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5500 12804 5549 12832
rect 5500 12792 5506 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7116 12832 7144 12872
rect 7745 12869 7757 12872
rect 7791 12869 7803 12903
rect 7745 12863 7803 12869
rect 7929 12903 7987 12909
rect 7929 12869 7941 12903
rect 7975 12900 7987 12903
rect 8202 12900 8208 12912
rect 7975 12872 8208 12900
rect 7975 12869 7987 12872
rect 7929 12863 7987 12869
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 9766 12900 9772 12912
rect 8312 12872 9772 12900
rect 7466 12832 7472 12844
rect 6687 12804 7144 12832
rect 7427 12804 7472 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 8312 12832 8340 12872
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 7576 12804 8340 12832
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2314 12764 2320 12776
rect 2275 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4387 12736 4813 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 4948 12736 5120 12764
rect 4948 12724 4954 12736
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 5092 12696 5120 12736
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5350 12764 5356 12776
rect 5224 12736 5356 12764
rect 5224 12724 5230 12736
rect 5350 12724 5356 12736
rect 5408 12764 5414 12776
rect 7576 12764 7604 12804
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9640 12804 9873 12832
rect 9640 12792 9646 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 10962 12832 10968 12844
rect 9861 12795 9919 12801
rect 10888 12804 10968 12832
rect 5408 12736 5488 12764
rect 5408 12724 5414 12736
rect 5460 12705 5488 12736
rect 6840 12736 7604 12764
rect 5445 12699 5503 12705
rect 3375 12668 5028 12696
rect 5092 12668 5396 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 5000 12637 5028 12668
rect 5368 12637 5396 12668
rect 5445 12665 5457 12699
rect 5491 12665 5503 12699
rect 5445 12659 5503 12665
rect 2409 12631 2467 12637
rect 2409 12597 2421 12631
rect 2455 12628 2467 12631
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2455 12600 2973 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 2961 12591 3019 12597
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3467 12600 3985 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 3973 12597 3985 12600
rect 4019 12597 4031 12631
rect 3973 12591 4031 12597
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12597 5043 12631
rect 4985 12591 5043 12597
rect 5353 12631 5411 12637
rect 5353 12597 5365 12631
rect 5399 12628 5411 12631
rect 6840 12628 6868 12736
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 10134 12773 10140 12776
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 7708 12736 8125 12764
rect 7708 12724 7714 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 10128 12764 10140 12773
rect 10047 12736 10140 12764
rect 8113 12727 8171 12733
rect 10128 12727 10140 12736
rect 10192 12764 10198 12776
rect 10888 12764 10916 12804
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12158 12832 12164 12844
rect 11756 12804 12164 12832
rect 11756 12792 11762 12804
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 14200 12832 14228 12928
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14200 12804 15025 12832
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 16022 12832 16028 12844
rect 15983 12804 16028 12832
rect 15013 12795 15071 12801
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 12250 12764 12256 12776
rect 10192 12736 10916 12764
rect 12211 12736 12256 12764
rect 10134 12724 10140 12727
rect 10192 12724 10198 12736
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12452 12736 12817 12764
rect 12452 12708 12480 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 15194 12764 15200 12776
rect 12805 12727 12863 12733
rect 12912 12736 15200 12764
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 10686 12696 10692 12708
rect 7331 12668 10692 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 12434 12696 12440 12708
rect 11204 12668 12440 12696
rect 11204 12656 11210 12668
rect 12434 12656 12440 12668
rect 12492 12656 12498 12708
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12912 12696 12940 12736
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15838 12764 15844 12776
rect 15799 12736 15844 12764
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 12584 12668 12940 12696
rect 13072 12699 13130 12705
rect 12584 12656 12590 12668
rect 13072 12665 13084 12699
rect 13118 12696 13130 12699
rect 13722 12696 13728 12708
rect 13118 12668 13728 12696
rect 13118 12665 13130 12668
rect 13072 12659 13130 12665
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 14921 12699 14979 12705
rect 14921 12696 14933 12699
rect 13872 12668 14933 12696
rect 13872 12656 13878 12668
rect 14921 12665 14933 12668
rect 14967 12665 14979 12699
rect 14921 12659 14979 12665
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 15933 12699 15991 12705
rect 15933 12696 15945 12699
rect 15804 12668 15945 12696
rect 15804 12656 15810 12668
rect 15933 12665 15945 12668
rect 15979 12665 15991 12699
rect 15933 12659 15991 12665
rect 5399 12600 6868 12628
rect 7377 12631 7435 12637
rect 5399 12597 5411 12600
rect 5353 12591 5411 12597
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7558 12628 7564 12640
rect 7423 12600 7564 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 10134 12628 10140 12640
rect 7791 12600 10140 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 11238 12628 11244 12640
rect 11199 12600 11244 12628
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12158 12628 12164 12640
rect 11848 12600 12164 12628
rect 11848 12588 11854 12600
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 14550 12588 14556 12640
rect 14608 12628 14614 12640
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 14608 12600 14841 12628
rect 14608 12588 14614 12600
rect 14829 12597 14841 12600
rect 14875 12597 14887 12631
rect 14829 12591 14887 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 5445 12427 5503 12433
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5534 12424 5540 12436
rect 5491 12396 5540 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 7098 12424 7104 12436
rect 7059 12396 7104 12424
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 7558 12424 7564 12436
rect 7515 12396 7564 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 8527 12396 10057 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 10045 12393 10057 12396
rect 10091 12393 10103 12427
rect 10045 12387 10103 12393
rect 10137 12427 10195 12433
rect 10137 12393 10149 12427
rect 10183 12424 10195 12427
rect 10410 12424 10416 12436
rect 10183 12396 10416 12424
rect 10183 12393 10195 12396
rect 10137 12387 10195 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 10928 12396 12725 12424
rect 10928 12384 10934 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13357 12427 13415 12433
rect 12860 12396 12905 12424
rect 12860 12384 12866 12396
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 13814 12424 13820 12436
rect 13403 12396 13820 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 1670 12316 1676 12368
rect 1728 12365 1734 12368
rect 1728 12359 1792 12365
rect 1728 12325 1746 12359
rect 1780 12325 1792 12359
rect 4062 12356 4068 12368
rect 3975 12328 4068 12356
rect 1728 12319 1792 12325
rect 1728 12316 1734 12319
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12288 1547 12291
rect 3988 12288 4016 12328
rect 4062 12316 4068 12328
rect 4120 12356 4126 12368
rect 5718 12356 5724 12368
rect 4120 12328 5724 12356
rect 4120 12316 4126 12328
rect 5718 12316 5724 12328
rect 5776 12316 5782 12368
rect 7929 12359 7987 12365
rect 7929 12325 7941 12359
rect 7975 12356 7987 12359
rect 8386 12356 8392 12368
rect 7975 12328 8392 12356
rect 7975 12325 7987 12328
rect 7929 12319 7987 12325
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 10594 12356 10600 12368
rect 8628 12328 10600 12356
rect 8628 12316 8634 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 10956 12359 11014 12365
rect 10956 12325 10968 12359
rect 11002 12356 11014 12359
rect 11238 12356 11244 12368
rect 11002 12328 11244 12356
rect 11002 12325 11014 12328
rect 10956 12319 11014 12325
rect 11238 12316 11244 12328
rect 11296 12356 11302 12368
rect 11296 12328 12940 12356
rect 11296 12316 11302 12328
rect 1535 12260 4016 12288
rect 1535 12257 1547 12260
rect 1489 12251 1547 12257
rect 3988 12220 4016 12260
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4332 12291 4390 12297
rect 4332 12288 4344 12291
rect 4212 12260 4344 12288
rect 4212 12248 4218 12260
rect 4332 12257 4344 12260
rect 4378 12288 4390 12291
rect 5442 12288 5448 12300
rect 4378 12260 5448 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5988 12291 6046 12297
rect 5988 12257 6000 12291
rect 6034 12288 6046 12291
rect 6454 12288 6460 12300
rect 6034 12260 6460 12288
rect 6034 12257 6046 12260
rect 5988 12251 6046 12257
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 7883 12260 8248 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3988 12192 4077 12220
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 5718 12220 5724 12232
rect 5679 12192 5724 12220
rect 4065 12183 4123 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 8018 12180 8024 12232
rect 8076 12220 8082 12232
rect 8220 12220 8248 12260
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 8849 12291 8907 12297
rect 8849 12288 8861 12291
rect 8352 12260 8861 12288
rect 8352 12248 8358 12260
rect 8849 12257 8861 12260
rect 8895 12257 8907 12291
rect 8849 12251 8907 12257
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10468 12260 10701 12288
rect 10468 12248 10474 12260
rect 10689 12257 10701 12260
rect 10735 12288 10747 12291
rect 10778 12288 10784 12300
rect 10735 12260 10784 12288
rect 10735 12257 10747 12260
rect 10689 12251 10747 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 8478 12220 8484 12232
rect 8076 12192 8121 12220
rect 8220 12192 8484 12220
rect 8076 12180 8082 12192
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 10042 12220 10048 12232
rect 9171 12192 10048 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12220 12219 12223
rect 12802 12220 12808 12232
rect 12207 12192 12808 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 12912 12229 12940 12328
rect 13538 12316 13544 12368
rect 13596 12356 13602 12368
rect 14274 12356 14280 12368
rect 13596 12328 14280 12356
rect 13596 12316 13602 12328
rect 14274 12316 14280 12328
rect 14332 12356 14338 12368
rect 15102 12356 15108 12368
rect 14332 12328 15108 12356
rect 14332 12316 14338 12328
rect 15102 12316 15108 12328
rect 15160 12356 15166 12368
rect 15160 12328 15332 12356
rect 15160 12316 15166 12328
rect 15304 12297 15332 12328
rect 13725 12291 13783 12297
rect 13725 12288 13737 12291
rect 13004 12260 13737 12288
rect 13004 12232 13032 12260
rect 13725 12257 13737 12260
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15556 12291 15614 12297
rect 15556 12257 15568 12291
rect 15602 12288 15614 12291
rect 17310 12288 17316 12300
rect 15602 12260 17316 12288
rect 15602 12257 15614 12260
rect 15556 12251 15614 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13817 12223 13875 12229
rect 13817 12220 13829 12223
rect 13087 12192 13829 12220
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 13087 12152 13115 12192
rect 13817 12189 13829 12192
rect 13863 12189 13875 12223
rect 13817 12183 13875 12189
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12189 13967 12223
rect 13909 12183 13967 12189
rect 12032 12124 13115 12152
rect 12032 12112 12038 12124
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 13924 12152 13952 12183
rect 13780 12124 13952 12152
rect 13780 12112 13786 12124
rect 2498 12044 2504 12096
rect 2556 12084 2562 12096
rect 2682 12084 2688 12096
rect 2556 12056 2688 12084
rect 2556 12044 2562 12056
rect 2682 12044 2688 12056
rect 2740 12084 2746 12096
rect 2869 12087 2927 12093
rect 2869 12084 2881 12087
rect 2740 12056 2881 12084
rect 2740 12044 2746 12056
rect 2869 12053 2881 12056
rect 2915 12053 2927 12087
rect 2869 12047 2927 12053
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 5258 12084 5264 12096
rect 3476 12056 5264 12084
rect 3476 12044 3482 12056
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 11882 12084 11888 12096
rect 9723 12056 11888 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 12115 12056 12173 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 12161 12047 12219 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 16850 12084 16856 12096
rect 16715 12056 16856 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 3326 11880 3332 11892
rect 2639 11852 3332 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 3602 11880 3608 11892
rect 3563 11852 3608 11880
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 6454 11880 6460 11892
rect 4120 11852 6316 11880
rect 6367 11852 6460 11880
rect 4120 11840 4126 11852
rect 6288 11812 6316 11852
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 8018 11880 8024 11892
rect 6512 11852 8024 11880
rect 6512 11840 6518 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8294 11880 8300 11892
rect 8255 11852 8300 11880
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 11606 11880 11612 11892
rect 9784 11852 11612 11880
rect 9674 11812 9680 11824
rect 6288 11784 9680 11812
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 4154 11744 4160 11756
rect 3283 11716 4160 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 5000 11716 5212 11744
rect 1670 11676 1676 11688
rect 1631 11648 1676 11676
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3970 11676 3976 11688
rect 2924 11648 3976 11676
rect 2924 11636 2930 11648
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 5000 11676 5028 11716
rect 4120 11648 5028 11676
rect 5077 11679 5135 11685
rect 4120 11636 4126 11648
rect 5077 11645 5089 11679
rect 5123 11645 5135 11679
rect 5184 11676 5212 11716
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 7800 11716 8769 11744
rect 7800 11704 7806 11716
rect 8757 11713 8769 11716
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 9122 11744 9128 11756
rect 8987 11716 9128 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9784 11753 9812 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 12066 11880 12072 11892
rect 11848 11852 12072 11880
rect 11848 11840 11854 11852
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 13538 11880 13544 11892
rect 12452 11852 13544 11880
rect 10321 11815 10379 11821
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 11146 11812 11152 11824
rect 10367 11784 11152 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 12158 11812 12164 11824
rect 11808 11784 12164 11812
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9950 11744 9956 11756
rect 9911 11716 9956 11744
rect 9769 11707 9827 11713
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10962 11744 10968 11756
rect 10923 11716 10968 11744
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11808 11744 11836 11784
rect 12158 11772 12164 11784
rect 12216 11772 12222 11824
rect 12452 11756 12480 11852
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13780 11852 13829 11880
rect 13780 11840 13786 11852
rect 13817 11849 13829 11852
rect 13863 11849 13875 11883
rect 13817 11843 13875 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14550 11880 14556 11892
rect 14139 11852 14556 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 11716 11716 11836 11744
rect 11977 11747 12035 11753
rect 7466 11676 7472 11688
rect 5184 11648 7472 11676
rect 5077 11639 5135 11645
rect 1486 11568 1492 11620
rect 1544 11608 1550 11620
rect 1949 11611 2007 11617
rect 1949 11608 1961 11611
rect 1544 11580 1961 11608
rect 1544 11568 1550 11580
rect 1949 11577 1961 11580
rect 1995 11577 2007 11611
rect 1949 11571 2007 11577
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 4617 11611 4675 11617
rect 4617 11608 4629 11611
rect 3007 11580 4629 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 4617 11577 4629 11580
rect 4663 11577 4675 11611
rect 4617 11571 4675 11577
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3418 11540 3424 11552
rect 3099 11512 3424 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 4062 11540 4068 11552
rect 3660 11512 4068 11540
rect 3660 11500 3666 11512
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 5092 11540 5120 11639
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10318 11676 10324 11688
rect 9723 11648 10324 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 5350 11617 5356 11620
rect 5344 11608 5356 11617
rect 5311 11580 5356 11608
rect 5344 11571 5356 11580
rect 5350 11568 5356 11571
rect 5408 11568 5414 11620
rect 8036 11608 8064 11639
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 11716 11685 11744 11716
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12066 11744 12072 11756
rect 12023 11716 12072 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12066 11704 12072 11716
rect 12124 11744 12130 11756
rect 12124 11716 12296 11744
rect 12124 11704 12130 11716
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11882 11676 11888 11688
rect 11839 11648 11888 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12268 11676 12296 11716
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 13832 11744 13860 11843
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 12492 11716 12537 11744
rect 13832 11716 14657 11744
rect 12492 11704 12498 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 14645 11707 14703 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 17310 11744 17316 11756
rect 17271 11716 17316 11744
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 12268 11648 14780 11676
rect 10689 11611 10747 11617
rect 8036 11580 10640 11608
rect 6822 11540 6828 11552
rect 4212 11512 5120 11540
rect 6783 11512 6828 11540
rect 4212 11500 4218 11512
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7650 11540 7656 11552
rect 7156 11512 7656 11540
rect 7156 11500 7162 11512
rect 7650 11500 7656 11512
rect 7708 11540 7714 11552
rect 7837 11543 7895 11549
rect 7837 11540 7849 11543
rect 7708 11512 7849 11540
rect 7708 11500 7714 11512
rect 7837 11509 7849 11512
rect 7883 11509 7895 11543
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 7837 11503 7895 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9272 11512 9321 11540
rect 9272 11500 9278 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 10612 11540 10640 11580
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 12526 11608 12532 11620
rect 10735 11580 12532 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12704 11611 12762 11617
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 12802 11608 12808 11620
rect 12750 11580 12808 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 14366 11608 14372 11620
rect 13596 11580 14372 11608
rect 13596 11568 13602 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14553 11611 14611 11617
rect 14553 11577 14565 11611
rect 14599 11608 14611 11611
rect 14642 11608 14648 11620
rect 14599 11580 14648 11608
rect 14599 11577 14611 11580
rect 14553 11571 14611 11577
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 11054 11540 11060 11552
rect 10612 11512 11060 11540
rect 9309 11503 9367 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11330 11540 11336 11552
rect 11291 11512 11336 11540
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 12544 11540 12572 11568
rect 13262 11540 13268 11552
rect 12544 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14752 11540 14780 11648
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 15712 11648 17141 11676
rect 15712 11636 15718 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 17218 11636 17224 11688
rect 17276 11676 17282 11688
rect 17276 11648 17321 11676
rect 17276 11636 17282 11648
rect 15372 11611 15430 11617
rect 15372 11577 15384 11611
rect 15418 11608 15430 11611
rect 16850 11608 16856 11620
rect 15418 11580 16856 11608
rect 15418 11577 15430 11580
rect 15372 11571 15430 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 14752 11512 16497 11540
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16758 11540 16764 11552
rect 16719 11512 16764 11540
rect 16485 11503 16543 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 2774 11336 2780 11348
rect 1719 11308 2780 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 6270 11336 6276 11348
rect 4120 11308 6276 11336
rect 4120 11296 4126 11308
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6822 11336 6828 11348
rect 6503 11308 6828 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 9214 11336 9220 11348
rect 9175 11308 9220 11336
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11112 11308 11437 11336
rect 11112 11296 11118 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11974 11336 11980 11348
rect 11935 11308 11980 11336
rect 11425 11299 11483 11305
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12400 11308 12449 11336
rect 12400 11296 12406 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 12986 11336 12992 11348
rect 12851 11308 12992 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13262 11336 13268 11348
rect 13223 11308 13268 11336
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 14458 11336 14464 11348
rect 13679 11308 14464 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15654 11336 15660 11348
rect 15335 11308 15660 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16298 11336 16304 11348
rect 16259 11308 16304 11336
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 16758 11336 16764 11348
rect 16719 11308 16764 11336
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 2308 11271 2366 11277
rect 2308 11237 2320 11271
rect 2354 11268 2366 11271
rect 2498 11268 2504 11280
rect 2354 11240 2504 11268
rect 2354 11237 2366 11240
rect 2308 11231 2366 11237
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 4332 11271 4390 11277
rect 3936 11240 4292 11268
rect 3936 11228 3942 11240
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 2056 11172 4077 11200
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2056 11141 2084 11172
rect 4065 11169 4077 11172
rect 4111 11200 4123 11203
rect 4154 11200 4160 11212
rect 4111 11172 4160 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4264 11200 4292 11240
rect 4332 11237 4344 11271
rect 4378 11268 4390 11271
rect 6178 11268 6184 11280
rect 4378 11240 6184 11268
rect 4378 11237 4390 11240
rect 4332 11231 4390 11237
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 8662 11228 8668 11280
rect 8720 11268 8726 11280
rect 9677 11271 9735 11277
rect 9677 11268 9689 11271
rect 8720 11240 9689 11268
rect 8720 11228 8726 11240
rect 9677 11237 9689 11240
rect 9723 11237 9735 11271
rect 9677 11231 9735 11237
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 10502 11268 10508 11280
rect 10183 11240 10508 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 10502 11228 10508 11240
rect 10560 11228 10566 11280
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12584 11240 13185 11268
rect 12584 11228 12590 11240
rect 13173 11237 13185 11240
rect 13219 11268 13231 11271
rect 13538 11268 13544 11280
rect 13219 11240 13544 11268
rect 13219 11237 13231 11240
rect 13173 11231 13231 11237
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 13648 11240 14136 11268
rect 4890 11200 4896 11212
rect 4264 11172 4896 11200
rect 4890 11160 4896 11172
rect 4948 11200 4954 11212
rect 4948 11172 5120 11200
rect 4948 11160 4954 11172
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 2004 11104 2053 11132
rect 2004 11092 2010 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 5092 11132 5120 11172
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 5776 11172 7113 11200
rect 5776 11160 5782 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 7368 11203 7426 11209
rect 7368 11169 7380 11203
rect 7414 11200 7426 11203
rect 9125 11203 9183 11209
rect 7414 11172 8248 11200
rect 7414 11169 7426 11172
rect 7368 11163 7426 11169
rect 8220 11144 8248 11172
rect 9125 11169 9137 11203
rect 9171 11200 9183 11203
rect 10042 11200 10048 11212
rect 9171 11172 10048 11200
rect 9171 11169 9183 11172
rect 9125 11163 9183 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 12158 11160 12164 11212
rect 12216 11200 12222 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 12216 11172 12357 11200
rect 12216 11160 12222 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13648 11200 13676 11240
rect 13998 11200 14004 11212
rect 13320 11172 13676 11200
rect 13959 11172 14004 11200
rect 13320 11160 13326 11172
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14108 11200 14136 11240
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 15528 11240 15792 11268
rect 15528 11228 15534 11240
rect 15764 11209 15792 11240
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 14108 11172 15669 11200
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 15838 11200 15844 11212
rect 15795 11172 15844 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 5092 11104 6561 11132
rect 2041 11095 2099 11101
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6549 11095 6607 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8260 11104 9321 11132
rect 8260 11092 8266 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 12802 11132 12808 11144
rect 12667 11104 12808 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 12802 11092 12808 11104
rect 12860 11132 12866 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 12860 11104 13369 11132
rect 12860 11092 12866 11104
rect 13357 11101 13369 11104
rect 13403 11132 13415 11135
rect 13538 11132 13544 11144
rect 13403 11104 13544 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13872 11104 14105 11132
rect 13872 11092 13878 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14240 11104 14289 11132
rect 14240 11092 14246 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 15672 11132 15700 11163
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16666 11200 16672 11212
rect 16627 11172 16672 11200
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 15930 11132 15936 11144
rect 15672 11104 15792 11132
rect 15891 11104 15936 11132
rect 14277 11095 14335 11101
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5920 11036 6224 11064
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3292 10968 3433 10996
rect 3292 10956 3298 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 3421 10959 3479 10965
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 5920 10996 5948 11036
rect 6086 10996 6092 11008
rect 4120 10968 5948 10996
rect 6047 10968 6092 10996
rect 4120 10956 4126 10968
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 6196 10996 6224 11036
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10502 11064 10508 11076
rect 9732 11036 10508 11064
rect 9732 11024 9738 11036
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 12894 11064 12900 11076
rect 11388 11036 12900 11064
rect 11388 11024 11394 11036
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 15764 11064 15792 11104
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16850 11132 16856 11144
rect 16811 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 17402 11064 17408 11076
rect 15764 11036 17408 11064
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 7466 10996 7472 11008
rect 6196 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10996 7530 11008
rect 7742 10996 7748 11008
rect 7524 10968 7748 10996
rect 7524 10956 7530 10968
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 8570 10996 8576 11008
rect 8527 10968 8576 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 16942 10996 16948 11008
rect 11664 10968 16948 10996
rect 11664 10956 11670 10968
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1670 10792 1676 10804
rect 1627 10764 1676 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 3568 10764 3801 10792
rect 3568 10752 3574 10764
rect 3789 10761 3801 10764
rect 3835 10761 3847 10795
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 3789 10755 3847 10761
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 6549 10795 6607 10801
rect 6549 10761 6561 10795
rect 6595 10792 6607 10795
rect 8202 10792 8208 10804
rect 6595 10764 8208 10792
rect 6595 10761 6607 10764
rect 6549 10755 6607 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 13449 10795 13507 10801
rect 10284 10764 13400 10792
rect 10284 10752 10290 10764
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 9861 10727 9919 10733
rect 9861 10724 9873 10727
rect 9732 10696 9873 10724
rect 9732 10684 9738 10696
rect 9861 10693 9873 10696
rect 9907 10724 9919 10727
rect 10962 10724 10968 10736
rect 9907 10696 10968 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10693 12495 10727
rect 13372 10724 13400 10764
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 14550 10792 14556 10804
rect 13495 10764 14556 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 15841 10795 15899 10801
rect 15841 10761 15853 10795
rect 15887 10792 15899 10795
rect 16666 10792 16672 10804
rect 15887 10764 16672 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 13372 10696 14780 10724
rect 12437 10687 12495 10693
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 3234 10656 3240 10668
rect 3195 10628 3240 10656
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4982 10656 4988 10668
rect 4764 10628 4988 10656
rect 4764 10616 4770 10628
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5350 10656 5356 10668
rect 5311 10628 5356 10656
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6411 10628 6561 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10008 10628 10793 10656
rect 10008 10616 10014 10628
rect 10781 10625 10793 10628
rect 10827 10656 10839 10659
rect 11974 10656 11980 10668
rect 10827 10628 11980 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12452 10656 12480 10687
rect 12894 10656 12900 10668
rect 12452 10628 12756 10656
rect 12855 10628 12900 10656
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 3970 10588 3976 10600
rect 3651 10560 3976 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 6086 10588 6092 10600
rect 6047 10560 6092 10588
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 2041 10523 2099 10529
rect 2041 10489 2053 10523
rect 2087 10520 2099 10523
rect 2866 10520 2872 10532
rect 2087 10492 2872 10520
rect 2087 10489 2099 10492
rect 2041 10483 2099 10489
rect 2866 10480 2872 10492
rect 2924 10480 2930 10532
rect 2961 10523 3019 10529
rect 2961 10489 2973 10523
rect 3007 10520 3019 10523
rect 3694 10520 3700 10532
rect 3007 10492 3700 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3694 10480 3700 10492
rect 3752 10480 3758 10532
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5442 10520 5448 10532
rect 5040 10492 5448 10520
rect 5040 10480 5046 10492
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 6914 10520 6920 10532
rect 5736 10492 6920 10520
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1636 10424 1961 10452
rect 1636 10412 1642 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 1949 10415 2007 10421
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 2188 10424 2605 10452
rect 2188 10412 2194 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3326 10452 3332 10464
rect 3099 10424 3332 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3326 10412 3332 10424
rect 3384 10452 3390 10464
rect 3786 10452 3792 10464
rect 3384 10424 3792 10452
rect 3384 10412 3390 10424
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5626 10452 5632 10464
rect 5215 10424 5632 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5736 10461 5764 10492
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 7092 10523 7150 10529
rect 7092 10520 7104 10523
rect 7024 10492 7104 10520
rect 5721 10455 5779 10461
rect 5721 10421 5733 10455
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 6086 10412 6092 10464
rect 6144 10452 6150 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6144 10424 6193 10452
rect 6144 10412 6150 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7024 10452 7052 10492
rect 7092 10489 7104 10492
rect 7138 10520 7150 10523
rect 8496 10520 8524 10551
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 8737 10591 8795 10597
rect 8737 10588 8749 10591
rect 8628 10560 8749 10588
rect 8628 10548 8634 10560
rect 8737 10557 8749 10560
rect 8783 10557 8795 10591
rect 8737 10551 8795 10557
rect 10410 10520 10416 10532
rect 7138 10492 8432 10520
rect 8496 10492 10416 10520
rect 7138 10489 7150 10492
rect 7092 10483 7150 10489
rect 6788 10424 7052 10452
rect 8404 10452 8432 10492
rect 10410 10480 10416 10492
rect 10468 10480 10474 10532
rect 10505 10523 10563 10529
rect 10505 10489 10517 10523
rect 10551 10520 10563 10523
rect 12158 10520 12164 10532
rect 10551 10492 12164 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 12728 10520 12756 10628
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13044 10628 13089 10656
rect 13044 10616 13050 10628
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13596 10628 14013 10656
rect 13596 10616 13602 10628
rect 14001 10625 14013 10628
rect 14047 10656 14059 10659
rect 14182 10656 14188 10668
rect 14047 10628 14188 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 14752 10656 14780 10696
rect 16114 10684 16120 10736
rect 16172 10724 16178 10736
rect 16850 10724 16856 10736
rect 16172 10696 16856 10724
rect 16172 10684 16178 10696
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 15286 10656 15292 10668
rect 14752 10628 15292 10656
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 13906 10588 13912 10600
rect 13863 10560 13912 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 14550 10520 14556 10532
rect 12728 10492 14556 10520
rect 14550 10480 14556 10492
rect 14608 10480 14614 10532
rect 9950 10452 9956 10464
rect 8404 10424 9956 10452
rect 6788 10412 6794 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10594 10452 10600 10464
rect 10555 10424 10600 10452
rect 10594 10412 10600 10424
rect 10652 10452 10658 10464
rect 12618 10452 12624 10464
rect 10652 10424 12624 10452
rect 10652 10412 10658 10424
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 13722 10452 13728 10464
rect 13596 10424 13728 10452
rect 13596 10412 13602 10424
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 13909 10455 13967 10461
rect 13909 10421 13921 10455
rect 13955 10452 13967 10455
rect 14752 10452 14780 10628
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 15930 10656 15936 10668
rect 15519 10628 15936 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16666 10656 16672 10668
rect 16531 10628 16672 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16666 10616 16672 10628
rect 16724 10656 16730 10668
rect 17310 10656 17316 10668
rect 16724 10628 17316 10656
rect 16724 10616 16730 10628
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 16209 10523 16267 10529
rect 16209 10520 16221 10523
rect 14844 10492 16221 10520
rect 14844 10461 14872 10492
rect 16209 10489 16221 10492
rect 16255 10489 16267 10523
rect 16209 10483 16267 10489
rect 13955 10424 14780 10452
rect 14829 10455 14887 10461
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14829 10421 14841 10455
rect 14875 10421 14887 10455
rect 14829 10415 14887 10421
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 15160 10424 15209 10452
rect 15160 10412 15166 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15378 10452 15384 10464
rect 15335 10424 15384 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 16298 10452 16304 10464
rect 16259 10424 16304 10452
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2041 10251 2099 10257
rect 2041 10217 2053 10251
rect 2087 10248 2099 10251
rect 2593 10251 2651 10257
rect 2593 10248 2605 10251
rect 2087 10220 2605 10248
rect 2087 10217 2099 10220
rect 2041 10211 2099 10217
rect 2593 10217 2605 10220
rect 2639 10217 2651 10251
rect 2958 10248 2964 10260
rect 2871 10220 2964 10248
rect 2593 10211 2651 10217
rect 2958 10208 2964 10220
rect 3016 10248 3022 10260
rect 3142 10248 3148 10260
rect 3016 10220 3148 10248
rect 3016 10208 3022 10220
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 4798 10248 4804 10260
rect 3528 10220 4804 10248
rect 1949 10183 2007 10189
rect 1949 10149 1961 10183
rect 1995 10180 2007 10183
rect 2130 10180 2136 10192
rect 1995 10152 2136 10180
rect 1995 10149 2007 10152
rect 1949 10143 2007 10149
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 3053 10183 3111 10189
rect 3053 10149 3065 10183
rect 3099 10180 3111 10183
rect 3528 10180 3556 10220
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5408 10220 5825 10248
rect 5408 10208 5414 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 5813 10211 5871 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 6972 10220 8493 10248
rect 6972 10208 6978 10220
rect 8481 10217 8493 10220
rect 8527 10217 8539 10251
rect 8481 10211 8539 10217
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8754 10248 8760 10260
rect 8619 10220 8760 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12250 10248 12256 10260
rect 12207 10220 12256 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 12676 10220 13952 10248
rect 12676 10208 12682 10220
rect 3099 10152 3556 10180
rect 3099 10149 3111 10152
rect 3053 10143 3111 10149
rect 3160 10124 3188 10152
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 13538 10180 13544 10192
rect 4120 10152 13544 10180
rect 4120 10140 4126 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 3142 10072 3148 10124
rect 3200 10072 3206 10124
rect 4700 10115 4758 10121
rect 4700 10081 4712 10115
rect 4746 10112 4758 10115
rect 5258 10112 5264 10124
rect 4746 10084 5264 10112
rect 4746 10081 4758 10084
rect 4700 10075 4758 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 6457 10115 6515 10121
rect 6457 10112 6469 10115
rect 5500 10084 6469 10112
rect 5500 10072 5506 10084
rect 6457 10081 6469 10084
rect 6503 10081 6515 10115
rect 6457 10075 6515 10081
rect 7469 10115 7527 10121
rect 7469 10081 7481 10115
rect 7515 10112 7527 10115
rect 9030 10112 9036 10124
rect 7515 10084 9036 10112
rect 7515 10081 7527 10084
rect 7469 10075 7527 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10778 10121 10784 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10468 10084 10517 10112
rect 10468 10072 10474 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10772 10112 10784 10121
rect 10739 10084 10784 10112
rect 10505 10075 10563 10081
rect 10772 10075 10784 10084
rect 10778 10072 10784 10075
rect 10836 10072 10842 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 11112 10084 12357 10112
rect 11112 10072 11118 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12492 10084 12633 10112
rect 12492 10072 12498 10084
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 12888 10115 12946 10121
rect 12888 10081 12900 10115
rect 12934 10112 12946 10115
rect 13814 10112 13820 10124
rect 12934 10084 13820 10112
rect 12934 10081 12946 10084
rect 12888 10075 12946 10081
rect 13814 10072 13820 10084
rect 13872 10072 13878 10124
rect 13924 10112 13952 10220
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 14056 10220 14289 10248
rect 14056 10208 14062 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 14277 10211 14335 10217
rect 14737 10251 14795 10257
rect 14737 10217 14749 10251
rect 14783 10248 14795 10251
rect 15102 10248 15108 10260
rect 14783 10220 15108 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 16666 10248 16672 10260
rect 16627 10220 16672 10248
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 15556 10183 15614 10189
rect 14200 10152 15516 10180
rect 14200 10112 14228 10152
rect 13924 10084 14228 10112
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 15378 10112 15384 10124
rect 15335 10084 15384 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 15378 10072 15384 10084
rect 15436 10072 15442 10124
rect 15488 10112 15516 10152
rect 15556 10149 15568 10183
rect 15602 10180 15614 10183
rect 15930 10180 15936 10192
rect 15602 10152 15936 10180
rect 15602 10149 15614 10152
rect 15556 10143 15614 10149
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 17034 10112 17040 10124
rect 15488 10084 17040 10112
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 3234 10044 3240 10056
rect 3195 10016 3240 10044
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4212 10016 4445 10044
rect 4212 10004 4218 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4448 9908 4476 10007
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 5592 10016 6561 10044
rect 5592 10004 5598 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6730 10044 6736 10056
rect 6691 10016 6736 10044
rect 6549 10007 6607 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7558 10044 7564 10056
rect 7519 10016 7564 10044
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8202 10044 8208 10056
rect 7791 10016 8208 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8628 10016 8677 10044
rect 8628 10004 8634 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 5684 9948 7113 9976
rect 5684 9936 5690 9948
rect 7101 9945 7113 9948
rect 7147 9945 7159 9979
rect 7101 9939 7159 9945
rect 11885 9979 11943 9985
rect 11885 9945 11897 9979
rect 11931 9976 11943 9979
rect 12342 9976 12348 9988
rect 11931 9948 12348 9976
rect 11931 9945 11943 9948
rect 11885 9939 11943 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 5350 9908 5356 9920
rect 4448 9880 5356 9908
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 11606 9908 11612 9920
rect 8159 9880 11612 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 12032 9880 14013 9908
rect 12032 9868 12038 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 14001 9871 14059 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 7469 9707 7527 9713
rect 4120 9676 7420 9704
rect 4120 9664 4126 9676
rect 4617 9639 4675 9645
rect 4617 9605 4629 9639
rect 4663 9636 4675 9639
rect 5074 9636 5080 9648
rect 4663 9608 5080 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6914 9636 6920 9648
rect 5868 9608 6920 9636
rect 5868 9596 5874 9608
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 7392 9636 7420 9676
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7558 9704 7564 9716
rect 7515 9676 7564 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 14366 9704 14372 9716
rect 7668 9676 14372 9704
rect 7668 9636 7696 9676
rect 14366 9664 14372 9676
rect 14424 9704 14430 9716
rect 15746 9704 15752 9716
rect 14424 9676 15752 9704
rect 14424 9664 14430 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 7392 9608 7696 9636
rect 10045 9639 10103 9645
rect 10045 9605 10057 9639
rect 10091 9636 10103 9639
rect 12434 9636 12440 9648
rect 10091 9608 10171 9636
rect 10091 9605 10103 9608
rect 10045 9599 10103 9605
rect 10143 9580 10171 9608
rect 10244 9608 12440 9636
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 5258 9568 5264 9580
rect 5171 9540 5264 9568
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 6144 9540 6193 9568
rect 6144 9528 6150 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7800 9540 8033 9568
rect 7800 9528 7806 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 2004 9472 2053 9500
rect 2004 9460 2010 9472
rect 2041 9469 2053 9472
rect 2087 9469 2099 9503
rect 2041 9463 2099 9469
rect 2308 9503 2366 9509
rect 2308 9469 2320 9503
rect 2354 9500 2366 9503
rect 3234 9500 3240 9512
rect 2354 9472 3240 9500
rect 2354 9469 2366 9472
rect 2308 9463 2366 9469
rect 3234 9460 3240 9472
rect 3292 9500 3298 9512
rect 4706 9500 4712 9512
rect 3292 9472 4712 9500
rect 3292 9460 3298 9472
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5276 9500 5304 9528
rect 5276 9472 6500 9500
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4120 9404 5089 9432
rect 4120 9392 4126 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 6362 9432 6368 9444
rect 6043 9404 6368 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 6472 9432 6500 9472
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 7156 9472 7205 9500
rect 7156 9460 7162 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7432 9472 7941 9500
rect 7432 9460 7438 9472
rect 7929 9469 7941 9472
rect 7975 9500 7987 9503
rect 8665 9503 8723 9509
rect 7975 9472 8616 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 8202 9432 8208 9444
rect 6472 9404 8208 9432
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 8588 9432 8616 9472
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 8754 9500 8760 9512
rect 8711 9472 8760 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 8932 9503 8990 9509
rect 8932 9469 8944 9503
rect 8978 9500 8990 9503
rect 9674 9500 9680 9512
rect 8978 9472 9680 9500
rect 8978 9469 8990 9472
rect 8932 9463 8990 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10244 9500 10272 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9636 13878 9648
rect 15105 9639 15163 9645
rect 13872 9608 14688 9636
rect 13872 9596 13878 9608
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11112 9540 11529 9568
rect 11112 9528 11118 9540
rect 11517 9537 11529 9540
rect 11563 9568 11575 9571
rect 12066 9568 12072 9580
rect 11563 9540 12072 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12066 9528 12072 9540
rect 12124 9568 12130 9580
rect 14550 9568 14556 9580
rect 12124 9540 12572 9568
rect 14511 9540 14556 9568
rect 12124 9528 12130 9540
rect 10008 9472 10272 9500
rect 10008 9460 10014 9472
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 11333 9503 11391 9509
rect 11333 9500 11345 9503
rect 10560 9472 11345 9500
rect 10560 9460 10566 9472
rect 11333 9469 11345 9472
rect 11379 9469 11391 9503
rect 11333 9463 11391 9469
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 11664 9472 12449 9500
rect 11664 9460 11670 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 14660 9577 14688 9608
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 16298 9636 16304 9648
rect 15151 9608 16304 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9568 15807 9571
rect 15930 9568 15936 9580
rect 15795 9540 15936 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 13078 9500 13084 9512
rect 12544 9472 13084 9500
rect 12437 9463 12495 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 14332 9472 15485 9500
rect 14332 9460 14338 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 11241 9435 11299 9441
rect 8588 9404 11008 9432
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 4982 9364 4988 9376
rect 4943 9336 4988 9364
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5626 9364 5632 9376
rect 5587 9336 5632 9364
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5776 9336 6101 9364
rect 5776 9324 5782 9336
rect 6089 9333 6101 9336
rect 6135 9333 6147 9367
rect 6089 9327 6147 9333
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6696 9336 7021 9364
rect 6696 9324 6702 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 7837 9367 7895 9373
rect 7837 9333 7849 9367
rect 7883 9364 7895 9367
rect 8386 9364 8392 9376
rect 7883 9336 8392 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 8386 9324 8392 9336
rect 8444 9364 8450 9376
rect 10594 9364 10600 9376
rect 8444 9336 10600 9364
rect 8444 9324 8450 9336
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10870 9364 10876 9376
rect 10831 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 10980 9364 11008 9404
rect 11241 9401 11253 9435
rect 11287 9432 11299 9435
rect 11885 9435 11943 9441
rect 11885 9432 11897 9435
rect 11287 9404 11897 9432
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 11885 9401 11897 9404
rect 11931 9401 11943 9435
rect 11885 9395 11943 9401
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 12682 9435 12740 9441
rect 12682 9432 12694 9435
rect 12400 9404 12694 9432
rect 12400 9392 12406 9404
rect 12682 9401 12694 9404
rect 12728 9401 12740 9435
rect 15010 9432 15016 9444
rect 12682 9395 12740 9401
rect 14108 9404 15016 9432
rect 11974 9364 11980 9376
rect 10980 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 14108 9373 14136 9404
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 14093 9367 14151 9373
rect 14093 9333 14105 9367
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14240 9336 14473 9364
rect 14240 9324 14246 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15252 9336 15577 9364
rect 15252 9324 15258 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2280 9132 2789 9160
rect 2280 9120 2286 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 5040 9132 5089 9160
rect 5040 9120 5046 9132
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5077 9123 5135 9129
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5408 9132 5549 9160
rect 5408 9120 5414 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 7193 9163 7251 9169
rect 5537 9123 5595 9129
rect 5644 9132 7144 9160
rect 1664 9095 1722 9101
rect 1664 9061 1676 9095
rect 1710 9092 1722 9095
rect 2130 9092 2136 9104
rect 1710 9064 2136 9092
rect 1710 9061 1722 9064
rect 1664 9055 1722 9061
rect 2130 9052 2136 9064
rect 2188 9092 2194 9104
rect 3418 9092 3424 9104
rect 2188 9064 3424 9092
rect 2188 9052 2194 9064
rect 3418 9052 3424 9064
rect 3476 9052 3482 9104
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 5644 9092 5672 9132
rect 6638 9092 6644 9104
rect 3844 9064 5672 9092
rect 5736 9064 6644 9092
rect 3844 9052 3850 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1946 9024 1952 9036
rect 1443 8996 1952 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 5736 9033 5764 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 4028 8996 4445 9024
rect 4028 8984 4034 8996
rect 4433 8993 4445 8996
rect 4479 8993 4491 9027
rect 4433 8987 4491 8993
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 9024 4583 9027
rect 5721 9027 5779 9033
rect 4571 8996 5672 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5644 8956 5672 8996
rect 5721 8993 5733 9027
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 5902 9024 5908 9036
rect 5859 8996 5908 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6086 9033 6092 9036
rect 6080 9024 6092 9033
rect 6047 8996 6092 9024
rect 6080 8987 6092 8996
rect 6086 8984 6092 8987
rect 6144 8984 6150 9036
rect 7116 9024 7144 9132
rect 7193 9129 7205 9163
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 7208 9092 7236 9123
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7432 9132 7880 9160
rect 7432 9120 7438 9132
rect 7742 9101 7748 9104
rect 7736 9092 7748 9101
rect 7208 9064 7748 9092
rect 7736 9055 7748 9064
rect 7742 9052 7748 9055
rect 7800 9052 7806 9104
rect 7852 9092 7880 9132
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8849 9163 8907 9169
rect 8849 9160 8861 9163
rect 8260 9132 8861 9160
rect 8260 9120 8266 9132
rect 8849 9129 8861 9132
rect 8895 9129 8907 9163
rect 8849 9123 8907 9129
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 10275 9132 10824 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 7852 9064 10057 9092
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 10137 9095 10195 9101
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 10689 9095 10747 9101
rect 10689 9092 10701 9095
rect 10183 9064 10701 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 10689 9061 10701 9064
rect 10735 9061 10747 9095
rect 10796 9092 10824 9132
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 10928 9132 11621 9160
rect 10928 9120 10934 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 11609 9123 11667 9129
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12802 9160 12808 9172
rect 12575 9132 12808 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 14366 9160 14372 9172
rect 14323 9132 14372 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 10796 9064 11713 9092
rect 10689 9055 10747 9061
rect 11701 9061 11713 9064
rect 11747 9061 11759 9095
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 11701 9055 11759 9061
rect 11808 9064 13001 9092
rect 9950 9024 9956 9036
rect 7116 8996 9956 9024
rect 9950 8984 9956 8996
rect 10008 9024 10014 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 10008 8996 10609 9024
rect 10008 8984 10014 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 11808 9024 11836 9064
rect 12989 9061 13001 9064
rect 13035 9092 13047 9095
rect 16206 9092 16212 9104
rect 13035 9064 16212 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 10597 8987 10655 8993
rect 10796 8996 11836 9024
rect 5644 8928 5856 8956
rect 5828 8900 5856 8928
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 6880 8928 7481 8956
rect 6880 8916 6886 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 8720 8928 9781 8956
rect 8720 8916 8726 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10091 8928 10456 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 3936 8860 5672 8888
rect 3936 8848 3942 8860
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3384 8792 4077 8820
rect 3384 8780 3390 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 5644 8820 5672 8860
rect 5810 8848 5816 8900
rect 5868 8848 5874 8900
rect 10318 8888 10324 8900
rect 8404 8860 10324 8888
rect 8404 8820 8432 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 10428 8888 10456 8928
rect 10796 8888 10824 8996
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12526 9024 12532 9036
rect 12032 8996 12532 9024
rect 12032 8984 12038 8996
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8956 10931 8959
rect 11054 8956 11060 8968
rect 10919 8928 11060 8956
rect 10919 8925 10931 8928
rect 10873 8919 10931 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12342 8956 12348 8968
rect 11931 8928 12348 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 12912 8956 12940 8987
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14366 9024 14372 9036
rect 14148 8996 14372 9024
rect 14148 8984 14154 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 13078 8956 13084 8968
rect 12768 8928 12940 8956
rect 13039 8928 13084 8956
rect 12768 8916 12774 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 14461 8959 14519 8965
rect 13596 8928 14320 8956
rect 13596 8916 13602 8928
rect 10428 8860 10824 8888
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 14182 8888 14188 8900
rect 11287 8860 14188 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 14182 8848 14188 8860
rect 14240 8848 14246 8900
rect 14292 8888 14320 8928
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14476 8888 14504 8919
rect 14292 8860 14504 8888
rect 5644 8792 8432 8820
rect 4065 8783 4123 8789
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 9456 8792 10149 8820
rect 9456 8780 9462 8792
rect 10137 8789 10149 8792
rect 10183 8789 10195 8823
rect 10137 8783 10195 8789
rect 13909 8823 13967 8829
rect 13909 8789 13921 8823
rect 13955 8820 13967 8823
rect 15746 8820 15752 8832
rect 13955 8792 15752 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5445 8619 5503 8625
rect 5445 8585 5457 8619
rect 5491 8616 5503 8619
rect 5718 8616 5724 8628
rect 5491 8588 5724 8616
rect 5491 8585 5503 8588
rect 5445 8579 5503 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6454 8616 6460 8628
rect 5960 8588 6460 8616
rect 5960 8576 5966 8588
rect 6454 8576 6460 8588
rect 6512 8616 6518 8628
rect 7098 8616 7104 8628
rect 6512 8588 7104 8616
rect 6512 8576 6518 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 7248 8588 7297 8616
rect 7248 8576 7254 8588
rect 7285 8585 7297 8588
rect 7331 8585 7343 8619
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 7285 8579 7343 8585
rect 7760 8588 10977 8616
rect 5258 8548 5264 8560
rect 4356 8520 5264 8548
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 1912 8452 2145 8480
rect 1912 8440 1918 8452
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 2133 8443 2191 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3476 8452 3521 8480
rect 3476 8440 3482 8452
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4062 8480 4068 8492
rect 3752 8452 4068 8480
rect 3752 8440 3758 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4356 8489 4384 8520
rect 5258 8508 5264 8520
rect 5316 8548 5322 8560
rect 5810 8548 5816 8560
rect 5316 8520 5816 8548
rect 5316 8508 5322 8520
rect 5810 8508 5816 8520
rect 5868 8508 5874 8560
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4706 8480 4712 8492
rect 4571 8452 4712 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5592 8452 6009 8480
rect 5592 8440 5598 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 7374 8480 7380 8492
rect 5997 8443 6055 8449
rect 6472 8452 7380 8480
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8412 2007 8415
rect 5626 8412 5632 8424
rect 1995 8384 5632 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 6472 8412 6500 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7760 8489 7788 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 15010 8616 15016 8628
rect 13311 8588 15016 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 8297 8551 8355 8557
rect 8297 8517 8309 8551
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8480 7987 8483
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 7975 8452 8217 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 6638 8412 6644 8424
rect 5859 8384 6500 8412
rect 6599 8384 6644 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 7653 8415 7711 8421
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 8312 8412 8340 8511
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 14274 8548 14280 8560
rect 10376 8520 14280 8548
rect 10376 8508 10382 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8480 8999 8483
rect 8987 8452 9444 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 8662 8412 8668 8424
rect 7699 8384 8340 8412
rect 8623 8384 8668 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 9306 8412 9312 8424
rect 8812 8384 9312 8412
rect 8812 8372 8818 8384
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9416 8412 9444 8452
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11425 8483 11483 8489
rect 11425 8480 11437 8483
rect 11204 8452 11437 8480
rect 11204 8440 11210 8452
rect 11425 8449 11437 8452
rect 11471 8449 11483 8483
rect 11425 8443 11483 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 9576 8415 9634 8421
rect 9576 8412 9588 8415
rect 9416 8384 9588 8412
rect 9576 8381 9588 8384
rect 9622 8412 9634 8415
rect 10134 8412 10140 8424
rect 9622 8384 10140 8412
rect 9622 8381 9634 8384
rect 9576 8375 9634 8381
rect 10134 8372 10140 8384
rect 10192 8412 10198 8424
rect 11532 8412 11560 8443
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13688 8452 13737 8480
rect 13688 8440 13694 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 10192 8384 11560 8412
rect 10192 8372 10198 8384
rect 12250 8372 12256 8424
rect 12308 8412 12314 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12308 8384 12817 8412
rect 12308 8372 12314 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 13832 8412 13860 8443
rect 13596 8384 13860 8412
rect 14277 8415 14335 8421
rect 13596 8372 13602 8384
rect 14277 8381 14289 8415
rect 14323 8412 14335 8415
rect 15378 8412 15384 8424
rect 14323 8384 15384 8412
rect 14323 8381 14335 8384
rect 14277 8375 14335 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 3237 8347 3295 8353
rect 3237 8313 3249 8347
rect 3283 8344 3295 8347
rect 3283 8316 3924 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 3896 8285 3924 8316
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4249 8347 4307 8353
rect 4249 8344 4261 8347
rect 4120 8316 4261 8344
rect 4120 8304 4126 8316
rect 4249 8313 4261 8316
rect 4295 8313 4307 8347
rect 4249 8307 4307 8313
rect 4985 8347 5043 8353
rect 4985 8313 4997 8347
rect 5031 8344 5043 8347
rect 6730 8344 6736 8356
rect 5031 8316 6736 8344
rect 5031 8313 5043 8316
rect 4985 8307 5043 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 8205 8347 8263 8353
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8251 8316 10732 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 3881 8279 3939 8285
rect 3881 8245 3893 8279
rect 3927 8245 3939 8279
rect 3881 8239 3939 8245
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 5350 8276 5356 8288
rect 4856 8248 5356 8276
rect 4856 8236 4862 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 6052 8248 6469 8276
rect 6052 8236 6058 8248
rect 6457 8245 6469 8248
rect 6503 8276 6515 8279
rect 6638 8276 6644 8288
rect 6503 8248 6644 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 6638 8236 6644 8248
rect 6696 8276 6702 8288
rect 6822 8276 6828 8288
rect 6696 8248 6828 8276
rect 6696 8236 6702 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 10704 8285 10732 8316
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11606 8344 11612 8356
rect 11204 8316 11612 8344
rect 11204 8304 11210 8316
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 13633 8347 13691 8353
rect 12584 8316 13584 8344
rect 12584 8304 12590 8316
rect 10689 8279 10747 8285
rect 8812 8248 8857 8276
rect 8812 8236 8818 8248
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10962 8276 10968 8288
rect 10735 8248 10968 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12618 8276 12624 8288
rect 12579 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 13556 8276 13584 8316
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 14366 8344 14372 8356
rect 13679 8316 14372 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 14366 8304 14372 8316
rect 14424 8304 14430 8356
rect 14550 8353 14556 8356
rect 14544 8344 14556 8353
rect 14511 8316 14556 8344
rect 14544 8307 14556 8316
rect 14550 8304 14556 8307
rect 14608 8304 14614 8356
rect 17218 8344 17224 8356
rect 14660 8316 17224 8344
rect 14660 8276 14688 8316
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 13556 8248 14688 8276
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 15657 8279 15715 8285
rect 15657 8276 15669 8279
rect 15620 8248 15669 8276
rect 15620 8236 15626 8248
rect 15657 8245 15669 8248
rect 15703 8245 15715 8279
rect 15657 8239 15715 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 5442 8072 5448 8084
rect 3936 8044 5448 8072
rect 3936 8032 3942 8044
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6086 8072 6092 8084
rect 6047 8044 6092 8072
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 6362 8072 6368 8084
rect 6323 8044 6368 8072
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 6730 8072 6736 8084
rect 6691 8044 6736 8072
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7524 8044 7941 8072
rect 7524 8032 7530 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8938 8072 8944 8084
rect 8619 8044 8944 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9677 8075 9735 8081
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 11330 8072 11336 8084
rect 9723 8044 11336 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14424 8044 14565 8072
rect 14424 8032 14430 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 15010 8032 15016 8084
rect 15068 8072 15074 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15068 8044 15669 8072
rect 15068 8032 15074 8044
rect 15657 8041 15669 8044
rect 15703 8041 15715 8075
rect 15657 8035 15715 8041
rect 15746 8032 15752 8084
rect 15804 8072 15810 8084
rect 15804 8044 15849 8072
rect 15804 8032 15810 8044
rect 1765 8007 1823 8013
rect 1765 7973 1777 8007
rect 1811 8004 1823 8007
rect 2038 8004 2044 8016
rect 1811 7976 2044 8004
rect 1811 7973 1823 7976
rect 1765 7967 1823 7973
rect 2038 7964 2044 7976
rect 2096 7964 2102 8016
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2470 8007 2528 8013
rect 2470 8004 2482 8007
rect 2280 7976 2482 8004
rect 2280 7964 2286 7976
rect 2470 7973 2482 7976
rect 2516 7973 2528 8007
rect 2470 7967 2528 7973
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 8021 8007 8079 8013
rect 8021 8004 8033 8007
rect 4120 7976 8033 8004
rect 4120 7964 4126 7976
rect 8021 7973 8033 7976
rect 8067 8004 8079 8007
rect 12618 8004 12624 8016
rect 8067 7976 8984 8004
rect 8067 7973 8079 7976
rect 8021 7967 8079 7973
rect 1486 7936 1492 7948
rect 1447 7908 1492 7936
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 4976 7939 5034 7945
rect 4976 7905 4988 7939
rect 5022 7936 5034 7939
rect 5534 7936 5540 7948
rect 5022 7908 5540 7936
rect 5022 7905 5034 7908
rect 4976 7899 5034 7905
rect 5534 7896 5540 7908
rect 5592 7936 5598 7948
rect 8956 7945 8984 7976
rect 9876 7976 10548 8004
rect 8941 7939 8999 7945
rect 5592 7908 6960 7936
rect 5592 7896 5598 7908
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 6932 7877 6960 7908
rect 8941 7905 8953 7939
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 6917 7831 6975 7837
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3605 7735 3663 7741
rect 3605 7732 3617 7735
rect 2924 7704 3617 7732
rect 2924 7692 2930 7704
rect 3605 7701 3617 7704
rect 3651 7701 3663 7735
rect 3605 7695 3663 7701
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 6840 7732 6868 7831
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 7561 7803 7619 7809
rect 7561 7769 7573 7803
rect 7607 7800 7619 7803
rect 8938 7800 8944 7812
rect 7607 7772 8944 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 8938 7760 8944 7772
rect 8996 7760 9002 7812
rect 5408 7704 6868 7732
rect 5408 7692 5414 7704
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 9048 7732 9076 7831
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 9180 7840 9229 7868
rect 9180 7828 9186 7840
rect 9217 7837 9229 7840
rect 9263 7868 9275 7871
rect 9876 7868 9904 7976
rect 10042 7936 10048 7948
rect 10003 7908 10048 7936
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 10134 7868 10140 7880
rect 9263 7840 9904 7868
rect 10095 7840 10140 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 10244 7800 10272 7831
rect 9732 7772 10272 7800
rect 9732 7760 9738 7772
rect 7708 7704 9076 7732
rect 7708 7692 7714 7704
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10410 7732 10416 7744
rect 9824 7704 10416 7732
rect 9824 7692 9830 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 10520 7732 10548 7976
rect 10980 7976 12624 8004
rect 10980 7945 11008 7976
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 11416 7939 11474 7945
rect 11416 7905 11428 7939
rect 11462 7936 11474 7939
rect 11698 7936 11704 7948
rect 11462 7908 11704 7936
rect 11462 7905 11474 7908
rect 11416 7899 11474 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 13072 7939 13130 7945
rect 13072 7905 13084 7939
rect 13118 7936 13130 7939
rect 13630 7936 13636 7948
rect 13118 7908 13636 7936
rect 13118 7905 13130 7908
rect 13072 7899 13130 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 11146 7868 11152 7880
rect 10796 7840 11152 7868
rect 10796 7809 10824 7840
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 14550 7868 14556 7880
rect 12805 7831 12863 7837
rect 14200 7840 14556 7868
rect 10781 7803 10839 7809
rect 10781 7769 10793 7803
rect 10827 7769 10839 7803
rect 10781 7763 10839 7769
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 10520 7704 12541 7732
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12820 7732 12848 7831
rect 14200 7809 14228 7840
rect 14550 7828 14556 7840
rect 14608 7868 14614 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 14608 7840 15853 7868
rect 14608 7828 14614 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 14185 7803 14243 7809
rect 14185 7769 14197 7803
rect 14231 7769 14243 7803
rect 14185 7763 14243 7769
rect 13538 7732 13544 7744
rect 12820 7704 13544 7732
rect 12529 7695 12587 7701
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15654 7732 15660 7744
rect 15335 7704 15660 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 1964 7500 4016 7528
rect 1964 7404 1992 7500
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3988 7401 4016 7500
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4304 7500 4445 7528
rect 4304 7488 4310 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 5721 7531 5779 7537
rect 5721 7497 5733 7531
rect 5767 7528 5779 7531
rect 5902 7528 5908 7540
rect 5767 7500 5908 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 6236 7500 8217 7528
rect 6236 7488 6242 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7528 8723 7531
rect 8754 7528 8760 7540
rect 8711 7500 8760 7528
rect 8711 7497 8723 7500
rect 8665 7491 8723 7497
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 11054 7528 11060 7540
rect 9723 7500 11060 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 8478 7420 8484 7472
rect 8536 7460 8542 7472
rect 10134 7460 10140 7472
rect 8536 7432 10140 7460
rect 8536 7420 8542 7432
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 14826 7460 14832 7472
rect 13872 7432 14832 7460
rect 13872 7420 13878 7432
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2924 7364 2973 7392
rect 2924 7352 2930 7364
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 4798 7392 4804 7404
rect 4672 7364 4804 7392
rect 4672 7352 4678 7364
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 5000 7324 5028 7355
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 5316 7364 6285 7392
rect 5316 7352 5322 7364
rect 6273 7361 6285 7364
rect 6319 7361 6331 7395
rect 9309 7395 9367 7401
rect 6273 7355 6331 7361
rect 6564 7364 6960 7392
rect 3384 7296 5028 7324
rect 6181 7327 6239 7333
rect 3384 7284 3390 7296
rect 6181 7293 6193 7327
rect 6227 7324 6239 7327
rect 6564 7324 6592 7364
rect 6227 7296 6592 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6832 7327 6890 7333
rect 6832 7324 6844 7327
rect 6788 7296 6844 7324
rect 6788 7284 6794 7296
rect 6832 7293 6844 7296
rect 6878 7293 6890 7327
rect 6932 7324 6960 7364
rect 7852 7364 9260 7392
rect 7852 7324 7880 7364
rect 6932 7296 7880 7324
rect 6832 7287 6890 7293
rect 7300 7268 7328 7296
rect 8846 7284 8852 7336
rect 8904 7324 8910 7336
rect 9122 7324 9128 7336
rect 8904 7296 9128 7324
rect 8904 7284 8910 7296
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9232 7324 9260 7364
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9674 7392 9680 7404
rect 9355 7364 9680 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 10318 7392 10324 7404
rect 10279 7364 10324 7392
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 13688 7364 15025 7392
rect 13688 7352 13694 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 10962 7333 10968 7336
rect 10689 7327 10747 7333
rect 9232 7296 10272 7324
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7256 2927 7259
rect 3602 7256 3608 7268
rect 2915 7228 3608 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 3786 7256 3792 7268
rect 3747 7228 3792 7256
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6454 7256 6460 7268
rect 6135 7228 6460 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 7098 7265 7104 7268
rect 7092 7256 7104 7265
rect 7059 7228 7104 7256
rect 7092 7219 7104 7228
rect 7098 7216 7104 7219
rect 7156 7216 7162 7268
rect 7282 7216 7288 7268
rect 7340 7216 7346 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9048 7228 10149 7256
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 1903 7160 2421 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 2409 7151 2467 7157
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2832 7160 2877 7188
rect 2832 7148 2838 7160
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 3108 7160 3433 7188
rect 3108 7148 3114 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3421 7151 3479 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4798 7188 4804 7200
rect 4759 7160 4804 7188
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 4948 7160 4993 7188
rect 4948 7148 4954 7160
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 9048 7197 9076 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 6328 7160 9045 7188
rect 6328 7148 6334 7160
rect 9033 7157 9045 7160
rect 9079 7157 9091 7191
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 9033 7151 9091 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10244 7188 10272 7296
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10956 7324 10968 7333
rect 10923 7296 10968 7324
rect 10689 7287 10747 7293
rect 10956 7287 10968 7296
rect 10704 7256 10732 7287
rect 10962 7284 10968 7287
rect 11020 7284 11026 7336
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 12676 7296 14013 7324
rect 12676 7284 12682 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14826 7324 14832 7336
rect 14787 7296 14832 7324
rect 14001 7287 14059 7293
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15436 7296 15485 7324
rect 15436 7284 15442 7296
rect 15473 7293 15485 7296
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 15729 7327 15787 7333
rect 15729 7324 15741 7327
rect 15620 7296 15741 7324
rect 15620 7284 15626 7296
rect 15729 7293 15741 7296
rect 15775 7293 15787 7327
rect 15729 7287 15787 7293
rect 11146 7256 11152 7268
rect 10704 7228 11152 7256
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 14844 7256 14872 7284
rect 16666 7256 16672 7268
rect 11256 7228 14780 7256
rect 14844 7228 16672 7256
rect 11256 7188 11284 7228
rect 12066 7188 12072 7200
rect 10244 7160 11284 7188
rect 12027 7160 12072 7188
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13596 7160 13829 7188
rect 13596 7148 13602 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 13817 7151 13875 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14752 7188 14780 7228
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 17678 7256 17684 7268
rect 16776 7228 17684 7256
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14752 7160 14933 7188
rect 14921 7157 14933 7160
rect 14967 7188 14979 7191
rect 16776 7188 16804 7228
rect 17678 7216 17684 7228
rect 17736 7216 17742 7268
rect 14967 7160 16804 7188
rect 16853 7191 16911 7197
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 17034 7188 17040 7200
rect 16899 7160 17040 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 5534 6984 5540 6996
rect 5495 6956 5540 6984
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 6181 6987 6239 6993
rect 6181 6953 6193 6987
rect 6227 6984 6239 6987
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 6227 6956 8493 6984
rect 6227 6953 6239 6956
rect 6181 6947 6239 6953
rect 8481 6953 8493 6956
rect 8527 6953 8539 6987
rect 8481 6947 8539 6953
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10100 6956 10701 6984
rect 10100 6944 10106 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 13446 6984 13452 6996
rect 13407 6956 13452 6984
rect 10689 6947 10747 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 14516 6956 14657 6984
rect 14516 6944 14522 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 14645 6947 14703 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 2222 6876 2228 6928
rect 2280 6916 2286 6928
rect 4706 6916 4712 6928
rect 2280 6888 4712 6916
rect 2280 6876 2286 6888
rect 2308 6851 2366 6857
rect 2308 6817 2320 6851
rect 2354 6848 2366 6851
rect 2866 6848 2872 6860
rect 2354 6820 2872 6848
rect 2354 6817 2366 6820
rect 2308 6811 2366 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4172 6857 4200 6888
rect 4706 6876 4712 6888
rect 4764 6916 4770 6928
rect 6730 6916 6736 6928
rect 4764 6888 6736 6916
rect 4764 6876 4770 6888
rect 6730 6876 6736 6888
rect 6788 6916 6794 6928
rect 6788 6888 6868 6916
rect 6788 6876 6794 6888
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4424 6851 4482 6857
rect 4424 6848 4436 6851
rect 4304 6820 4436 6848
rect 4304 6808 4310 6820
rect 4424 6817 4436 6820
rect 4470 6848 4482 6851
rect 5258 6848 5264 6860
rect 4470 6820 5264 6848
rect 4470 6817 4482 6820
rect 4424 6811 4482 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 6178 6808 6184 6860
rect 6236 6848 6242 6860
rect 6840 6857 6868 6888
rect 9122 6876 9128 6928
rect 9180 6916 9186 6928
rect 11692 6919 11750 6925
rect 9180 6888 10088 6916
rect 9180 6876 9186 6888
rect 6825 6851 6883 6857
rect 6236 6820 6408 6848
rect 6236 6808 6242 6820
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1912 6752 2053 6780
rect 1912 6740 1918 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 2041 6743 2099 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6380 6789 6408 6820
rect 6825 6817 6837 6851
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 7092 6851 7150 6857
rect 7092 6817 7104 6851
rect 7138 6848 7150 6851
rect 8202 6848 8208 6860
rect 7138 6820 8208 6848
rect 7138 6817 7150 6820
rect 7092 6811 7150 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8846 6848 8852 6860
rect 8807 6820 8852 6848
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 10060 6857 10088 6888
rect 11692 6885 11704 6919
rect 11738 6916 11750 6919
rect 12066 6916 12072 6928
rect 11738 6888 12072 6916
rect 11738 6885 11750 6888
rect 11692 6879 11750 6885
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 14553 6919 14611 6925
rect 14553 6916 14565 6919
rect 12584 6888 14565 6916
rect 12584 6876 12590 6888
rect 14553 6885 14565 6888
rect 14599 6885 14611 6919
rect 14553 6879 14611 6885
rect 15488 6888 15976 6916
rect 10045 6851 10103 6857
rect 8996 6820 9041 6848
rect 8996 6808 9002 6820
rect 10045 6817 10057 6851
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 10836 6820 13553 6848
rect 10836 6808 10842 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 15488 6848 15516 6888
rect 13541 6811 13599 6817
rect 13740 6820 15516 6848
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 6365 6743 6423 6749
rect 8220 6752 9045 6780
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 3292 6684 3556 6712
rect 3292 6672 3298 6684
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2004 6616 3433 6644
rect 2004 6604 2010 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3528 6644 3556 6684
rect 5626 6644 5632 6656
rect 3528 6616 5632 6644
rect 3421 6607 3479 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5810 6644 5816 6656
rect 5771 6616 5816 6644
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 8220 6653 8248 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 9033 6743 9091 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6780 10324 6792
rect 10231 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6780 10382 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 10376 6752 11345 6780
rect 10376 6740 10382 6752
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 9306 6712 9312 6724
rect 9180 6684 9312 6712
rect 9180 6672 9186 6684
rect 9306 6672 9312 6684
rect 9364 6712 9370 6724
rect 11146 6712 11152 6724
rect 9364 6684 11152 6712
rect 9364 6672 9370 6684
rect 11146 6672 11152 6684
rect 11204 6712 11210 6724
rect 11440 6712 11468 6743
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12492 6752 13492 6780
rect 12492 6740 12498 6752
rect 11204 6684 11468 6712
rect 11204 6672 11210 6684
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 7248 6616 8217 6644
rect 7248 6604 7254 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 10962 6644 10968 6656
rect 9723 6616 10968 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 12158 6644 12164 6656
rect 11379 6616 12164 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 12158 6604 12164 6616
rect 12216 6644 12222 6656
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12216 6616 12817 6644
rect 12216 6604 12222 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 13081 6647 13139 6653
rect 13081 6613 13093 6647
rect 13127 6644 13139 6647
rect 13354 6644 13360 6656
rect 13127 6616 13360 6644
rect 13127 6613 13139 6616
rect 13081 6607 13139 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13464 6644 13492 6752
rect 13556 6712 13584 6811
rect 13740 6792 13768 6820
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15948 6848 15976 6888
rect 17034 6848 17040 6860
rect 15620 6820 15884 6848
rect 15948 6820 17040 6848
rect 15620 6808 15626 6820
rect 13722 6780 13728 6792
rect 13635 6752 13728 6780
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 15856 6789 15884 6820
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 19150 6857 19156 6860
rect 19144 6848 19156 6857
rect 19111 6820 19156 6848
rect 19144 6811 19156 6820
rect 19150 6808 19156 6811
rect 19208 6808 19214 6860
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14700 6752 14749 6780
rect 14700 6740 14706 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 14737 6743 14795 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 18874 6780 18880 6792
rect 18835 6752 18880 6780
rect 15841 6743 15899 6749
rect 13906 6712 13912 6724
rect 13556 6684 13912 6712
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 14185 6715 14243 6721
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 15764 6712 15792 6743
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 14231 6684 15792 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 14090 6644 14096 6656
rect 13464 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 15194 6644 15200 6656
rect 14516 6616 15200 6644
rect 14516 6604 14522 6616
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15654 6644 15660 6656
rect 15335 6616 15660 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 20254 6644 20260 6656
rect 20215 6616 20260 6644
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 1397 6443 1455 6449
rect 1397 6409 1409 6443
rect 1443 6440 1455 6443
rect 1486 6440 1492 6452
rect 1443 6412 1492 6440
rect 1443 6409 1455 6412
rect 1397 6403 1455 6409
rect 1486 6400 1492 6412
rect 1544 6400 1550 6452
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 1820 6412 2421 6440
rect 1820 6400 1826 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 3878 6440 3884 6452
rect 3839 6412 3884 6440
rect 2409 6403 2467 6409
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 11146 6440 11152 6452
rect 5868 6412 11152 6440
rect 5868 6400 5874 6412
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 15746 6440 15752 6452
rect 14231 6412 15752 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 6822 6372 6828 6384
rect 5031 6344 6828 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 10778 6372 10784 6384
rect 10244 6344 10784 6372
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2924 6276 2973 6304
rect 2924 6264 2930 6276
rect 2961 6273 2973 6276
rect 3007 6304 3019 6307
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 3007 6276 4537 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 4525 6273 4537 6276
rect 4571 6304 4583 6307
rect 4614 6304 4620 6316
rect 4571 6276 4620 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8202 6304 8208 6316
rect 8159 6276 8208 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6304 8539 6307
rect 8846 6304 8852 6316
rect 8527 6276 8852 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 1452 6208 1777 6236
rect 1452 6196 1458 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 3050 6236 3056 6248
rect 1903 6208 3056 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 7466 6236 7472 6248
rect 5684 6208 7472 6236
rect 5684 6196 5690 6208
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7616 6208 7941 6236
rect 7616 6196 7622 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 9122 6236 9128 6248
rect 9083 6208 9128 6236
rect 7929 6199 7987 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10244 6236 10272 6344
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12437 6375 12495 6381
rect 12437 6372 12449 6375
rect 12400 6344 12449 6372
rect 12400 6332 12406 6344
rect 12437 6341 12449 6344
rect 12483 6341 12495 6375
rect 20254 6372 20260 6384
rect 12437 6335 12495 6341
rect 13004 6344 20260 6372
rect 10962 6264 10968 6316
rect 11020 6304 11026 6316
rect 11241 6307 11299 6313
rect 11241 6304 11253 6307
rect 11020 6276 11253 6304
rect 11020 6264 11026 6276
rect 11241 6273 11253 6276
rect 11287 6273 11299 6307
rect 11241 6267 11299 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 9232 6208 10272 6236
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 3421 6171 3479 6177
rect 3421 6168 3433 6171
rect 2823 6140 3433 6168
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 3421 6137 3433 6140
rect 3467 6137 3479 6171
rect 5350 6168 5356 6180
rect 5311 6140 5356 6168
rect 3421 6131 3479 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 9232 6168 9260 6208
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 11112 6208 11161 6236
rect 11112 6196 11118 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 6052 6140 9260 6168
rect 9392 6171 9450 6177
rect 6052 6128 6058 6140
rect 9392 6137 9404 6171
rect 9438 6168 9450 6171
rect 10962 6168 10968 6180
rect 9438 6140 10968 6168
rect 9438 6137 9450 6140
rect 9392 6131 9450 6137
rect 10962 6128 10968 6140
rect 11020 6168 11026 6180
rect 11348 6168 11376 6267
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12032 6276 12909 6304
rect 12032 6264 12038 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 13004 6236 13032 6344
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13722 6304 13728 6316
rect 13127 6276 13728 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14458 6264 14464 6316
rect 14516 6304 14522 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14516 6276 14657 6304
rect 14516 6264 14522 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6304 14887 6307
rect 15102 6304 15108 6316
rect 14875 6276 15108 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15657 6307 15715 6313
rect 15657 6304 15669 6307
rect 15344 6276 15669 6304
rect 15344 6264 15350 6276
rect 15657 6273 15669 6276
rect 15703 6273 15715 6307
rect 15838 6304 15844 6316
rect 15799 6276 15844 6304
rect 15657 6267 15715 6273
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 17126 6304 17132 6316
rect 17087 6276 17132 6304
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 11756 6208 13032 6236
rect 11756 6196 11762 6208
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 17037 6239 17095 6245
rect 17037 6236 17049 6239
rect 13412 6208 17049 6236
rect 13412 6196 13418 6208
rect 17037 6205 17049 6208
rect 17083 6205 17095 6239
rect 17037 6199 17095 6205
rect 18969 6239 19027 6245
rect 18969 6205 18981 6239
rect 19015 6205 19027 6239
rect 18969 6199 19027 6205
rect 18984 6168 19012 6199
rect 11020 6140 11376 6168
rect 11440 6140 19012 6168
rect 19245 6171 19303 6177
rect 11020 6128 11026 6140
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 3510 6100 3516 6112
rect 2915 6072 3516 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3510 6060 3516 6072
rect 3568 6060 3574 6112
rect 4246 6100 4252 6112
rect 4207 6072 4252 6100
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4396 6072 4441 6100
rect 4396 6060 4402 6072
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 5040 6072 5457 6100
rect 5040 6060 5046 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7469 6103 7527 6109
rect 7469 6100 7481 6103
rect 6972 6072 7481 6100
rect 6972 6060 6978 6072
rect 7469 6069 7481 6072
rect 7515 6069 7527 6103
rect 7469 6063 7527 6069
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7708 6072 7849 6100
rect 7708 6060 7714 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 7837 6063 7895 6069
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 9582 6100 9588 6112
rect 8352 6072 9588 6100
rect 8352 6060 8358 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10652 6072 10793 6100
rect 10652 6060 10658 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 11440 6100 11468 6140
rect 19245 6137 19257 6171
rect 19291 6168 19303 6171
rect 19794 6168 19800 6180
rect 19291 6140 19800 6168
rect 19291 6137 19303 6140
rect 19245 6131 19303 6137
rect 19794 6128 19800 6140
rect 19852 6128 19858 6180
rect 11204 6072 11468 6100
rect 11204 6060 11210 6072
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 11664 6072 12817 6100
rect 11664 6060 11670 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14553 6103 14611 6109
rect 14553 6100 14565 6103
rect 14332 6072 14565 6100
rect 14332 6060 14338 6072
rect 14553 6069 14565 6072
rect 14599 6069 14611 6103
rect 15194 6100 15200 6112
rect 15155 6072 15200 6100
rect 14553 6063 14611 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 16577 6103 16635 6109
rect 16577 6069 16589 6103
rect 16623 6100 16635 6103
rect 16758 6100 16764 6112
rect 16623 6072 16764 6100
rect 16623 6069 16635 6072
rect 16577 6063 16635 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 2038 5856 2044 5908
rect 2096 5896 2102 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2096 5868 2789 5896
rect 2096 5856 2102 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 2777 5859 2835 5865
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3844 5868 4077 5896
rect 3844 5856 3850 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4706 5896 4712 5908
rect 4479 5868 4712 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5408 5868 6101 5896
rect 5408 5856 5414 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6328 5868 6561 5896
rect 6328 5856 6334 5868
rect 6549 5865 6561 5868
rect 6595 5865 6607 5899
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6549 5859 6607 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7524 5868 10824 5896
rect 7524 5856 7530 5868
rect 1664 5831 1722 5837
rect 1664 5797 1676 5831
rect 1710 5828 1722 5831
rect 1946 5828 1952 5840
rect 1710 5800 1952 5828
rect 1710 5797 1722 5800
rect 1664 5791 1722 5797
rect 1946 5788 1952 5800
rect 2004 5788 2010 5840
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 6178 5828 6184 5840
rect 4571 5800 6184 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 6178 5788 6184 5800
rect 6236 5828 6242 5840
rect 6236 5800 8064 5828
rect 6236 5788 6242 5800
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 5316 5732 5457 5760
rect 5316 5720 5322 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 6788 5732 7941 5760
rect 6788 5720 6794 5732
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 8036 5760 8064 5800
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 10042 5828 10048 5840
rect 8168 5800 10048 5828
rect 8168 5788 8174 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10796 5828 10824 5868
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 12434 5896 12440 5908
rect 11057 5859 11115 5865
rect 11164 5868 12440 5896
rect 11164 5828 11192 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 13998 5896 14004 5908
rect 12544 5868 14004 5896
rect 10796 5800 11192 5828
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 12544 5828 12572 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 15562 5896 15568 5908
rect 14783 5868 15568 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 20257 5899 20315 5905
rect 20257 5865 20269 5899
rect 20303 5865 20315 5899
rect 20257 5859 20315 5865
rect 11940 5800 12572 5828
rect 11940 5788 11946 5800
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 20272 5828 20300 5859
rect 15988 5800 20300 5828
rect 15988 5788 15994 5800
rect 9766 5760 9772 5772
rect 8036 5732 9772 5760
rect 7929 5723 7987 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 10318 5760 10324 5772
rect 9990 5732 10324 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 13072 5763 13130 5769
rect 11756 5732 11801 5760
rect 11756 5720 11762 5732
rect 13072 5729 13084 5763
rect 13118 5760 13130 5763
rect 15102 5760 15108 5772
rect 13118 5732 15108 5760
rect 13118 5729 13130 5732
rect 13072 5723 13130 5729
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15832 5763 15890 5769
rect 15832 5729 15844 5763
rect 15878 5760 15890 5763
rect 17034 5760 17040 5772
rect 15878 5732 17040 5760
rect 15878 5729 15890 5732
rect 15832 5723 15890 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 17126 5720 17132 5772
rect 17184 5760 17190 5772
rect 17477 5763 17535 5769
rect 17477 5760 17489 5763
rect 17184 5732 17489 5760
rect 17184 5720 17190 5732
rect 17477 5729 17489 5732
rect 17523 5729 17535 5763
rect 17477 5723 17535 5729
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 18785 5763 18843 5769
rect 17920 5732 18552 5760
rect 17920 5720 17926 5732
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5132 5664 5549 5692
rect 5132 5652 5138 5664
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5684 5664 5733 5692
rect 5684 5652 5690 5664
rect 5721 5661 5733 5664
rect 5767 5692 5779 5695
rect 6362 5692 6368 5704
rect 5767 5664 6368 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 7009 5655 7067 5661
rect 4338 5584 4344 5636
rect 4396 5624 4402 5636
rect 7024 5624 7052 5655
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8202 5692 8208 5704
rect 8115 5664 8208 5692
rect 8021 5655 8079 5661
rect 7561 5627 7619 5633
rect 7561 5624 7573 5627
rect 4396 5596 6776 5624
rect 7024 5596 7573 5624
rect 4396 5584 4402 5596
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 6638 5556 6644 5568
rect 5123 5528 6644 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6748 5556 6776 5596
rect 7561 5593 7573 5596
rect 7607 5593 7619 5627
rect 8036 5624 8064 5655
rect 8202 5652 8208 5664
rect 8260 5692 8266 5704
rect 8260 5664 8800 5692
rect 8260 5652 8266 5664
rect 8294 5624 8300 5636
rect 8036 5596 8300 5624
rect 7561 5587 7619 5593
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 7006 5556 7012 5568
rect 6748 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5556 7070 5568
rect 8662 5556 8668 5568
rect 7064 5528 8668 5556
rect 7064 5516 7070 5528
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8772 5556 8800 5664
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9180 5664 9689 5692
rect 9180 5652 9186 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11112 5664 11805 5692
rect 11112 5652 11118 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12158 5692 12164 5704
rect 12023 5664 12164 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12802 5692 12808 5704
rect 12763 5664 12808 5692
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 15436 5664 15577 5692
rect 15436 5652 15442 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 15565 5655 15623 5661
rect 16592 5664 17233 5692
rect 10778 5556 10784 5568
rect 8772 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11204 5528 11345 5556
rect 11204 5516 11210 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 14182 5556 14188 5568
rect 14143 5528 14188 5556
rect 11333 5519 11391 5525
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 15838 5556 15844 5568
rect 15160 5528 15844 5556
rect 15160 5516 15166 5528
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 16592 5556 16620 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 18524 5692 18552 5732
rect 18785 5729 18797 5763
rect 18831 5760 18843 5763
rect 19133 5763 19191 5769
rect 19133 5760 19145 5763
rect 18831 5732 19145 5760
rect 18831 5729 18843 5732
rect 18785 5723 18843 5729
rect 19133 5729 19145 5732
rect 19179 5729 19191 5763
rect 19133 5723 19191 5729
rect 18874 5692 18880 5704
rect 18524 5664 18880 5692
rect 17221 5655 17279 5661
rect 15988 5528 16620 5556
rect 16945 5559 17003 5565
rect 15988 5516 15994 5528
rect 16945 5525 16957 5559
rect 16991 5556 17003 5559
rect 17126 5556 17132 5568
rect 16991 5528 17132 5556
rect 16991 5525 17003 5528
rect 16945 5519 17003 5525
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17236 5556 17264 5655
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 17862 5556 17868 5568
rect 17236 5528 17868 5556
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18601 5559 18659 5565
rect 18601 5556 18613 5559
rect 18012 5528 18613 5556
rect 18012 5516 18018 5528
rect 18601 5525 18613 5528
rect 18647 5556 18659 5559
rect 18785 5559 18843 5565
rect 18785 5556 18797 5559
rect 18647 5528 18797 5556
rect 18647 5525 18659 5528
rect 18601 5519 18659 5525
rect 18785 5525 18797 5528
rect 18831 5525 18843 5559
rect 18785 5519 18843 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 1765 5355 1823 5361
rect 1765 5321 1777 5355
rect 1811 5352 1823 5355
rect 4154 5352 4160 5364
rect 1811 5324 3740 5352
rect 4115 5324 4160 5352
rect 1811 5321 1823 5324
rect 1765 5315 1823 5321
rect 3712 5284 3740 5324
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 10134 5352 10140 5364
rect 5000 5324 10140 5352
rect 4798 5284 4804 5296
rect 3712 5256 4804 5284
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2004 5188 2329 5216
rect 2004 5176 2010 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4706 5216 4712 5228
rect 4212 5188 4712 5216
rect 4212 5176 4218 5188
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 2222 5148 2228 5160
rect 1452 5120 2228 5148
rect 1452 5108 1458 5120
rect 2222 5108 2228 5120
rect 2280 5148 2286 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 2280 5120 2789 5148
rect 2280 5108 2286 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 2777 5111 2835 5117
rect 3044 5151 3102 5157
rect 3044 5117 3056 5151
rect 3090 5148 3102 5151
rect 3326 5148 3332 5160
rect 3090 5120 3332 5148
rect 3090 5117 3102 5120
rect 3044 5111 3102 5117
rect 2792 5080 2820 5111
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 5000 5148 5028 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10042 5244 10048 5296
rect 10100 5284 10106 5296
rect 10686 5284 10692 5296
rect 10100 5256 10692 5284
rect 10100 5244 10106 5256
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 10778 5244 10784 5296
rect 10836 5284 10842 5296
rect 11698 5284 11704 5296
rect 10836 5256 11704 5284
rect 10836 5244 10842 5256
rect 11698 5244 11704 5256
rect 11756 5284 11762 5296
rect 13998 5284 14004 5296
rect 11756 5256 14004 5284
rect 11756 5244 11762 5256
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9232 5188 9873 5216
rect 3936 5120 5028 5148
rect 5077 5151 5135 5157
rect 3936 5108 3942 5120
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5718 5148 5724 5160
rect 5123 5120 5724 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5092 5080 5120 5111
rect 5718 5108 5724 5120
rect 5776 5148 5782 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 5776 5120 7113 5148
rect 5776 5108 5782 5120
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7368 5151 7426 5157
rect 7368 5117 7380 5151
rect 7414 5148 7426 5151
rect 9232 5148 9260 5188
rect 9861 5185 9873 5188
rect 9907 5216 9919 5219
rect 10502 5216 10508 5228
rect 9907 5188 10508 5216
rect 9907 5185 9919 5188
rect 9861 5179 9919 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 7414 5120 9260 5148
rect 9677 5151 9735 5157
rect 7414 5117 7426 5120
rect 7368 5111 7426 5117
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 10594 5148 10600 5160
rect 9723 5120 10600 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 10594 5108 10600 5120
rect 10652 5108 10658 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 11146 5148 11152 5160
rect 10735 5120 11152 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 11992 5148 12020 5179
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12342 5216 12348 5228
rect 12124 5188 12348 5216
rect 12124 5176 12130 5188
rect 12342 5176 12348 5188
rect 12400 5216 12406 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12400 5188 13001 5216
rect 12400 5176 12406 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 12989 5179 13047 5185
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 12158 5148 12164 5160
rect 11992 5120 12164 5148
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 13538 5148 13544 5160
rect 12860 5120 13544 5148
rect 12860 5108 12866 5120
rect 13538 5108 13544 5120
rect 13596 5148 13602 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 13596 5120 14381 5148
rect 13596 5108 13602 5120
rect 14369 5117 14381 5120
rect 14415 5148 14427 5151
rect 15378 5148 15384 5160
rect 14415 5120 15384 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 15378 5108 15384 5120
rect 15436 5148 15442 5160
rect 15930 5148 15936 5160
rect 15436 5120 15936 5148
rect 15436 5108 15442 5120
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17218 5148 17224 5160
rect 16899 5120 17224 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17218 5108 17224 5120
rect 17276 5148 17282 5160
rect 17862 5148 17868 5160
rect 17276 5120 17868 5148
rect 17276 5108 17282 5120
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 2792 5052 5120 5080
rect 5344 5083 5402 5089
rect 5344 5049 5356 5083
rect 5390 5080 5402 5083
rect 6914 5080 6920 5092
rect 5390 5052 6920 5080
rect 5390 5049 5402 5052
rect 5344 5043 5402 5049
rect 6914 5040 6920 5052
rect 6972 5080 6978 5092
rect 6972 5052 8524 5080
rect 6972 5040 6978 5052
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 2280 4984 2325 5012
rect 2280 4972 2286 4984
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 5074 5012 5080 5024
rect 4120 4984 5080 5012
rect 4120 4972 4126 4984
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6420 4984 6469 5012
rect 6420 4972 6426 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7374 5012 7380 5024
rect 6880 4984 7380 5012
rect 6880 4972 6886 4984
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 8496 5021 8524 5052
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 10502 5080 10508 5092
rect 8720 5052 10508 5080
rect 8720 5040 8726 5052
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 12894 5080 12900 5092
rect 12807 5052 12900 5080
rect 12894 5040 12900 5052
rect 12952 5080 12958 5092
rect 13814 5080 13820 5092
rect 12952 5052 13820 5080
rect 12952 5040 12958 5052
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 14636 5083 14694 5089
rect 14636 5049 14648 5083
rect 14682 5080 14694 5083
rect 15010 5080 15016 5092
rect 14682 5052 15016 5080
rect 14682 5049 14694 5052
rect 14636 5043 14694 5049
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 16942 5040 16948 5092
rect 17000 5080 17006 5092
rect 17405 5083 17463 5089
rect 17405 5080 17417 5083
rect 17000 5052 17417 5080
rect 17000 5040 17006 5052
rect 17405 5049 17417 5052
rect 17451 5049 17463 5083
rect 17405 5043 17463 5049
rect 8481 5015 8539 5021
rect 8481 4981 8493 5015
rect 8527 4981 8539 5015
rect 8481 4975 8539 4981
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 5012 9367 5015
rect 9674 5012 9680 5024
rect 9355 4984 9680 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 9815 4984 10333 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10321 4981 10333 4984
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 10827 4984 11345 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 11333 4981 11345 4984
rect 11379 4981 11391 5015
rect 11698 5012 11704 5024
rect 11659 4984 11704 5012
rect 11333 4975 11391 4981
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 11793 5015 11851 5021
rect 11793 4981 11805 5015
rect 11839 5012 11851 5015
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 11839 4984 12449 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 12437 4975 12495 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 13780 4984 15761 5012
rect 13780 4972 13786 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 16390 5012 16396 5024
rect 16351 4984 16396 5012
rect 15749 4975 15807 4981
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 16850 5012 16856 5024
rect 16807 4984 16856 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20622 5012 20628 5024
rect 20027 4984 20628 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 6696 4780 7849 4808
rect 6696 4768 6702 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 10008 4780 10241 4808
rect 10008 4768 10014 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 11054 4808 11060 4820
rect 10827 4780 11060 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11756 4780 11805 4808
rect 11756 4768 11762 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12492 4780 14596 4808
rect 12492 4768 12498 4780
rect 2038 4700 2044 4752
rect 2096 4749 2102 4752
rect 2096 4743 2160 4749
rect 2096 4709 2114 4743
rect 2148 4709 2160 4743
rect 2096 4703 2160 4709
rect 2096 4700 2102 4703
rect 3786 4700 3792 4752
rect 3844 4740 3850 4752
rect 3844 4712 6868 4740
rect 3844 4700 3850 4712
rect 1854 4672 1860 4684
rect 1767 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4672 1918 4684
rect 4332 4675 4390 4681
rect 1912 4644 4108 4672
rect 1912 4632 1918 4644
rect 4080 4616 4108 4644
rect 4332 4641 4344 4675
rect 4378 4672 4390 4675
rect 5626 4672 5632 4684
rect 4378 4644 5632 4672
rect 4378 4641 4390 4644
rect 4332 4635 4390 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6840 4672 6868 4712
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 7432 4712 7757 4740
rect 7432 4700 7438 4712
rect 7745 4709 7757 4712
rect 7791 4709 7803 4743
rect 9398 4740 9404 4752
rect 7745 4703 7803 4709
rect 7852 4712 9404 4740
rect 7852 4672 7880 4712
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 12710 4700 12716 4752
rect 12768 4740 12774 4752
rect 13262 4740 13268 4752
rect 12768 4712 13268 4740
rect 12768 4700 12774 4712
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 13808 4743 13866 4749
rect 13808 4709 13820 4743
rect 13854 4740 13866 4743
rect 14182 4740 14188 4752
rect 13854 4712 14188 4740
rect 13854 4709 13866 4712
rect 13808 4703 13866 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 14568 4740 14596 4780
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15252 4780 15669 4808
rect 15252 4768 15258 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 15804 4780 15849 4808
rect 15804 4768 15810 4780
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 16761 4811 16819 4817
rect 16761 4808 16773 4811
rect 16448 4780 16773 4808
rect 16448 4768 16454 4780
rect 16761 4777 16773 4780
rect 16807 4777 16819 4811
rect 16761 4771 16819 4777
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4777 17371 4811
rect 17313 4771 17371 4777
rect 16669 4743 16727 4749
rect 16669 4740 16681 4743
rect 14568 4712 16681 4740
rect 16669 4709 16681 4712
rect 16715 4709 16727 4743
rect 17328 4740 17356 4771
rect 17328 4712 18368 4740
rect 16669 4703 16727 4709
rect 8754 4672 8760 4684
rect 6840 4644 7880 4672
rect 8715 4644 8760 4672
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 9272 4644 9720 4672
rect 9272 4632 9278 4644
rect 4062 4604 4068 4616
rect 4023 4576 4068 4604
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 6822 4604 6828 4616
rect 5276 4576 6828 4604
rect 3068 4508 4108 4536
rect 198 4428 204 4480
rect 256 4468 262 4480
rect 3068 4468 3096 4508
rect 3234 4468 3240 4480
rect 256 4440 3096 4468
rect 3195 4440 3240 4468
rect 256 4428 262 4440
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4080 4468 4108 4508
rect 5276 4468 5304 4576
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7929 4607 7987 4613
rect 6972 4576 7017 4604
rect 6972 4564 6978 4576
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 8846 4604 8852 4616
rect 8807 4576 8852 4604
rect 7929 4567 7987 4573
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 5445 4539 5503 4545
rect 5445 4536 5457 4539
rect 5408 4508 5457 4536
rect 5408 4496 5414 4508
rect 5445 4505 5457 4508
rect 5491 4536 5503 4539
rect 7944 4536 7972 4567
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9582 4604 9588 4616
rect 9079 4576 9588 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9692 4604 9720 4644
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 10100 4644 10149 4672
rect 10100 4632 10106 4644
rect 10137 4641 10149 4644
rect 10183 4641 10195 4675
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 10137 4635 10195 4641
rect 11146 4632 11152 4644
rect 11204 4672 11210 4684
rect 11606 4672 11612 4684
rect 11204 4644 11612 4672
rect 11204 4632 11210 4644
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 12066 4632 12072 4684
rect 12124 4672 12130 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 12124 4644 12173 4672
rect 12124 4632 12130 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 14200 4672 14228 4700
rect 12308 4644 12353 4672
rect 14200 4644 15884 4672
rect 12308 4632 12314 4644
rect 15856 4616 15884 4644
rect 16758 4632 16764 4684
rect 16816 4672 16822 4684
rect 18340 4681 18368 4712
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 16816 4644 17693 4672
rect 16816 4632 16822 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 17681 4635 17739 4641
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 9692 4576 10333 4604
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11112 4576 11253 4604
rect 11112 4564 11118 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 11425 4567 11483 4573
rect 5491 4508 7972 4536
rect 8389 4539 8447 4545
rect 5491 4505 5503 4508
rect 5445 4499 5503 4505
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 10962 4536 10968 4548
rect 8435 4508 10968 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11440 4536 11468 4567
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 16945 4607 17003 4613
rect 15896 4576 15989 4604
rect 16316 4576 16896 4604
rect 15896 4564 15902 4576
rect 12360 4536 12388 4564
rect 16316 4545 16344 4576
rect 11440 4508 12388 4536
rect 16301 4539 16359 4545
rect 16301 4505 16313 4539
rect 16347 4505 16359 4539
rect 16868 4536 16896 4576
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 17126 4604 17132 4616
rect 16991 4576 17132 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 17126 4564 17132 4576
rect 17184 4564 17190 4616
rect 17773 4607 17831 4613
rect 17773 4573 17785 4607
rect 17819 4573 17831 4607
rect 17954 4604 17960 4616
rect 17915 4576 17960 4604
rect 17773 4567 17831 4573
rect 17788 4536 17816 4567
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 16868 4508 17816 4536
rect 16301 4499 16359 4505
rect 4080 4440 5304 4468
rect 6270 4428 6276 4480
rect 6328 4468 6334 4480
rect 6365 4471 6423 4477
rect 6365 4468 6377 4471
rect 6328 4440 6377 4468
rect 6328 4428 6334 4440
rect 6365 4437 6377 4440
rect 6411 4437 6423 4471
rect 6365 4431 6423 4437
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7377 4471 7435 4477
rect 7377 4468 7389 4471
rect 7248 4440 7389 4468
rect 7248 4428 7254 4440
rect 7377 4437 7389 4440
rect 7423 4437 7435 4471
rect 9766 4468 9772 4480
rect 9727 4440 9772 4468
rect 7377 4431 7435 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 12618 4468 12624 4480
rect 11848 4440 12624 4468
rect 11848 4428 11854 4440
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 14918 4468 14924 4480
rect 14879 4440 14924 4468
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15289 4471 15347 4477
rect 15289 4437 15301 4471
rect 15335 4468 15347 4471
rect 16666 4468 16672 4480
rect 15335 4440 16672 4468
rect 15335 4437 15347 4440
rect 15289 4431 15347 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 2501 4267 2559 4273
rect 2501 4264 2513 4267
rect 2280 4236 2513 4264
rect 2280 4224 2286 4236
rect 2501 4233 2513 4236
rect 2547 4233 2559 4267
rect 8573 4267 8631 4273
rect 2501 4227 2559 4233
rect 5184 4236 7512 4264
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4196 1547 4199
rect 1535 4168 2268 4196
rect 1535 4165 1547 4168
rect 1489 4159 1547 4165
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 2004 4100 2053 4128
rect 2004 4088 2010 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2240 4128 2268 4168
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 2682 4196 2688 4208
rect 2372 4168 2688 4196
rect 2372 4156 2378 4168
rect 2682 4156 2688 4168
rect 2740 4196 2746 4208
rect 3234 4196 3240 4208
rect 2740 4168 3240 4196
rect 2740 4156 2746 4168
rect 3160 4137 3188 4168
rect 3234 4156 3240 4168
rect 3292 4196 3298 4208
rect 3292 4168 4108 4196
rect 3292 4156 3298 4168
rect 3145 4131 3203 4137
rect 2240 4100 3096 4128
rect 2041 4091 2099 4097
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 1820 4032 2881 4060
rect 1820 4020 1826 4032
rect 2869 4029 2881 4032
rect 2915 4060 2927 4063
rect 2958 4060 2964 4072
rect 2915 4032 2964 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3068 4060 3096 4100
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 4080 4128 4108 4168
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4080 4100 4261 4128
rect 3145 4091 3203 4097
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 5184 4128 5212 4236
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 6972 4168 7420 4196
rect 6972 4156 6978 4168
rect 5350 4128 5356 4140
rect 4488 4100 5212 4128
rect 5311 4100 5356 4128
rect 4488 4088 4494 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6362 4128 6368 4140
rect 5684 4100 6368 4128
rect 5684 4088 5690 4100
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7392 4137 7420 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7484 4128 7512 4236
rect 8573 4233 8585 4267
rect 8619 4264 8631 4267
rect 8754 4264 8760 4276
rect 8619 4236 8760 4264
rect 8619 4233 8631 4236
rect 8573 4227 8631 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 12066 4264 12072 4276
rect 8864 4236 12072 4264
rect 7834 4156 7840 4208
rect 7892 4196 7898 4208
rect 8864 4196 8892 4236
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 14976 4236 16896 4264
rect 14976 4224 14982 4236
rect 7892 4168 8892 4196
rect 7892 4156 7898 4168
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 11146 4196 11152 4208
rect 9640 4168 10180 4196
rect 9640 4156 9646 4168
rect 8938 4128 8944 4140
rect 7484 4100 8944 4128
rect 7377 4091 7435 4097
rect 8938 4088 8944 4100
rect 8996 4128 9002 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8996 4100 9045 4128
rect 8996 4088 9002 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9214 4128 9220 4140
rect 9175 4100 9220 4128
rect 9033 4091 9091 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10152 4137 10180 4168
rect 10888 4168 11152 4196
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9824 4100 10057 4128
rect 9824 4088 9830 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10888 4128 10916 4168
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 13722 4196 13728 4208
rect 13096 4168 13728 4196
rect 10459 4100 10916 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 11020 4100 11069 4128
rect 11020 4088 11026 4100
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11238 4128 11244 4140
rect 11199 4100 11244 4128
rect 11057 4091 11115 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 12250 4128 12256 4140
rect 11756 4100 12256 4128
rect 11756 4088 11762 4100
rect 12250 4088 12256 4100
rect 12308 4128 12314 4140
rect 13096 4137 13124 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 15289 4199 15347 4205
rect 15289 4165 15301 4199
rect 15335 4165 15347 4199
rect 15289 4159 15347 4165
rect 13081 4131 13139 4137
rect 12308 4100 13032 4128
rect 12308 4088 12314 4100
rect 4890 4060 4896 4072
rect 3068 4032 4896 4060
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6270 4060 6276 4072
rect 6135 4032 6276 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 7282 4060 7288 4072
rect 7243 4032 7288 4060
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 9732 4032 11621 4060
rect 9732 4020 9738 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 11609 4023 11667 4029
rect 11716 4032 12909 4060
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 8941 3995 8999 4001
rect 1903 3964 3740 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3924 2007 3927
rect 2774 3924 2780 3936
rect 1995 3896 2780 3924
rect 1995 3893 2007 3896
rect 1949 3887 2007 3893
rect 2774 3884 2780 3896
rect 2832 3884 2838 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 3142 3924 3148 3936
rect 3007 3896 3148 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3712 3933 3740 3964
rect 8941 3961 8953 3995
rect 8987 3992 8999 3995
rect 9398 3992 9404 4004
rect 8987 3964 9404 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 9600 3964 10977 3992
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3893 3755 3927
rect 3697 3887 3755 3893
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3844 3896 4077 3924
rect 3844 3884 3850 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4522 3924 4528 3936
rect 4203 3896 4528 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3924 5227 3927
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 5215 3896 5733 3924
rect 5215 3893 5227 3896
rect 5169 3887 5227 3893
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6227 3896 6837 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 9306 3924 9312 3936
rect 7239 3896 9312 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9600 3933 9628 3964
rect 10965 3961 10977 3964
rect 11011 3961 11023 3995
rect 10965 3955 11023 3961
rect 9585 3927 9643 3933
rect 9585 3893 9597 3927
rect 9631 3893 9643 3927
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9585 3887 9643 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10100 3896 10425 3924
rect 10100 3884 10106 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10413 3887 10471 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11716 3924 11744 4032
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 13004 4060 13032 4100
rect 13081 4097 13093 4131
rect 13127 4097 13139 4131
rect 14550 4128 14556 4140
rect 13081 4091 13139 4097
rect 13188 4100 14556 4128
rect 13188 4060 13216 4100
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15102 4128 15108 4140
rect 14967 4100 15108 4128
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 13446 4060 13452 4072
rect 13004 4032 13216 4060
rect 13407 4032 13452 4060
rect 12897 4023 12955 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 15304 4060 15332 4159
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 15896 4168 15976 4196
rect 15896 4156 15902 4168
rect 15948 4137 15976 4168
rect 16868 4137 16896 4236
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 15304 4032 16773 4060
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18506 4060 18512 4072
rect 18095 4032 18512 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 11885 3995 11943 4001
rect 11885 3961 11897 3995
rect 11931 3992 11943 3995
rect 13354 3992 13360 4004
rect 11931 3964 13360 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 13354 3952 13360 3964
rect 13412 3952 13418 4004
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 14292 3964 15761 3992
rect 10836 3896 11744 3924
rect 10836 3884 10842 3896
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12805 3927 12863 3933
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12805 3893 12817 3927
rect 12851 3924 12863 3927
rect 12986 3924 12992 3936
rect 12851 3896 12992 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13633 3927 13691 3933
rect 13633 3893 13645 3927
rect 13679 3924 13691 3927
rect 14090 3924 14096 3936
rect 13679 3896 14096 3924
rect 13679 3893 13691 3896
rect 13633 3887 13691 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14292 3933 14320 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 16666 3992 16672 4004
rect 16627 3964 16672 3992
rect 15749 3955 15807 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 14277 3927 14335 3933
rect 14277 3893 14289 3927
rect 14323 3893 14335 3927
rect 14277 3887 14335 3893
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14608 3896 14657 3924
rect 14608 3884 14614 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 14645 3887 14703 3893
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 15194 3924 15200 3936
rect 14783 3896 15200 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15344 3896 15669 3924
rect 15344 3884 15350 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 15657 3887 15715 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 18782 3924 18788 3936
rect 18279 3896 18788 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3326 3720 3332 3732
rect 3099 3692 3332 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4430 3720 4436 3732
rect 3476 3692 4436 3720
rect 3476 3680 3482 3692
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3720 4767 3723
rect 5074 3720 5080 3732
rect 4755 3692 5080 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 7558 3720 7564 3732
rect 6288 3692 7564 3720
rect 6288 3652 6316 3692
rect 7558 3680 7564 3692
rect 7616 3720 7622 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 7616 3692 8493 3720
rect 7616 3680 7622 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8846 3720 8852 3732
rect 8619 3692 8852 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8846 3680 8852 3692
rect 8904 3680 8910 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9766 3720 9772 3732
rect 9548 3692 9772 3720
rect 9548 3680 9554 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10226 3720 10232 3732
rect 9916 3692 10232 3720
rect 9916 3680 9922 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 10652 3692 13001 3720
rect 10652 3680 10658 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 12989 3683 13047 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 15194 3680 15200 3732
rect 15252 3720 15258 3732
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 15252 3692 15301 3720
rect 15252 3680 15258 3692
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 22462 3720 22468 3732
rect 15289 3683 15347 3689
rect 15396 3692 22468 3720
rect 5092 3624 6316 3652
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1946 3593 1952 3596
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1452 3556 1685 3584
rect 1452 3544 1458 3556
rect 1673 3553 1685 3556
rect 1719 3553 1731 3587
rect 1940 3584 1952 3593
rect 1907 3556 1952 3584
rect 1673 3547 1731 3553
rect 1940 3547 1952 3556
rect 1946 3544 1952 3547
rect 2004 3544 2010 3596
rect 5092 3593 5120 3624
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 7929 3655 7987 3661
rect 7929 3652 7941 3655
rect 6788 3624 7941 3652
rect 6788 3612 6794 3624
rect 7929 3621 7941 3624
rect 7975 3621 7987 3655
rect 9674 3652 9680 3664
rect 7929 3615 7987 3621
rect 8496 3624 9680 3652
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 2976 3556 5089 3584
rect 2976 3528 3004 3556
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 5077 3547 5135 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5994 3593 6000 3596
rect 5988 3547 6000 3593
rect 6052 3584 6058 3596
rect 6052 3556 6088 3584
rect 5994 3544 6000 3547
rect 6052 3544 6058 3556
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 8496 3584 8524 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 11238 3661 11244 3664
rect 11232 3652 11244 3661
rect 9968 3624 11008 3652
rect 11199 3624 11244 3652
rect 6880 3556 8524 3584
rect 8941 3587 8999 3593
rect 6880 3544 6886 3556
rect 8941 3553 8953 3587
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 2958 3476 2964 3528
rect 3016 3476 3022 3528
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 3752 3488 5181 3516
rect 3752 3476 3758 3488
rect 5169 3485 5181 3488
rect 5215 3516 5227 3519
rect 5258 3516 5264 3528
rect 5215 3488 5264 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5626 3516 5632 3528
rect 5399 3488 5632 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7742 3516 7748 3528
rect 6972 3488 7748 3516
rect 6972 3476 6978 3488
rect 7742 3476 7748 3488
rect 7800 3516 7806 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7800 3488 8033 3516
rect 7800 3476 7806 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3516 8539 3519
rect 8956 3516 8984 3547
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 9968 3584 9996 3624
rect 10134 3584 10140 3596
rect 9180 3556 9996 3584
rect 10095 3556 10140 3584
rect 9180 3544 9186 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10980 3593 11008 3624
rect 11232 3615 11244 3624
rect 11238 3612 11244 3615
rect 11296 3612 11302 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 12912 3624 14105 3652
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 8527 3488 8984 3516
rect 9033 3519 9091 3525
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9033 3479 9091 3485
rect 8220 3448 8248 3479
rect 8754 3448 8760 3460
rect 8220 3420 8760 3448
rect 8754 3408 8760 3420
rect 8812 3408 8818 3460
rect 8938 3408 8944 3460
rect 8996 3448 9002 3460
rect 9048 3448 9076 3479
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 10042 3516 10048 3528
rect 9324 3488 10048 3516
rect 9324 3448 9352 3488
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 8996 3420 9352 3448
rect 8996 3408 9002 3420
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 10336 3448 10364 3479
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12912 3516 12940 3624
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 15396 3652 15424 3692
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 14608 3624 15424 3652
rect 14608 3612 14614 3624
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 15657 3655 15715 3661
rect 15657 3652 15669 3655
rect 15528 3624 15669 3652
rect 15528 3612 15534 3624
rect 15657 3621 15669 3624
rect 15703 3652 15715 3655
rect 15703 3624 16528 3652
rect 15703 3621 15715 3624
rect 15657 3615 15715 3621
rect 15102 3584 15108 3596
rect 14292 3556 15108 3584
rect 13078 3516 13084 3528
rect 12124 3488 12940 3516
rect 13039 3488 13084 3516
rect 12124 3476 12130 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14292 3525 14320 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 15804 3556 16313 3584
rect 15804 3544 15810 3556
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 16301 3547 16359 3553
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 15286 3516 15292 3528
rect 14277 3479 14335 3485
rect 14384 3488 15292 3516
rect 9640 3420 10364 3448
rect 12345 3451 12403 3457
rect 9640 3408 9646 3420
rect 12345 3417 12357 3451
rect 12391 3448 12403 3451
rect 12802 3448 12808 3460
rect 12391 3420 12808 3448
rect 12391 3417 12403 3420
rect 12345 3411 12403 3417
rect 12802 3408 12808 3420
rect 12860 3448 12866 3460
rect 13188 3448 13216 3479
rect 12860 3420 13216 3448
rect 13633 3451 13691 3457
rect 12860 3408 12866 3420
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 14384 3448 14412 3488
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 16500 3516 16528 3624
rect 16758 3544 16764 3596
rect 16816 3584 16822 3596
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16816 3556 16865 3584
rect 16816 3544 16822 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 16853 3547 16911 3553
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17405 3587 17463 3593
rect 17405 3584 17417 3587
rect 17000 3556 17417 3584
rect 17000 3544 17006 3556
rect 17405 3553 17417 3556
rect 17451 3553 17463 3587
rect 17405 3547 17463 3553
rect 20254 3516 20260 3528
rect 16500 3488 20260 3516
rect 15841 3479 15899 3485
rect 13679 3420 14412 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 14458 3408 14464 3460
rect 14516 3448 14522 3460
rect 15856 3448 15884 3479
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 14516 3420 15884 3448
rect 17037 3451 17095 3457
rect 14516 3408 14522 3420
rect 17037 3417 17049 3451
rect 17083 3448 17095 3451
rect 21542 3448 21548 3460
rect 17083 3420 21548 3448
rect 17083 3417 17095 3420
rect 17037 3411 17095 3417
rect 21542 3408 21548 3420
rect 21600 3408 21606 3460
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 7374 3380 7380 3392
rect 7147 3352 7380 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 11882 3380 11888 3392
rect 9815 3352 11888 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 15930 3380 15936 3392
rect 12952 3352 15936 3380
rect 12952 3340 12958 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16482 3380 16488 3392
rect 16443 3352 16488 3380
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 17589 3383 17647 3389
rect 17589 3349 17601 3383
rect 17635 3380 17647 3383
rect 22002 3380 22008 3392
rect 17635 3352 22008 3380
rect 17635 3349 17647 3352
rect 17589 3343 17647 3349
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 2004 3148 3433 3176
rect 2004 3136 2010 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 5994 3176 6000 3188
rect 5951 3148 6000 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 8570 3176 8576 3188
rect 6696 3148 8576 3176
rect 6696 3136 6702 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 8720 3148 10180 3176
rect 8720 3136 8726 3148
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6656 3108 6684 3136
rect 8754 3108 8760 3120
rect 5592 3080 6684 3108
rect 8128 3080 8760 3108
rect 5592 3068 5598 3080
rect 4062 3040 4068 3052
rect 3344 3012 4068 3040
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2087 2944 2728 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2314 2913 2320 2916
rect 2308 2904 2320 2913
rect 2275 2876 2320 2904
rect 2308 2867 2320 2876
rect 2314 2864 2320 2867
rect 2372 2864 2378 2916
rect 2700 2904 2728 2944
rect 3344 2904 3372 3012
rect 4062 3000 4068 3012
rect 4120 3040 4126 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4120 3012 4537 3040
rect 4120 3000 4126 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 5776 3012 7113 3040
rect 5776 3000 5782 3012
rect 7101 3009 7113 3012
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 4792 2975 4850 2981
rect 4792 2941 4804 2975
rect 4838 2972 4850 2975
rect 5350 2972 5356 2984
rect 4838 2944 5356 2972
rect 4838 2941 4850 2944
rect 4792 2935 4850 2941
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 7374 2981 7380 2984
rect 7368 2972 7380 2981
rect 7287 2944 7380 2972
rect 7368 2935 7380 2944
rect 7432 2972 7438 2984
rect 8128 2972 8156 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 10152 3108 10180 3148
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10284 3148 10885 3176
rect 10284 3136 10290 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 11054 3176 11060 3188
rect 10873 3139 10931 3145
rect 10980 3148 11060 3176
rect 10597 3111 10655 3117
rect 10152 3080 10548 3108
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 10520 3040 10548 3080
rect 10597 3077 10609 3111
rect 10643 3108 10655 3111
rect 10689 3111 10747 3117
rect 10689 3108 10701 3111
rect 10643 3080 10701 3108
rect 10643 3077 10655 3080
rect 10597 3071 10655 3077
rect 10689 3077 10701 3080
rect 10735 3077 10747 3111
rect 10689 3071 10747 3077
rect 10980 3040 11008 3148
rect 11054 3136 11060 3148
rect 11112 3176 11118 3188
rect 12066 3176 12072 3188
rect 11112 3148 12072 3176
rect 11112 3136 11118 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 19426 3176 19432 3188
rect 12299 3148 19432 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 12526 3108 12532 3120
rect 11532 3080 12532 3108
rect 8260 3012 9352 3040
rect 10520 3012 11008 3040
rect 8260 3000 8266 3012
rect 8662 2972 8668 2984
rect 7432 2944 8156 2972
rect 8220 2944 8668 2972
rect 7374 2932 7380 2935
rect 7432 2932 7438 2944
rect 2700 2876 3372 2904
rect 3436 2876 3832 2904
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 3436 2836 3464 2876
rect 1636 2808 3464 2836
rect 1636 2796 1642 2808
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3697 2839 3755 2845
rect 3697 2836 3709 2839
rect 3568 2808 3709 2836
rect 3568 2796 3574 2808
rect 3697 2805 3709 2808
rect 3743 2805 3755 2839
rect 3804 2836 3832 2876
rect 5258 2864 5264 2916
rect 5316 2904 5322 2916
rect 8110 2904 8116 2916
rect 5316 2876 8116 2904
rect 5316 2864 5322 2876
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 8220 2836 8248 2944
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9180 2944 9229 2972
rect 9180 2932 9186 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9324 2972 9352 3012
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 11112 3012 11437 3040
rect 11112 3000 11118 3012
rect 11425 3009 11437 3012
rect 11471 3009 11483 3043
rect 11425 3003 11483 3009
rect 11532 2972 11560 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 15562 3068 15568 3120
rect 15620 3108 15626 3120
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 15620 3080 16773 3108
rect 15620 3068 15626 3080
rect 16761 3077 16773 3080
rect 16807 3077 16819 3111
rect 16761 3071 16819 3077
rect 15212 3012 18920 3040
rect 12802 2981 12808 2984
rect 9324 2944 11560 2972
rect 12529 2975 12587 2981
rect 9217 2935 9275 2941
rect 12529 2941 12541 2975
rect 12575 2941 12587 2975
rect 12796 2972 12808 2981
rect 12763 2944 12808 2972
rect 12529 2935 12587 2941
rect 12796 2935 12808 2944
rect 9462 2907 9520 2913
rect 9462 2904 9474 2907
rect 8496 2876 9474 2904
rect 3804 2808 8248 2836
rect 3697 2799 3755 2805
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8496 2845 8524 2876
rect 9462 2873 9474 2876
rect 9508 2904 9520 2907
rect 9582 2904 9588 2916
rect 9508 2876 9588 2904
rect 9508 2873 9520 2876
rect 9462 2867 9520 2873
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 10689 2907 10747 2913
rect 10689 2873 10701 2907
rect 10735 2904 10747 2907
rect 11146 2904 11152 2916
rect 10735 2876 11152 2904
rect 10735 2873 10747 2876
rect 10689 2867 10747 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 11241 2907 11299 2913
rect 11241 2873 11253 2907
rect 11287 2904 11299 2907
rect 11974 2904 11980 2916
rect 11287 2876 11980 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 11974 2864 11980 2876
rect 12032 2904 12038 2916
rect 12253 2907 12311 2913
rect 12253 2904 12265 2907
rect 12032 2876 12265 2904
rect 12032 2864 12038 2876
rect 12253 2873 12265 2876
rect 12299 2873 12311 2907
rect 12544 2904 12572 2935
rect 12802 2932 12808 2935
rect 12860 2932 12866 2984
rect 13538 2972 13544 2984
rect 12912 2944 13544 2972
rect 12912 2904 12940 2944
rect 13538 2932 13544 2944
rect 13596 2972 13602 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13596 2944 14197 2972
rect 13596 2932 13602 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 15212 2972 15240 3012
rect 14185 2935 14243 2941
rect 14292 2944 15240 2972
rect 14292 2904 14320 2944
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15712 2944 15853 2972
rect 15712 2932 15718 2944
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16577 2975 16635 2981
rect 16577 2972 16589 2975
rect 15988 2944 16589 2972
rect 15988 2932 15994 2944
rect 16577 2941 16589 2944
rect 16623 2941 16635 2975
rect 16577 2935 16635 2941
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 14458 2913 14464 2916
rect 14452 2904 14464 2913
rect 12544 2876 12940 2904
rect 13004 2876 14320 2904
rect 14384 2876 14464 2904
rect 12253 2867 12311 2873
rect 8481 2839 8539 2845
rect 8481 2836 8493 2839
rect 8352 2808 8493 2836
rect 8352 2796 8358 2808
rect 8481 2805 8493 2808
rect 8527 2805 8539 2839
rect 8481 2799 8539 2805
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9214 2836 9220 2848
rect 8812 2808 9220 2836
rect 8812 2796 8818 2808
rect 9214 2796 9220 2808
rect 9272 2836 9278 2848
rect 11054 2836 11060 2848
rect 9272 2808 11060 2836
rect 9272 2796 9278 2808
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11330 2836 11336 2848
rect 11291 2808 11336 2836
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 13004 2836 13032 2876
rect 12492 2808 13032 2836
rect 13909 2839 13967 2845
rect 12492 2796 12498 2808
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 14384 2836 14412 2876
rect 14452 2867 14464 2876
rect 14458 2864 14464 2867
rect 14516 2864 14522 2916
rect 15010 2864 15016 2916
rect 15068 2904 15074 2916
rect 16117 2907 16175 2913
rect 15068 2876 15700 2904
rect 15068 2864 15074 2876
rect 13955 2808 14412 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 15565 2839 15623 2845
rect 15565 2836 15577 2839
rect 15160 2808 15577 2836
rect 15160 2796 15166 2808
rect 15565 2805 15577 2808
rect 15611 2805 15623 2839
rect 15672 2836 15700 2876
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 17144 2904 17172 2935
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 18892 2981 18920 3012
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17368 2944 18061 2972
rect 17368 2932 17374 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 16163 2876 17172 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 16666 2836 16672 2848
rect 15672 2808 16672 2836
rect 15565 2799 15623 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 17313 2839 17371 2845
rect 17313 2836 17325 2839
rect 17000 2808 17325 2836
rect 17000 2796 17006 2808
rect 17313 2805 17325 2808
rect 17359 2805 17371 2839
rect 17313 2799 17371 2805
rect 18233 2839 18291 2845
rect 18233 2805 18245 2839
rect 18279 2836 18291 2839
rect 18506 2836 18512 2848
rect 18279 2808 18512 2836
rect 18279 2805 18291 2808
rect 18233 2799 18291 2805
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 19061 2839 19119 2845
rect 19061 2805 19073 2839
rect 19107 2836 19119 2839
rect 19702 2836 19708 2848
rect 19107 2808 19708 2836
rect 19107 2805 19119 2808
rect 19061 2799 19119 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2130 2632 2136 2644
rect 1995 2604 2136 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3421 2635 3479 2641
rect 2363 2604 3280 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 3142 2564 3148 2576
rect 2455 2536 3148 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 3252 2564 3280 2604
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 3970 2632 3976 2644
rect 3467 2604 3976 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 4764 2604 5457 2632
rect 4764 2592 4770 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7558 2632 7564 2644
rect 7423 2604 7564 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7929 2635 7987 2641
rect 7929 2601 7941 2635
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 3510 2564 3516 2576
rect 3252 2536 3516 2564
rect 3510 2524 3516 2536
rect 3568 2524 3574 2576
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 7190 2564 7196 2576
rect 5399 2536 7196 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 7944 2564 7972 2595
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 8297 2635 8355 2641
rect 8297 2632 8309 2635
rect 8260 2604 8309 2632
rect 8260 2592 8266 2604
rect 8297 2601 8309 2604
rect 8343 2601 8355 2635
rect 8297 2595 8355 2601
rect 9861 2635 9919 2641
rect 9861 2601 9873 2635
rect 9907 2632 9919 2635
rect 9950 2632 9956 2644
rect 9907 2604 9956 2632
rect 9907 2601 9919 2604
rect 9861 2595 9919 2601
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10192 2604 10425 2632
rect 10192 2592 10198 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 10873 2635 10931 2641
rect 10873 2601 10885 2635
rect 10919 2632 10931 2635
rect 11698 2632 11704 2644
rect 10919 2604 11704 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 14550 2592 14556 2644
rect 14608 2632 14614 2644
rect 16209 2635 16267 2641
rect 16209 2632 16221 2635
rect 14608 2604 16221 2632
rect 14608 2592 14614 2604
rect 16209 2601 16221 2604
rect 16255 2601 16267 2635
rect 16209 2595 16267 2601
rect 16666 2592 16672 2644
rect 16724 2632 16730 2644
rect 16761 2635 16819 2641
rect 16761 2632 16773 2635
rect 16724 2604 16773 2632
rect 16724 2592 16730 2604
rect 16761 2601 16773 2604
rect 16807 2601 16819 2635
rect 16761 2595 16819 2601
rect 7331 2536 7972 2564
rect 8312 2536 9628 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 2682 2496 2688 2508
rect 2608 2468 2688 2496
rect 2608 2437 2636 2468
rect 2682 2456 2688 2468
rect 2740 2496 2746 2508
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2740 2468 2789 2496
rect 2740 2456 2746 2468
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 3329 2499 3387 2505
rect 3329 2465 3341 2499
rect 3375 2496 3387 2499
rect 5258 2496 5264 2508
rect 3375 2468 5264 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2496 6331 2499
rect 8312 2496 8340 2536
rect 6319 2468 8340 2496
rect 8389 2499 8447 2505
rect 6319 2465 6331 2468
rect 6273 2459 6331 2465
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8662 2496 8668 2508
rect 8435 2468 8668 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2915 2400 3525 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5902 2428 5908 2440
rect 5675 2400 5908 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 2961 2363 3019 2369
rect 2961 2360 2973 2363
rect 2832 2332 2973 2360
rect 2832 2320 2838 2332
rect 2961 2329 2973 2332
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 6012 2360 6040 2459
rect 8662 2456 8668 2468
rect 8720 2456 8726 2508
rect 9600 2496 9628 2536
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10778 2564 10784 2576
rect 9732 2536 10784 2564
rect 9732 2524 9738 2536
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 12897 2567 12955 2573
rect 11716 2536 12112 2564
rect 11716 2496 11744 2536
rect 9600 2468 11744 2496
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 11882 2496 11888 2508
rect 11839 2468 11888 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 8294 2428 8300 2440
rect 7607 2400 8300 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9214 2428 9220 2440
rect 8619 2400 9220 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11054 2428 11060 2440
rect 11011 2400 11060 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11204 2400 11989 2428
rect 11204 2388 11210 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 12084 2428 12112 2536
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 13446 2564 13452 2576
rect 12943 2536 13452 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 13446 2524 13452 2536
rect 13504 2524 13510 2576
rect 16298 2564 16304 2576
rect 14292 2536 16304 2564
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13354 2496 13360 2508
rect 13315 2468 13360 2496
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 14292 2505 14320 2536
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 14277 2459 14335 2465
rect 14384 2468 15485 2496
rect 14384 2428 14412 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15887 2468 16037 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 16577 2499 16635 2505
rect 16577 2465 16589 2499
rect 16623 2465 16635 2499
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 16577 2459 16635 2465
rect 12084 2400 14412 2428
rect 14553 2431 14611 2437
rect 11977 2391 12035 2397
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 16592 2428 16620 2459
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 17678 2496 17684 2508
rect 17639 2468 17684 2496
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18012 2468 18337 2496
rect 18012 2456 18018 2468
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 18325 2459 18383 2465
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 20254 2496 20260 2508
rect 20215 2468 20260 2496
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 14599 2400 16620 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 5031 2332 6040 2360
rect 11425 2363 11483 2369
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 11425 2329 11437 2363
rect 11471 2360 11483 2363
rect 13078 2360 13084 2372
rect 11471 2332 13084 2360
rect 11471 2329 11483 2332
rect 11425 2323 11483 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 15841 2363 15899 2369
rect 15841 2360 15853 2363
rect 13872 2332 15853 2360
rect 13872 2320 13878 2332
rect 15841 2329 15853 2332
rect 15887 2329 15899 2363
rect 15841 2323 15899 2329
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 17313 2363 17371 2369
rect 17313 2360 17325 2363
rect 16080 2332 17325 2360
rect 16080 2320 16086 2332
rect 17313 2329 17325 2332
rect 17359 2329 17371 2363
rect 17313 2323 17371 2329
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 11882 2292 11888 2304
rect 6963 2264 11888 2292
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13228 2264 13553 2292
rect 13228 2252 13234 2264
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 13630 2252 13636 2304
rect 13688 2292 13694 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 13688 2264 15669 2292
rect 13688 2252 13694 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17460 2264 17877 2292
rect 17460 2252 17466 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 18012 2264 18521 2292
rect 18012 2252 18018 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 19061 2295 19119 2301
rect 19061 2261 19073 2295
rect 19107 2292 19119 2295
rect 19242 2292 19248 2304
rect 19107 2264 19248 2292
rect 19107 2261 19119 2264
rect 19061 2255 19119 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2292 19671 2295
rect 20162 2292 20168 2304
rect 19659 2264 20168 2292
rect 19659 2261 19671 2264
rect 19613 2255 19671 2261
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 20441 2295 20499 2301
rect 20441 2261 20453 2295
rect 20487 2292 20499 2295
rect 21082 2292 21088 2304
rect 20487 2264 21088 2292
rect 20487 2261 20499 2264
rect 20441 2255 20499 2261
rect 21082 2252 21088 2264
rect 21140 2252 21146 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 658 2048 664 2100
rect 716 2088 722 2100
rect 6914 2088 6920 2100
rect 716 2060 6920 2088
rect 716 2048 722 2060
rect 6914 2048 6920 2060
rect 6972 2048 6978 2100
rect 2038 1980 2044 2032
rect 2096 2020 2102 2032
rect 3694 2020 3700 2032
rect 2096 1992 3700 2020
rect 2096 1980 2102 1992
rect 3694 1980 3700 1992
rect 3752 1980 3758 2032
rect 2498 1912 2504 1964
rect 2556 1952 2562 1964
rect 8938 1952 8944 1964
rect 2556 1924 8944 1952
rect 2556 1912 2562 1924
rect 8938 1912 8944 1924
rect 8996 1912 9002 1964
rect 1118 1844 1124 1896
rect 1176 1884 1182 1896
rect 6730 1884 6736 1896
rect 1176 1856 6736 1884
rect 1176 1844 1182 1856
rect 6730 1844 6736 1856
rect 6788 1844 6794 1896
<< via1 >>
rect 4252 21904 4304 21956
rect 4620 21904 4672 21956
rect 6092 21904 6144 21956
rect 6276 21904 6328 21956
rect 7104 20272 7156 20324
rect 7932 20272 7984 20324
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 3608 20043 3660 20052
rect 3608 20009 3617 20043
rect 3617 20009 3651 20043
rect 3651 20009 3660 20043
rect 3608 20000 3660 20009
rect 12900 20000 12952 20052
rect 19340 20000 19392 20052
rect 20260 20000 20312 20052
rect 4988 19932 5040 19984
rect 13268 19932 13320 19984
rect 2688 19864 2740 19916
rect 5908 19907 5960 19916
rect 2044 19796 2096 19848
rect 5908 19873 5917 19907
rect 5917 19873 5951 19907
rect 5951 19873 5960 19907
rect 5908 19864 5960 19873
rect 7748 19907 7800 19916
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 13636 19864 13688 19916
rect 18604 19864 18656 19916
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 6920 19796 6972 19848
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 8208 19796 8260 19848
rect 9864 19796 9916 19848
rect 9036 19728 9088 19780
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 5632 19660 5684 19712
rect 6368 19660 6420 19712
rect 6828 19660 6880 19712
rect 8852 19660 8904 19712
rect 16672 19660 16724 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3332 19499 3384 19508
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 7840 19499 7892 19508
rect 2872 19388 2924 19440
rect 2688 19363 2740 19372
rect 2688 19329 2697 19363
rect 2697 19329 2731 19363
rect 2731 19329 2740 19363
rect 2688 19320 2740 19329
rect 2044 19252 2096 19304
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 2872 19116 2924 19168
rect 3792 19184 3844 19236
rect 4804 19252 4856 19304
rect 4988 19252 5040 19304
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 6092 19388 6144 19440
rect 6276 19388 6328 19440
rect 6828 19295 6880 19304
rect 4160 19159 4212 19168
rect 4160 19125 4169 19159
rect 4169 19125 4203 19159
rect 4203 19125 4212 19159
rect 4160 19116 4212 19125
rect 5448 19184 5500 19236
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 9036 19363 9088 19372
rect 7656 19252 7708 19304
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 8852 19295 8904 19304
rect 8484 19184 8536 19236
rect 8852 19261 8861 19295
rect 8861 19261 8895 19295
rect 8895 19261 8904 19295
rect 8852 19252 8904 19261
rect 9496 19252 9548 19304
rect 12164 19320 12216 19372
rect 9864 19227 9916 19236
rect 9864 19193 9898 19227
rect 9898 19193 9916 19227
rect 9864 19184 9916 19193
rect 12624 19252 12676 19304
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 7564 19116 7616 19168
rect 11888 19184 11940 19236
rect 11980 19184 12032 19236
rect 12808 19184 12860 19236
rect 14096 19252 14148 19304
rect 14464 19252 14516 19304
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 15476 19252 15528 19304
rect 16212 19295 16264 19304
rect 16212 19261 16221 19295
rect 16221 19261 16255 19295
rect 16255 19261 16264 19295
rect 16212 19252 16264 19261
rect 16948 19252 17000 19304
rect 12440 19116 12492 19168
rect 13360 19116 13412 19168
rect 14280 19116 14332 19168
rect 15200 19116 15252 19168
rect 15660 19116 15712 19168
rect 16120 19116 16172 19168
rect 17040 19184 17092 19236
rect 17224 19252 17276 19304
rect 17500 19252 17552 19304
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 22100 19184 22152 19236
rect 17408 19116 17460 19168
rect 17960 19116 18012 19168
rect 18512 19116 18564 19168
rect 20720 19116 20772 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 3148 18844 3200 18896
rect 1952 18776 2004 18828
rect 1676 18683 1728 18692
rect 1676 18649 1685 18683
rect 1685 18649 1719 18683
rect 1719 18649 1728 18683
rect 1676 18640 1728 18649
rect 2780 18776 2832 18828
rect 3884 18776 3936 18828
rect 3700 18708 3752 18760
rect 5540 18844 5592 18896
rect 5908 18912 5960 18964
rect 7748 18912 7800 18964
rect 8484 18912 8536 18964
rect 9680 18912 9732 18964
rect 9864 18912 9916 18964
rect 7012 18844 7064 18896
rect 7656 18887 7708 18896
rect 7656 18853 7690 18887
rect 7690 18853 7708 18887
rect 7656 18844 7708 18853
rect 8024 18844 8076 18896
rect 9496 18844 9548 18896
rect 12624 18912 12676 18964
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 14556 18912 14608 18964
rect 16580 18912 16632 18964
rect 18880 18912 18932 18964
rect 19800 18912 19852 18964
rect 6920 18776 6972 18828
rect 12532 18844 12584 18896
rect 12716 18844 12768 18896
rect 14004 18844 14056 18896
rect 14188 18844 14240 18896
rect 15108 18844 15160 18896
rect 16672 18844 16724 18896
rect 21640 18844 21692 18896
rect 4344 18708 4396 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 4252 18683 4304 18692
rect 4252 18649 4261 18683
rect 4261 18649 4295 18683
rect 4295 18649 4304 18683
rect 4252 18640 4304 18649
rect 10324 18776 10376 18828
rect 12348 18776 12400 18828
rect 13452 18776 13504 18828
rect 13636 18819 13688 18828
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 9128 18751 9180 18760
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 3240 18572 3292 18624
rect 5816 18572 5868 18624
rect 7288 18572 7340 18624
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 9496 18708 9548 18760
rect 12808 18708 12860 18760
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 16396 18776 16448 18828
rect 18972 18819 19024 18828
rect 18972 18785 18981 18819
rect 18981 18785 19015 18819
rect 19015 18785 19024 18819
rect 18972 18776 19024 18785
rect 16304 18708 16356 18760
rect 8024 18572 8076 18624
rect 8116 18572 8168 18624
rect 10324 18572 10376 18624
rect 15936 18640 15988 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1492 18368 1544 18420
rect 2504 18368 2556 18420
rect 1952 18164 2004 18216
rect 3700 18368 3752 18420
rect 6000 18368 6052 18420
rect 10140 18368 10192 18420
rect 13820 18368 13872 18420
rect 15292 18368 15344 18420
rect 22560 18368 22612 18420
rect 7288 18300 7340 18352
rect 6828 18232 6880 18284
rect 8576 18300 8628 18352
rect 10048 18300 10100 18352
rect 10600 18300 10652 18352
rect 12164 18300 12216 18352
rect 21180 18300 21232 18352
rect 8484 18232 8536 18284
rect 10324 18275 10376 18284
rect 4252 18164 4304 18216
rect 4712 18164 4764 18216
rect 7288 18164 7340 18216
rect 8116 18164 8168 18216
rect 9128 18164 9180 18216
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 12532 18232 12584 18284
rect 16028 18232 16080 18284
rect 17500 18232 17552 18284
rect 19340 18232 19392 18284
rect 12256 18164 12308 18216
rect 12900 18164 12952 18216
rect 15016 18207 15068 18216
rect 3792 18139 3844 18148
rect 3792 18105 3826 18139
rect 3826 18105 3844 18139
rect 3792 18096 3844 18105
rect 10692 18096 10744 18148
rect 11612 18096 11664 18148
rect 13084 18096 13136 18148
rect 15016 18173 15025 18207
rect 15025 18173 15059 18207
rect 15059 18173 15068 18207
rect 15016 18164 15068 18173
rect 18420 18207 18472 18216
rect 13820 18096 13872 18148
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 16856 18096 16908 18148
rect 3056 18028 3108 18080
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 4804 18028 4856 18080
rect 6828 18028 6880 18080
rect 9312 18028 9364 18080
rect 9956 18028 10008 18080
rect 10324 18028 10376 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 12808 18028 12860 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 2872 17867 2924 17876
rect 2872 17833 2881 17867
rect 2881 17833 2915 17867
rect 2915 17833 2924 17867
rect 2872 17824 2924 17833
rect 2964 17824 3016 17876
rect 4160 17824 4212 17876
rect 6920 17824 6972 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 12532 17867 12584 17876
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 12808 17867 12860 17876
rect 12808 17833 12817 17867
rect 12817 17833 12851 17867
rect 12851 17833 12860 17867
rect 12808 17824 12860 17833
rect 13820 17867 13872 17876
rect 13820 17833 13829 17867
rect 13829 17833 13863 17867
rect 13863 17833 13872 17867
rect 13820 17824 13872 17833
rect 2780 17756 2832 17808
rect 3056 17756 3108 17808
rect 5448 17756 5500 17808
rect 6828 17799 6880 17808
rect 6828 17765 6862 17799
rect 6862 17765 6880 17799
rect 6828 17756 6880 17765
rect 1768 17688 1820 17740
rect 1860 17688 1912 17740
rect 3148 17688 3200 17740
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 8760 17756 8812 17808
rect 10048 17799 10100 17808
rect 10048 17765 10057 17799
rect 10057 17765 10091 17799
rect 10091 17765 10100 17799
rect 10048 17756 10100 17765
rect 11796 17756 11848 17808
rect 13084 17756 13136 17808
rect 13636 17756 13688 17808
rect 3240 17620 3292 17672
rect 1032 17552 1084 17604
rect 5264 17620 5316 17672
rect 3608 17552 3660 17604
rect 7288 17688 7340 17740
rect 10784 17688 10836 17740
rect 5816 17620 5868 17672
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 12900 17688 12952 17740
rect 16120 17688 16172 17740
rect 14280 17663 14332 17672
rect 3884 17484 3936 17536
rect 7748 17484 7800 17536
rect 8208 17527 8260 17536
rect 8208 17493 8217 17527
rect 8217 17493 8251 17527
rect 8251 17493 8260 17527
rect 8208 17484 8260 17493
rect 9680 17484 9732 17536
rect 10784 17484 10836 17536
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 12348 17484 12400 17536
rect 12716 17484 12768 17536
rect 16396 17484 16448 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1860 17323 1912 17332
rect 1860 17289 1869 17323
rect 1869 17289 1903 17323
rect 1903 17289 1912 17323
rect 1860 17280 1912 17289
rect 8208 17280 8260 17332
rect 8576 17280 8628 17332
rect 6184 17212 6236 17264
rect 8760 17212 8812 17264
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 3976 17144 4028 17196
rect 4252 17144 4304 17196
rect 7104 17144 7156 17196
rect 7380 17144 7432 17196
rect 8576 17144 8628 17196
rect 11796 17280 11848 17332
rect 15108 17280 15160 17332
rect 12992 17187 13044 17196
rect 1952 17076 2004 17128
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 2964 17076 3016 17128
rect 3240 17008 3292 17060
rect 9496 17076 9548 17128
rect 4712 17008 4764 17060
rect 6920 17008 6972 17060
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 11796 17076 11848 17128
rect 13912 17076 13964 17128
rect 14372 17119 14424 17128
rect 14372 17085 14406 17119
rect 14406 17085 14424 17119
rect 14372 17076 14424 17085
rect 4252 16983 4304 16992
rect 4252 16949 4261 16983
rect 4261 16949 4295 16983
rect 4295 16949 4304 16983
rect 4252 16940 4304 16949
rect 5908 16940 5960 16992
rect 6000 16940 6052 16992
rect 7656 16940 7708 16992
rect 8852 16940 8904 16992
rect 11060 17008 11112 17060
rect 12348 17008 12400 17060
rect 13728 17008 13780 17060
rect 17960 17008 18012 17060
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 10508 16940 10560 16992
rect 11704 16940 11756 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 15844 16940 15896 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1492 16736 1544 16788
rect 2504 16736 2556 16788
rect 2964 16736 3016 16788
rect 1768 16668 1820 16720
rect 3240 16668 3292 16720
rect 3884 16668 3936 16720
rect 4252 16668 4304 16720
rect 4712 16736 4764 16788
rect 5908 16736 5960 16788
rect 6000 16668 6052 16720
rect 6184 16711 6236 16720
rect 6184 16677 6218 16711
rect 6218 16677 6236 16711
rect 6184 16668 6236 16677
rect 7656 16736 7708 16788
rect 7748 16736 7800 16788
rect 9312 16736 9364 16788
rect 11060 16779 11112 16788
rect 3332 16643 3384 16652
rect 3332 16609 3341 16643
rect 3341 16609 3375 16643
rect 3375 16609 3384 16643
rect 3332 16600 3384 16609
rect 2136 16532 2188 16584
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 4712 16600 4764 16652
rect 4896 16600 4948 16652
rect 2872 16464 2924 16516
rect 3976 16464 4028 16516
rect 2780 16396 2832 16448
rect 5816 16532 5868 16584
rect 8484 16600 8536 16652
rect 9680 16668 9732 16720
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11152 16736 11204 16788
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 13728 16668 13780 16720
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 10232 16600 10284 16652
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 13820 16600 13872 16652
rect 11888 16575 11940 16584
rect 8760 16464 8812 16516
rect 9496 16464 9548 16516
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 14372 16736 14424 16788
rect 5264 16396 5316 16448
rect 11704 16464 11756 16516
rect 11060 16396 11112 16448
rect 15568 16532 15620 16584
rect 13728 16396 13780 16448
rect 17408 16396 17460 16448
rect 20352 16396 20404 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1584 16192 1636 16244
rect 3424 16192 3476 16244
rect 6920 16192 6972 16244
rect 8576 16235 8628 16244
rect 8576 16201 8585 16235
rect 8585 16201 8619 16235
rect 8619 16201 8628 16235
rect 8576 16192 8628 16201
rect 10508 16235 10560 16244
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 14280 16192 14332 16244
rect 16120 16235 16172 16244
rect 16120 16201 16129 16235
rect 16129 16201 16163 16235
rect 16163 16201 16172 16235
rect 16120 16192 16172 16201
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 5724 16124 5776 16176
rect 2136 16056 2188 16108
rect 3148 16056 3200 16108
rect 3332 16056 3384 16108
rect 4252 16056 4304 16108
rect 5540 16056 5592 16108
rect 10232 16167 10284 16176
rect 10232 16133 10241 16167
rect 10241 16133 10275 16167
rect 10275 16133 10284 16167
rect 10232 16124 10284 16133
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 5172 15988 5224 16040
rect 8300 15988 8352 16040
rect 8760 15988 8812 16040
rect 4896 15920 4948 15972
rect 4988 15920 5040 15972
rect 5356 15920 5408 15972
rect 8208 15920 8260 15972
rect 10876 15963 10928 15972
rect 10876 15929 10885 15963
rect 10885 15929 10919 15963
rect 10919 15929 10928 15963
rect 10876 15920 10928 15929
rect 12992 15988 13044 16040
rect 15200 16056 15252 16108
rect 13820 15988 13872 16040
rect 15108 15988 15160 16040
rect 13912 15920 13964 15972
rect 5264 15852 5316 15904
rect 5632 15895 5684 15904
rect 5632 15861 5641 15895
rect 5641 15861 5675 15895
rect 5675 15861 5684 15895
rect 5632 15852 5684 15861
rect 11060 15852 11112 15904
rect 15660 15920 15712 15972
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 16488 15895 16540 15904
rect 16488 15861 16497 15895
rect 16497 15861 16531 15895
rect 16531 15861 16540 15895
rect 16488 15852 16540 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1676 15648 1728 15700
rect 3056 15691 3108 15700
rect 3056 15657 3065 15691
rect 3065 15657 3099 15691
rect 3099 15657 3108 15691
rect 3056 15648 3108 15657
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 8852 15648 8904 15700
rect 9864 15648 9916 15700
rect 10140 15691 10192 15700
rect 10140 15657 10149 15691
rect 10149 15657 10183 15691
rect 10183 15657 10192 15691
rect 10140 15648 10192 15657
rect 11704 15691 11756 15700
rect 1492 15580 1544 15632
rect 5540 15580 5592 15632
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 11888 15648 11940 15700
rect 12900 15648 12952 15700
rect 14096 15648 14148 15700
rect 14372 15648 14424 15700
rect 15200 15648 15252 15700
rect 16488 15648 16540 15700
rect 1860 15512 1912 15564
rect 3056 15512 3108 15564
rect 3976 15512 4028 15564
rect 4712 15376 4764 15428
rect 6460 15308 6512 15360
rect 9864 15512 9916 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 14464 15580 14516 15632
rect 10692 15512 10744 15564
rect 11796 15512 11848 15564
rect 12072 15512 12124 15564
rect 13636 15512 13688 15564
rect 14096 15512 14148 15564
rect 8208 15419 8260 15428
rect 8208 15385 8217 15419
rect 8217 15385 8251 15419
rect 8251 15385 8260 15419
rect 12256 15444 12308 15496
rect 12992 15444 13044 15496
rect 15752 15487 15804 15496
rect 8208 15376 8260 15385
rect 8300 15308 8352 15360
rect 10140 15308 10192 15360
rect 12072 15308 12124 15360
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 15936 15444 15988 15496
rect 13912 15308 13964 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 572 15036 624 15088
rect 13820 15104 13872 15156
rect 15660 15104 15712 15156
rect 12808 15036 12860 15088
rect 1860 14968 1912 15020
rect 3056 15011 3108 15020
rect 3056 14977 3065 15011
rect 3065 14977 3099 15011
rect 3099 14977 3108 15011
rect 3056 14968 3108 14977
rect 5632 14968 5684 15020
rect 1584 14943 1636 14952
rect 1584 14909 1593 14943
rect 1593 14909 1627 14943
rect 1627 14909 1636 14943
rect 1584 14900 1636 14909
rect 2964 14900 3016 14952
rect 3976 14900 4028 14952
rect 5540 14900 5592 14952
rect 9404 14968 9456 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 12992 14968 13044 15020
rect 13636 15036 13688 15088
rect 14096 14968 14148 15020
rect 14556 14968 14608 15020
rect 15936 14968 15988 15020
rect 8208 14900 8260 14952
rect 8944 14900 8996 14952
rect 11612 14900 11664 14952
rect 15384 14900 15436 14952
rect 5448 14832 5500 14884
rect 5080 14764 5132 14816
rect 10140 14832 10192 14884
rect 12256 14832 12308 14884
rect 12808 14875 12860 14884
rect 12808 14841 12817 14875
rect 12817 14841 12851 14875
rect 12851 14841 12860 14875
rect 12808 14832 12860 14841
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 8300 14764 8352 14816
rect 8668 14764 8720 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 11152 14764 11204 14816
rect 14280 14764 14332 14816
rect 15292 14764 15344 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14560 1728 14612
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 4896 14560 4948 14612
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 1860 14424 1912 14476
rect 3332 14467 3384 14476
rect 3332 14433 3341 14467
rect 3341 14433 3375 14467
rect 3375 14433 3384 14467
rect 3332 14424 3384 14433
rect 1584 14356 1636 14408
rect 5908 14424 5960 14476
rect 8300 14560 8352 14612
rect 9956 14560 10008 14612
rect 11060 14560 11112 14612
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 12624 14560 12676 14612
rect 15568 14560 15620 14612
rect 7656 14492 7708 14544
rect 8484 14492 8536 14544
rect 6920 14424 6972 14476
rect 8668 14424 8720 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 3976 14288 4028 14340
rect 7104 14356 7156 14408
rect 10600 14492 10652 14544
rect 10784 14492 10836 14544
rect 12164 14492 12216 14544
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 12164 14356 12216 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 13084 14356 13136 14408
rect 14556 14356 14608 14408
rect 5080 14288 5132 14340
rect 5632 14220 5684 14272
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 5908 14220 5960 14272
rect 10876 14288 10928 14340
rect 15108 14288 15160 14340
rect 15384 14424 15436 14476
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 18972 14288 19024 14340
rect 10784 14220 10836 14272
rect 11704 14220 11756 14272
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 2780 14016 2832 14025
rect 3332 14016 3384 14068
rect 4712 14016 4764 14068
rect 5632 14016 5684 14068
rect 4252 13948 4304 14000
rect 4620 13948 4672 14000
rect 4896 13948 4948 14000
rect 8484 14016 8536 14068
rect 9956 14016 10008 14068
rect 10968 14016 11020 14068
rect 5908 13880 5960 13932
rect 6460 13880 6512 13932
rect 10140 13948 10192 14000
rect 15200 14016 15252 14068
rect 18604 14016 18656 14068
rect 11612 13948 11664 14000
rect 10876 13923 10928 13932
rect 2044 13812 2096 13864
rect 3240 13812 3292 13864
rect 4804 13812 4856 13864
rect 6828 13812 6880 13864
rect 5724 13787 5776 13796
rect 5724 13753 5733 13787
rect 5733 13753 5767 13787
rect 5767 13753 5776 13787
rect 5724 13744 5776 13753
rect 7104 13812 7156 13864
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 12440 13948 12492 14000
rect 13176 13991 13228 14000
rect 13176 13957 13185 13991
rect 13185 13957 13219 13991
rect 13219 13957 13228 13991
rect 13176 13948 13228 13957
rect 13912 13948 13964 14000
rect 14280 13948 14332 14000
rect 12164 13880 12216 13932
rect 4436 13719 4488 13728
rect 4436 13685 4445 13719
rect 4445 13685 4479 13719
rect 4479 13685 4488 13719
rect 4436 13676 4488 13685
rect 9128 13744 9180 13796
rect 9588 13676 9640 13728
rect 9772 13676 9824 13728
rect 10232 13676 10284 13728
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 15844 13812 15896 13864
rect 13360 13744 13412 13796
rect 10784 13719 10836 13728
rect 10784 13685 10793 13719
rect 10793 13685 10827 13719
rect 10827 13685 10836 13719
rect 10784 13676 10836 13685
rect 11428 13676 11480 13728
rect 11888 13676 11940 13728
rect 12532 13676 12584 13728
rect 14188 13744 14240 13796
rect 15384 13676 15436 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 16396 13676 16448 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 4436 13515 4488 13524
rect 4436 13481 4445 13515
rect 4445 13481 4479 13515
rect 4479 13481 4488 13515
rect 4436 13472 4488 13481
rect 7104 13472 7156 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 9128 13472 9180 13524
rect 11520 13472 11572 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12256 13472 12308 13524
rect 12440 13472 12492 13524
rect 3608 13404 3660 13456
rect 3884 13404 3936 13456
rect 1952 13336 2004 13388
rect 3332 13379 3384 13388
rect 3332 13345 3341 13379
rect 3341 13345 3375 13379
rect 3375 13345 3384 13379
rect 3332 13336 3384 13345
rect 7104 13336 7156 13388
rect 7472 13336 7524 13388
rect 9956 13379 10008 13388
rect 9956 13345 9990 13379
rect 9990 13345 10008 13379
rect 9956 13336 10008 13345
rect 10324 13404 10376 13456
rect 10600 13404 10652 13456
rect 11428 13404 11480 13456
rect 12532 13404 12584 13456
rect 13176 13472 13228 13524
rect 15292 13472 15344 13524
rect 12716 13379 12768 13388
rect 1400 13268 1452 13320
rect 3700 13268 3752 13320
rect 5540 13268 5592 13320
rect 5724 13268 5776 13320
rect 7564 13268 7616 13320
rect 7472 13200 7524 13252
rect 9588 13268 9640 13320
rect 2320 13132 2372 13184
rect 5356 13132 5408 13184
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 14004 13404 14056 13456
rect 14556 13404 14608 13456
rect 15384 13404 15436 13456
rect 14188 13336 14240 13388
rect 11152 13200 11204 13252
rect 11520 13268 11572 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16396 13268 16448 13320
rect 12348 13200 12400 13252
rect 15108 13200 15160 13252
rect 16028 13200 16080 13252
rect 10968 13132 11020 13184
rect 17224 13132 17276 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 5172 12928 5224 12980
rect 6920 12971 6972 12980
rect 6920 12937 6929 12971
rect 6929 12937 6963 12971
rect 6963 12937 6972 12971
rect 6920 12928 6972 12937
rect 1676 12860 1728 12912
rect 2688 12792 2740 12844
rect 4068 12860 4120 12912
rect 10600 12928 10652 12980
rect 11612 12928 11664 12980
rect 11888 12928 11940 12980
rect 12808 12928 12860 12980
rect 14188 12971 14240 12980
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 14556 12928 14608 12980
rect 15752 12928 15804 12980
rect 3700 12792 3752 12844
rect 4160 12792 4212 12844
rect 5448 12792 5500 12844
rect 8208 12860 8260 12912
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 9772 12860 9824 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 4896 12724 4948 12776
rect 5172 12724 5224 12776
rect 5356 12724 5408 12776
rect 9588 12792 9640 12844
rect 7656 12724 7708 12776
rect 10140 12767 10192 12776
rect 10140 12733 10174 12767
rect 10174 12733 10192 12767
rect 10968 12792 11020 12844
rect 11704 12792 11756 12844
rect 12164 12792 12216 12844
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 12256 12767 12308 12776
rect 10140 12724 10192 12733
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 10692 12656 10744 12708
rect 11152 12656 11204 12708
rect 12440 12656 12492 12708
rect 12532 12656 12584 12708
rect 15200 12724 15252 12776
rect 15844 12767 15896 12776
rect 15844 12733 15853 12767
rect 15853 12733 15887 12767
rect 15887 12733 15896 12767
rect 15844 12724 15896 12733
rect 13728 12656 13780 12708
rect 13820 12656 13872 12708
rect 15752 12656 15804 12708
rect 7564 12588 7616 12640
rect 10140 12588 10192 12640
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 11796 12588 11848 12640
rect 12164 12588 12216 12640
rect 14556 12588 14608 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 5540 12384 5592 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 7564 12384 7616 12436
rect 10416 12384 10468 12436
rect 10876 12384 10928 12436
rect 12808 12427 12860 12436
rect 12808 12393 12817 12427
rect 12817 12393 12851 12427
rect 12851 12393 12860 12427
rect 12808 12384 12860 12393
rect 13820 12384 13872 12436
rect 1676 12316 1728 12368
rect 4068 12316 4120 12368
rect 5724 12316 5776 12368
rect 8392 12316 8444 12368
rect 8576 12316 8628 12368
rect 10600 12316 10652 12368
rect 11244 12316 11296 12368
rect 4160 12248 4212 12300
rect 5448 12248 5500 12300
rect 6460 12248 6512 12300
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8300 12248 8352 12300
rect 10416 12248 10468 12300
rect 10784 12248 10836 12300
rect 8024 12180 8076 12189
rect 8484 12180 8536 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 10048 12180 10100 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 12808 12180 12860 12232
rect 13544 12316 13596 12368
rect 14280 12316 14332 12368
rect 15108 12316 15160 12368
rect 17316 12248 17368 12300
rect 12992 12180 13044 12232
rect 11980 12112 12032 12164
rect 13728 12112 13780 12164
rect 2504 12044 2556 12096
rect 2688 12044 2740 12096
rect 3424 12044 3476 12096
rect 5264 12044 5316 12096
rect 11888 12044 11940 12096
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 16856 12044 16908 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 3332 11840 3384 11892
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 4068 11840 4120 11892
rect 6460 11883 6512 11892
rect 6460 11849 6469 11883
rect 6469 11849 6503 11883
rect 6503 11849 6512 11883
rect 6460 11840 6512 11849
rect 8024 11840 8076 11892
rect 8300 11883 8352 11892
rect 8300 11849 8309 11883
rect 8309 11849 8343 11883
rect 8343 11849 8352 11883
rect 8300 11840 8352 11849
rect 9680 11772 9732 11824
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 2872 11636 2924 11688
rect 3976 11679 4028 11688
rect 3976 11645 3985 11679
rect 3985 11645 4019 11679
rect 4019 11645 4028 11679
rect 3976 11636 4028 11645
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 7748 11704 7800 11756
rect 9128 11704 9180 11756
rect 11612 11840 11664 11892
rect 11796 11840 11848 11892
rect 12072 11840 12124 11892
rect 11152 11772 11204 11824
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 12164 11772 12216 11824
rect 13544 11840 13596 11892
rect 13728 11840 13780 11892
rect 1492 11568 1544 11620
rect 3424 11500 3476 11552
rect 3608 11500 3660 11552
rect 4068 11500 4120 11552
rect 4160 11500 4212 11552
rect 7472 11636 7524 11688
rect 5356 11611 5408 11620
rect 5356 11577 5390 11611
rect 5390 11577 5408 11611
rect 5356 11568 5408 11577
rect 10324 11636 10376 11688
rect 12072 11704 12124 11756
rect 11888 11636 11940 11688
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 14556 11840 14608 11892
rect 12440 11704 12492 11713
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7104 11500 7156 11552
rect 7656 11500 7708 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 9220 11500 9272 11552
rect 12532 11568 12584 11620
rect 12808 11568 12860 11620
rect 13544 11568 13596 11620
rect 14372 11568 14424 11620
rect 14648 11568 14700 11620
rect 11060 11500 11112 11552
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 13268 11500 13320 11552
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 15660 11636 15712 11688
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 16856 11568 16908 11620
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 4068 11296 4120 11348
rect 6276 11296 6328 11348
rect 6828 11296 6880 11348
rect 9220 11339 9272 11348
rect 9220 11305 9229 11339
rect 9229 11305 9263 11339
rect 9263 11305 9272 11339
rect 9220 11296 9272 11305
rect 11060 11296 11112 11348
rect 11980 11339 12032 11348
rect 11980 11305 11989 11339
rect 11989 11305 12023 11339
rect 12023 11305 12032 11339
rect 11980 11296 12032 11305
rect 12348 11296 12400 11348
rect 12992 11296 13044 11348
rect 13268 11339 13320 11348
rect 13268 11305 13277 11339
rect 13277 11305 13311 11339
rect 13311 11305 13320 11339
rect 13268 11296 13320 11305
rect 14464 11296 14516 11348
rect 15660 11296 15712 11348
rect 16304 11339 16356 11348
rect 16304 11305 16313 11339
rect 16313 11305 16347 11339
rect 16347 11305 16356 11339
rect 16304 11296 16356 11305
rect 16764 11339 16816 11348
rect 16764 11305 16773 11339
rect 16773 11305 16807 11339
rect 16807 11305 16816 11339
rect 16764 11296 16816 11305
rect 2504 11228 2556 11280
rect 3884 11228 3936 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 1952 11092 2004 11144
rect 4160 11160 4212 11212
rect 6184 11228 6236 11280
rect 8668 11228 8720 11280
rect 10508 11228 10560 11280
rect 12532 11228 12584 11280
rect 13544 11228 13596 11280
rect 4896 11160 4948 11212
rect 5724 11160 5776 11212
rect 10048 11160 10100 11212
rect 12164 11160 12216 11212
rect 13268 11160 13320 11212
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 15476 11228 15528 11280
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 8208 11092 8260 11144
rect 12808 11092 12860 11144
rect 13544 11092 13596 11144
rect 13820 11092 13872 11144
rect 14188 11092 14240 11144
rect 15844 11160 15896 11212
rect 16672 11203 16724 11212
rect 16672 11169 16681 11203
rect 16681 11169 16715 11203
rect 16715 11169 16724 11203
rect 16672 11160 16724 11169
rect 15936 11135 15988 11144
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 3240 10956 3292 11008
rect 4068 10956 4120 11008
rect 6092 10999 6144 11008
rect 6092 10965 6101 10999
rect 6101 10965 6135 10999
rect 6135 10965 6144 10999
rect 6092 10956 6144 10965
rect 9680 11024 9732 11076
rect 10508 11024 10560 11076
rect 11336 11024 11388 11076
rect 12900 11024 12952 11076
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 17408 11024 17460 11076
rect 7472 10956 7524 11008
rect 7748 10956 7800 11008
rect 8576 10956 8628 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 11612 10956 11664 11008
rect 16948 10956 17000 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1676 10752 1728 10804
rect 3516 10752 3568 10804
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 10048 10752 10100 10804
rect 10232 10752 10284 10804
rect 9680 10684 9732 10736
rect 10968 10684 11020 10736
rect 14556 10752 14608 10804
rect 16672 10752 16724 10804
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 4712 10616 4764 10668
rect 4988 10616 5040 10668
rect 5356 10659 5408 10668
rect 5356 10625 5365 10659
rect 5365 10625 5399 10659
rect 5399 10625 5408 10659
rect 5356 10616 5408 10625
rect 9956 10616 10008 10668
rect 11980 10616 12032 10668
rect 12900 10659 12952 10668
rect 3976 10548 4028 10600
rect 6092 10591 6144 10600
rect 6092 10557 6101 10591
rect 6101 10557 6135 10591
rect 6135 10557 6144 10591
rect 6092 10548 6144 10557
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 2872 10480 2924 10532
rect 3700 10480 3752 10532
rect 4988 10480 5040 10532
rect 5448 10480 5500 10532
rect 1584 10412 1636 10464
rect 2136 10412 2188 10464
rect 3332 10412 3384 10464
rect 3792 10412 3844 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5632 10412 5684 10464
rect 6920 10480 6972 10532
rect 6092 10412 6144 10464
rect 6736 10412 6788 10464
rect 8576 10548 8628 10600
rect 10416 10480 10468 10532
rect 12164 10480 12216 10532
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 13544 10616 13596 10668
rect 14188 10616 14240 10668
rect 16120 10684 16172 10736
rect 16856 10684 16908 10736
rect 13912 10548 13964 10600
rect 14556 10480 14608 10532
rect 9956 10412 10008 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 12624 10412 12676 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13544 10412 13596 10464
rect 13728 10412 13780 10464
rect 15292 10616 15344 10668
rect 15936 10616 15988 10668
rect 16672 10616 16724 10668
rect 17316 10616 17368 10668
rect 15108 10412 15160 10464
rect 15384 10412 15436 10464
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 3148 10208 3200 10260
rect 2136 10140 2188 10192
rect 4804 10208 4856 10260
rect 5356 10208 5408 10260
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 6920 10208 6972 10260
rect 8760 10208 8812 10260
rect 12256 10208 12308 10260
rect 12624 10208 12676 10260
rect 4068 10140 4120 10192
rect 13544 10140 13596 10192
rect 3148 10072 3200 10124
rect 5264 10072 5316 10124
rect 5448 10072 5500 10124
rect 9036 10072 9088 10124
rect 10416 10072 10468 10124
rect 10784 10115 10836 10124
rect 10784 10081 10818 10115
rect 10818 10081 10836 10115
rect 10784 10072 10836 10081
rect 11060 10072 11112 10124
rect 12440 10072 12492 10124
rect 13820 10072 13872 10124
rect 14004 10208 14056 10260
rect 15108 10208 15160 10260
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 15384 10072 15436 10124
rect 15936 10140 15988 10192
rect 17040 10072 17092 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 4160 10004 4212 10056
rect 5540 10004 5592 10056
rect 6736 10047 6788 10056
rect 6736 10013 6745 10047
rect 6745 10013 6779 10047
rect 6779 10013 6788 10047
rect 6736 10004 6788 10013
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8208 10004 8260 10056
rect 8576 10004 8628 10056
rect 5632 9936 5684 9988
rect 12348 9936 12400 9988
rect 5356 9868 5408 9920
rect 11612 9868 11664 9920
rect 11980 9868 12032 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 4068 9664 4120 9716
rect 5080 9596 5132 9648
rect 5816 9596 5868 9648
rect 6920 9596 6972 9648
rect 7564 9664 7616 9716
rect 14372 9664 14424 9716
rect 15752 9664 15804 9716
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 6092 9528 6144 9580
rect 7748 9528 7800 9580
rect 10140 9528 10192 9580
rect 1952 9460 2004 9512
rect 3240 9460 3292 9512
rect 4712 9460 4764 9512
rect 4068 9392 4120 9444
rect 6368 9392 6420 9444
rect 7104 9460 7156 9512
rect 7380 9460 7432 9512
rect 8208 9392 8260 9444
rect 8760 9460 8812 9512
rect 9680 9460 9732 9512
rect 9956 9460 10008 9512
rect 12440 9596 12492 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 11060 9528 11112 9580
rect 12072 9528 12124 9580
rect 14556 9571 14608 9580
rect 10508 9460 10560 9512
rect 11612 9460 11664 9512
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 16304 9596 16356 9648
rect 15936 9528 15988 9580
rect 13084 9460 13136 9512
rect 14280 9460 14332 9512
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 5632 9367 5684 9376
rect 5632 9333 5641 9367
rect 5641 9333 5675 9367
rect 5675 9333 5684 9367
rect 5632 9324 5684 9333
rect 5724 9324 5776 9376
rect 6644 9324 6696 9376
rect 8392 9324 8444 9376
rect 10600 9324 10652 9376
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 12348 9392 12400 9444
rect 11980 9324 12032 9376
rect 15016 9392 15068 9444
rect 14188 9324 14240 9376
rect 15200 9324 15252 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9120 2280 9172
rect 4988 9120 5040 9172
rect 5356 9120 5408 9172
rect 2136 9052 2188 9104
rect 3424 9052 3476 9104
rect 3792 9052 3844 9104
rect 1952 8984 2004 9036
rect 3976 8984 4028 9036
rect 6644 9052 6696 9104
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5908 8984 5960 9036
rect 6092 9027 6144 9036
rect 6092 8993 6126 9027
rect 6126 8993 6144 9027
rect 6092 8984 6144 8993
rect 7380 9120 7432 9172
rect 7748 9095 7800 9104
rect 7748 9061 7782 9095
rect 7782 9061 7800 9095
rect 7748 9052 7800 9061
rect 8208 9120 8260 9172
rect 10876 9120 10928 9172
rect 12808 9120 12860 9172
rect 14372 9120 14424 9172
rect 9956 8984 10008 9036
rect 16212 9052 16264 9104
rect 6828 8916 6880 8968
rect 8668 8916 8720 8968
rect 3884 8848 3936 8900
rect 3332 8780 3384 8832
rect 5816 8848 5868 8900
rect 10324 8848 10376 8900
rect 11980 8984 12032 9036
rect 12532 8984 12584 9036
rect 11060 8916 11112 8968
rect 12348 8916 12400 8968
rect 12716 8916 12768 8968
rect 14096 8984 14148 9036
rect 14372 9027 14424 9036
rect 14372 8993 14381 9027
rect 14381 8993 14415 9027
rect 14415 8993 14424 9027
rect 14372 8984 14424 8993
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 13544 8916 13596 8968
rect 14188 8848 14240 8900
rect 9404 8780 9456 8832
rect 15752 8780 15804 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 5724 8576 5776 8628
rect 5908 8576 5960 8628
rect 6460 8576 6512 8628
rect 7104 8576 7156 8628
rect 7196 8576 7248 8628
rect 1860 8440 1912 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 3700 8440 3752 8492
rect 4068 8440 4120 8492
rect 5264 8508 5316 8560
rect 5816 8508 5868 8560
rect 4712 8440 4764 8492
rect 5540 8440 5592 8492
rect 5632 8372 5684 8424
rect 7380 8440 7432 8492
rect 15016 8576 15068 8628
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 10324 8508 10376 8560
rect 14280 8508 14332 8560
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 8760 8372 8812 8424
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 11152 8440 11204 8492
rect 10140 8372 10192 8424
rect 13636 8440 13688 8492
rect 12256 8372 12308 8424
rect 13544 8372 13596 8424
rect 15384 8372 15436 8424
rect 4068 8304 4120 8356
rect 6736 8304 6788 8356
rect 4804 8236 4856 8288
rect 5356 8236 5408 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6000 8236 6052 8288
rect 6644 8236 6696 8288
rect 6828 8236 6880 8288
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 11152 8304 11204 8356
rect 11612 8304 11664 8356
rect 12532 8304 12584 8356
rect 8760 8236 8812 8245
rect 10968 8236 11020 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 14372 8304 14424 8356
rect 14556 8347 14608 8356
rect 14556 8313 14590 8347
rect 14590 8313 14608 8347
rect 14556 8304 14608 8313
rect 17224 8304 17276 8356
rect 15568 8236 15620 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3884 8032 3936 8084
rect 5448 8032 5500 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7472 8032 7524 8084
rect 8944 8032 8996 8084
rect 11336 8032 11388 8084
rect 14372 8032 14424 8084
rect 15016 8032 15068 8084
rect 15752 8075 15804 8084
rect 15752 8041 15761 8075
rect 15761 8041 15795 8075
rect 15795 8041 15804 8075
rect 15752 8032 15804 8041
rect 2044 7964 2096 8016
rect 2228 7964 2280 8016
rect 4068 7964 4120 8016
rect 1492 7939 1544 7948
rect 1492 7905 1501 7939
rect 1501 7905 1535 7939
rect 1535 7905 1544 7939
rect 1492 7896 1544 7905
rect 5540 7896 5592 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 8208 7871 8260 7880
rect 2872 7692 2924 7744
rect 5356 7692 5408 7744
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8944 7760 8996 7812
rect 7656 7692 7708 7744
rect 9128 7828 9180 7880
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 9680 7760 9732 7812
rect 9772 7692 9824 7744
rect 10416 7692 10468 7744
rect 12624 7964 12676 8016
rect 11704 7896 11756 7948
rect 13636 7896 13688 7948
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 14556 7828 14608 7880
rect 13544 7692 13596 7744
rect 15660 7692 15712 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2872 7352 2924 7404
rect 4252 7488 4304 7540
rect 5908 7488 5960 7540
rect 6184 7488 6236 7540
rect 8760 7488 8812 7540
rect 11060 7488 11112 7540
rect 8484 7420 8536 7472
rect 10140 7420 10192 7472
rect 13820 7420 13872 7472
rect 14832 7420 14884 7472
rect 4620 7352 4672 7404
rect 4804 7352 4856 7404
rect 3332 7284 3384 7336
rect 5264 7352 5316 7404
rect 6736 7284 6788 7336
rect 8852 7284 8904 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9680 7352 9732 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 13636 7352 13688 7404
rect 3608 7216 3660 7268
rect 3792 7259 3844 7268
rect 3792 7225 3801 7259
rect 3801 7225 3835 7259
rect 3835 7225 3844 7259
rect 3792 7216 3844 7225
rect 6460 7216 6512 7268
rect 7104 7259 7156 7268
rect 7104 7225 7138 7259
rect 7138 7225 7156 7259
rect 7104 7216 7156 7225
rect 7288 7216 7340 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 3056 7148 3108 7200
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 6276 7148 6328 7200
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 10968 7327 11020 7336
rect 10968 7293 11002 7327
rect 11002 7293 11020 7327
rect 10968 7284 11020 7293
rect 12624 7284 12676 7336
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 15384 7284 15436 7336
rect 15568 7284 15620 7336
rect 11152 7216 11204 7268
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 13544 7148 13596 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 16672 7216 16724 7268
rect 17684 7216 17736 7268
rect 17040 7148 17092 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 5540 6987 5592 6996
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 10048 6944 10100 6996
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 14464 6944 14516 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 2228 6876 2280 6928
rect 2872 6808 2924 6860
rect 4712 6876 4764 6928
rect 6736 6876 6788 6928
rect 4252 6808 4304 6860
rect 5264 6808 5316 6860
rect 6184 6808 6236 6860
rect 9128 6876 9180 6928
rect 1860 6740 1912 6792
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 8208 6808 8260 6860
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 12072 6876 12124 6928
rect 12532 6876 12584 6928
rect 8944 6808 8996 6817
rect 10784 6808 10836 6860
rect 3240 6672 3292 6724
rect 1952 6604 2004 6656
rect 5632 6604 5684 6656
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 7196 6604 7248 6656
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 9128 6672 9180 6724
rect 9312 6672 9364 6724
rect 11152 6672 11204 6724
rect 12440 6740 12492 6792
rect 10968 6604 11020 6656
rect 12164 6604 12216 6656
rect 13360 6604 13412 6656
rect 15568 6808 15620 6860
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14648 6740 14700 6792
rect 17040 6808 17092 6860
rect 19156 6851 19208 6860
rect 19156 6817 19190 6851
rect 19190 6817 19208 6851
rect 19156 6808 19208 6817
rect 18880 6783 18932 6792
rect 13912 6672 13964 6724
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 14096 6604 14148 6656
rect 14464 6604 14516 6656
rect 15200 6604 15252 6656
rect 15660 6604 15712 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 1492 6400 1544 6452
rect 1768 6400 1820 6452
rect 3884 6443 3936 6452
rect 3884 6409 3893 6443
rect 3893 6409 3927 6443
rect 3927 6409 3936 6443
rect 3884 6400 3936 6409
rect 5816 6400 5868 6452
rect 11152 6400 11204 6452
rect 15752 6400 15804 6452
rect 6828 6332 6880 6384
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2872 6264 2924 6316
rect 4620 6264 4672 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 8208 6264 8260 6316
rect 8852 6264 8904 6316
rect 1400 6196 1452 6248
rect 3056 6196 3108 6248
rect 5632 6196 5684 6248
rect 7472 6196 7524 6248
rect 7564 6196 7616 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10784 6332 10836 6384
rect 12348 6332 12400 6384
rect 10968 6264 11020 6316
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 6000 6128 6052 6180
rect 11060 6196 11112 6248
rect 10968 6128 11020 6180
rect 11980 6264 12032 6316
rect 11704 6196 11756 6248
rect 20260 6332 20312 6384
rect 13728 6264 13780 6316
rect 14464 6264 14516 6316
rect 15108 6264 15160 6316
rect 15292 6264 15344 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 17132 6307 17184 6316
rect 17132 6273 17141 6307
rect 17141 6273 17175 6307
rect 17175 6273 17184 6307
rect 17132 6264 17184 6273
rect 13360 6196 13412 6248
rect 3516 6060 3568 6112
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 4988 6060 5040 6112
rect 6920 6060 6972 6112
rect 7656 6060 7708 6112
rect 8300 6060 8352 6112
rect 9588 6060 9640 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 10600 6060 10652 6112
rect 11152 6060 11204 6112
rect 19800 6128 19852 6180
rect 11612 6060 11664 6112
rect 14280 6060 14332 6112
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15200 6060 15252 6069
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16764 6060 16816 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 2044 5856 2096 5908
rect 3792 5856 3844 5908
rect 4712 5856 4764 5908
rect 5356 5856 5408 5908
rect 6276 5856 6328 5908
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7472 5856 7524 5908
rect 1952 5788 2004 5840
rect 6184 5788 6236 5840
rect 5264 5720 5316 5772
rect 6736 5720 6788 5772
rect 8116 5788 8168 5840
rect 10048 5788 10100 5840
rect 10968 5856 11020 5908
rect 12440 5856 12492 5908
rect 11888 5788 11940 5840
rect 14004 5856 14056 5908
rect 15568 5856 15620 5908
rect 15936 5788 15988 5840
rect 9772 5720 9824 5772
rect 10324 5720 10376 5772
rect 11704 5763 11756 5772
rect 11704 5729 11713 5763
rect 11713 5729 11747 5763
rect 11747 5729 11756 5763
rect 11704 5720 11756 5729
rect 15108 5720 15160 5772
rect 17040 5720 17092 5772
rect 17132 5720 17184 5772
rect 17868 5720 17920 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 5080 5652 5132 5704
rect 5632 5652 5684 5704
rect 6368 5652 6420 5704
rect 7196 5695 7248 5704
rect 4344 5584 4396 5636
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 8208 5695 8260 5704
rect 6644 5516 6696 5568
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 8300 5584 8352 5636
rect 7012 5516 7064 5568
rect 8668 5516 8720 5568
rect 9128 5652 9180 5704
rect 11060 5652 11112 5704
rect 12164 5652 12216 5704
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 15384 5652 15436 5704
rect 10784 5516 10836 5568
rect 11152 5516 11204 5568
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 15108 5516 15160 5568
rect 15844 5516 15896 5568
rect 15936 5516 15988 5568
rect 18880 5695 18932 5704
rect 17132 5516 17184 5568
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 17868 5516 17920 5568
rect 17960 5516 18012 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 4804 5244 4856 5296
rect 1952 5176 2004 5228
rect 4160 5176 4212 5228
rect 4712 5176 4764 5228
rect 1400 5108 1452 5160
rect 2228 5108 2280 5160
rect 3332 5108 3384 5160
rect 3884 5108 3936 5160
rect 10140 5312 10192 5364
rect 10048 5244 10100 5296
rect 10692 5244 10744 5296
rect 10784 5244 10836 5296
rect 11704 5244 11756 5296
rect 14004 5244 14056 5296
rect 5724 5108 5776 5160
rect 10508 5176 10560 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 10600 5108 10652 5160
rect 11152 5108 11204 5160
rect 12072 5176 12124 5228
rect 12348 5176 12400 5228
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 12164 5108 12216 5160
rect 12808 5108 12860 5160
rect 13544 5108 13596 5160
rect 15384 5108 15436 5160
rect 15936 5108 15988 5160
rect 17224 5108 17276 5160
rect 17868 5108 17920 5160
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 6920 5040 6972 5092
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 4068 4972 4120 5024
rect 5080 4972 5132 5024
rect 6368 4972 6420 5024
rect 6828 4972 6880 5024
rect 7380 4972 7432 5024
rect 8668 5040 8720 5092
rect 10508 5040 10560 5092
rect 12900 5083 12952 5092
rect 12900 5049 12909 5083
rect 12909 5049 12943 5083
rect 12943 5049 12952 5083
rect 12900 5040 12952 5049
rect 13820 5040 13872 5092
rect 15016 5040 15068 5092
rect 16948 5040 17000 5092
rect 9680 4972 9732 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 13728 4972 13780 5024
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 16856 4972 16908 5024
rect 20628 4972 20680 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 6644 4768 6696 4820
rect 9956 4768 10008 4820
rect 11060 4768 11112 4820
rect 11704 4768 11756 4820
rect 12440 4768 12492 4820
rect 2044 4700 2096 4752
rect 3792 4700 3844 4752
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 5632 4632 5684 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 7380 4700 7432 4752
rect 9404 4700 9456 4752
rect 12716 4700 12768 4752
rect 13268 4700 13320 4752
rect 14188 4700 14240 4752
rect 15200 4768 15252 4820
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16396 4768 16448 4820
rect 8760 4675 8812 4684
rect 8760 4641 8769 4675
rect 8769 4641 8803 4675
rect 8803 4641 8812 4675
rect 8760 4632 8812 4641
rect 9220 4632 9272 4684
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 6828 4607 6880 4616
rect 204 4428 256 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 8852 4607 8904 4616
rect 5356 4496 5408 4548
rect 8852 4573 8861 4607
rect 8861 4573 8895 4607
rect 8895 4573 8904 4607
rect 8852 4564 8904 4573
rect 9588 4564 9640 4616
rect 10048 4632 10100 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 11612 4632 11664 4684
rect 12072 4632 12124 4684
rect 12256 4675 12308 4684
rect 12256 4641 12265 4675
rect 12265 4641 12299 4675
rect 12299 4641 12308 4675
rect 12256 4632 12308 4641
rect 16764 4632 16816 4684
rect 11060 4564 11112 4616
rect 12348 4607 12400 4616
rect 10968 4496 11020 4548
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 17132 4564 17184 4616
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 6276 4428 6328 4480
rect 7196 4428 7248 4480
rect 9772 4471 9824 4480
rect 9772 4437 9781 4471
rect 9781 4437 9815 4471
rect 9815 4437 9824 4471
rect 9772 4428 9824 4437
rect 11796 4428 11848 4480
rect 12624 4428 12676 4480
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 16672 4428 16724 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2228 4224 2280 4276
rect 1952 4088 2004 4140
rect 2320 4156 2372 4208
rect 2688 4156 2740 4208
rect 3240 4156 3292 4208
rect 1768 4020 1820 4072
rect 2964 4020 3016 4072
rect 4436 4088 4488 4140
rect 6920 4156 6972 4208
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5632 4088 5684 4140
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 8760 4224 8812 4276
rect 7840 4156 7892 4208
rect 12072 4224 12124 4276
rect 14924 4224 14976 4276
rect 9588 4156 9640 4208
rect 8944 4088 8996 4140
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9772 4088 9824 4140
rect 11152 4156 11204 4208
rect 10968 4088 11020 4140
rect 11244 4131 11296 4140
rect 11244 4097 11253 4131
rect 11253 4097 11287 4131
rect 11287 4097 11296 4131
rect 11244 4088 11296 4097
rect 11704 4088 11756 4140
rect 12256 4088 12308 4140
rect 13728 4156 13780 4208
rect 4896 4020 4948 4072
rect 6276 4020 6328 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 9680 4020 9732 4072
rect 2780 3884 2832 3936
rect 3148 3884 3200 3936
rect 9404 3952 9456 4004
rect 3792 3884 3844 3936
rect 4528 3884 4580 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 9312 3884 9364 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10048 3884 10100 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 10784 3884 10836 3936
rect 14556 4088 14608 4140
rect 15108 4088 15160 4140
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 15844 4156 15896 4208
rect 18512 4020 18564 4072
rect 13360 3952 13412 4004
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12992 3884 13044 3936
rect 14096 3884 14148 3936
rect 16672 3995 16724 4004
rect 16672 3961 16681 3995
rect 16681 3961 16715 3995
rect 16715 3961 16724 3995
rect 16672 3952 16724 3961
rect 14556 3884 14608 3936
rect 15200 3884 15252 3936
rect 15292 3884 15344 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 18788 3884 18840 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3332 3680 3384 3732
rect 3424 3680 3476 3732
rect 4436 3680 4488 3732
rect 5080 3680 5132 3732
rect 7564 3680 7616 3732
rect 8852 3680 8904 3732
rect 9496 3680 9548 3732
rect 9772 3680 9824 3732
rect 9864 3680 9916 3732
rect 10232 3680 10284 3732
rect 10600 3680 10652 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 15200 3680 15252 3732
rect 1400 3544 1452 3596
rect 1952 3587 2004 3596
rect 1952 3553 1986 3587
rect 1986 3553 2004 3587
rect 1952 3544 2004 3553
rect 6736 3612 6788 3664
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 6000 3587 6052 3596
rect 6000 3553 6034 3587
rect 6034 3553 6052 3587
rect 6000 3544 6052 3553
rect 6828 3544 6880 3596
rect 9680 3612 9732 3664
rect 11244 3655 11296 3664
rect 2964 3476 3016 3528
rect 3700 3476 3752 3528
rect 5264 3476 5316 3528
rect 5632 3476 5684 3528
rect 6920 3476 6972 3528
rect 7748 3476 7800 3528
rect 9128 3544 9180 3596
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 11244 3621 11278 3655
rect 11278 3621 11296 3655
rect 11244 3612 11296 3621
rect 9220 3519 9272 3528
rect 8760 3408 8812 3460
rect 8944 3408 8996 3460
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 10048 3476 10100 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 9588 3408 9640 3460
rect 12072 3476 12124 3528
rect 14556 3612 14608 3664
rect 22468 3680 22520 3732
rect 15476 3612 15528 3664
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 15108 3544 15160 3596
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 12808 3408 12860 3460
rect 15292 3476 15344 3528
rect 16764 3544 16816 3596
rect 16948 3544 17000 3596
rect 14464 3408 14516 3460
rect 20260 3476 20312 3528
rect 21548 3408 21600 3460
rect 7380 3340 7432 3392
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 11888 3340 11940 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 12900 3340 12952 3392
rect 15936 3340 15988 3392
rect 16488 3383 16540 3392
rect 16488 3349 16497 3383
rect 16497 3349 16531 3383
rect 16531 3349 16540 3383
rect 16488 3340 16540 3349
rect 22008 3340 22060 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 1952 3136 2004 3188
rect 6000 3136 6052 3188
rect 6644 3136 6696 3188
rect 8576 3136 8628 3188
rect 8668 3136 8720 3188
rect 5540 3068 5592 3120
rect 2320 2907 2372 2916
rect 2320 2873 2354 2907
rect 2354 2873 2372 2907
rect 2320 2864 2372 2873
rect 4068 3000 4120 3052
rect 5724 3000 5776 3052
rect 5356 2932 5408 2984
rect 7380 2975 7432 2984
rect 7380 2941 7414 2975
rect 7414 2941 7432 2975
rect 8760 3068 8812 3120
rect 10232 3136 10284 3188
rect 8208 3000 8260 3052
rect 11060 3136 11112 3188
rect 12072 3136 12124 3188
rect 19432 3136 19484 3188
rect 7380 2932 7432 2941
rect 1584 2796 1636 2848
rect 3516 2796 3568 2848
rect 5264 2864 5316 2916
rect 8116 2864 8168 2916
rect 8668 2932 8720 2984
rect 9128 2932 9180 2984
rect 11060 3000 11112 3052
rect 12532 3068 12584 3120
rect 15568 3068 15620 3120
rect 12808 2975 12860 2984
rect 12808 2941 12842 2975
rect 12842 2941 12860 2975
rect 8300 2796 8352 2848
rect 9588 2864 9640 2916
rect 11152 2864 11204 2916
rect 11980 2864 12032 2916
rect 12808 2932 12860 2941
rect 13544 2932 13596 2984
rect 15660 2932 15712 2984
rect 15936 2932 15988 2984
rect 14464 2907 14516 2916
rect 8760 2796 8812 2848
rect 9220 2796 9272 2848
rect 11060 2796 11112 2848
rect 11336 2839 11388 2848
rect 11336 2805 11345 2839
rect 11345 2805 11379 2839
rect 11379 2805 11388 2839
rect 11336 2796 11388 2805
rect 12440 2796 12492 2848
rect 14464 2873 14498 2907
rect 14498 2873 14516 2907
rect 14464 2864 14516 2873
rect 15016 2864 15068 2916
rect 15108 2796 15160 2848
rect 17316 2932 17368 2984
rect 16672 2796 16724 2848
rect 16948 2796 17000 2848
rect 18512 2796 18564 2848
rect 19708 2796 19760 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2136 2592 2188 2644
rect 3148 2524 3200 2576
rect 3976 2592 4028 2644
rect 4712 2592 4764 2644
rect 7564 2592 7616 2644
rect 3516 2524 3568 2576
rect 7196 2524 7248 2576
rect 8208 2592 8260 2644
rect 9956 2592 10008 2644
rect 10140 2592 10192 2644
rect 11704 2592 11756 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 14556 2592 14608 2644
rect 16672 2592 16724 2644
rect 2688 2456 2740 2508
rect 5264 2456 5316 2508
rect 5908 2388 5960 2440
rect 2780 2320 2832 2372
rect 8668 2456 8720 2508
rect 9680 2524 9732 2576
rect 10784 2567 10836 2576
rect 10784 2533 10793 2567
rect 10793 2533 10827 2567
rect 10827 2533 10836 2567
rect 10784 2524 10836 2533
rect 11888 2456 11940 2508
rect 8300 2388 8352 2440
rect 9220 2388 9272 2440
rect 11060 2388 11112 2440
rect 11152 2388 11204 2440
rect 13452 2524 13504 2576
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13360 2499 13412 2508
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 16304 2524 16356 2576
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 17684 2499 17736 2508
rect 17684 2465 17693 2499
rect 17693 2465 17727 2499
rect 17727 2465 17736 2499
rect 17684 2456 17736 2465
rect 17960 2456 18012 2508
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 20260 2499 20312 2508
rect 20260 2465 20269 2499
rect 20269 2465 20303 2499
rect 20303 2465 20312 2499
rect 20260 2456 20312 2465
rect 13084 2320 13136 2372
rect 13820 2320 13872 2372
rect 16028 2320 16080 2372
rect 11888 2252 11940 2304
rect 13176 2252 13228 2304
rect 13636 2252 13688 2304
rect 17408 2252 17460 2304
rect 17960 2252 18012 2304
rect 19248 2252 19300 2304
rect 20168 2252 20220 2304
rect 21088 2252 21140 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 664 2048 716 2100
rect 6920 2048 6972 2100
rect 2044 1980 2096 2032
rect 3700 1980 3752 2032
rect 2504 1912 2556 1964
rect 8944 1912 8996 1964
rect 1124 1844 1176 1896
rect 6736 1844 6788 1896
<< metal2 >>
rect 202 22000 258 22800
rect 570 22000 626 22800
rect 1030 22000 1086 22800
rect 1490 22000 1546 22800
rect 1950 22000 2006 22800
rect 2410 22000 2466 22800
rect 2870 22000 2926 22800
rect 3330 22000 3386 22800
rect 3514 22128 3570 22137
rect 3514 22063 3570 22072
rect 216 17105 244 22000
rect 202 17096 258 17105
rect 202 17031 258 17040
rect 584 15094 612 22000
rect 1044 17610 1072 22000
rect 1504 18426 1532 22000
rect 1964 19938 1992 22000
rect 1964 19910 2176 19938
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 19281 1992 19654
rect 2056 19310 2084 19790
rect 2044 19304 2096 19310
rect 1950 19272 2006 19281
rect 2044 19246 2096 19252
rect 1950 19207 2006 19216
rect 1950 18864 2006 18873
rect 1950 18799 1952 18808
rect 2004 18799 2006 18808
rect 1952 18770 2004 18776
rect 2148 18737 2176 19910
rect 1674 18728 1730 18737
rect 1674 18663 1676 18672
rect 1728 18663 1730 18672
rect 2134 18728 2190 18737
rect 2134 18663 2190 18672
rect 1676 18634 1728 18640
rect 1492 18420 1544 18426
rect 1492 18362 1544 18368
rect 1490 18320 1546 18329
rect 1490 18255 1546 18264
rect 1032 17604 1084 17610
rect 1032 17546 1084 17552
rect 1504 16794 1532 18255
rect 1952 18216 2004 18222
rect 2424 18193 2452 22000
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2792 20058 2820 20159
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2700 19378 2728 19858
rect 2884 19446 2912 22000
rect 3054 21176 3110 21185
rect 3054 21111 3110 21120
rect 3068 20058 3096 21111
rect 3344 20754 3372 22000
rect 3252 20726 3372 20754
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 1952 18158 2004 18164
rect 2410 18184 2466 18193
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1688 17785 1716 17818
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1582 17368 1638 17377
rect 1582 17303 1638 17312
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 1596 16250 1624 17303
rect 1780 16726 1808 17682
rect 1872 17338 1900 17682
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1964 17134 1992 18158
rect 2410 18119 2466 18128
rect 2516 17785 2544 18362
rect 2792 17814 2820 18770
rect 2884 17882 2912 19110
rect 3160 18902 3188 19246
rect 3148 18896 3200 18902
rect 3148 18838 3200 18844
rect 3252 18630 3280 20726
rect 3330 20632 3386 20641
rect 3330 20567 3386 20576
rect 3344 19514 3372 20567
rect 3422 19680 3478 19689
rect 3422 19615 3478 19624
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 2976 17882 3004 18566
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3068 17814 3096 18022
rect 2780 17808 2832 17814
rect 2502 17776 2558 17785
rect 2780 17750 2832 17756
rect 3056 17808 3108 17814
rect 3056 17750 3108 17756
rect 2502 17711 2558 17720
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2516 16794 2544 17138
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 1674 16416 1730 16425
rect 1674 16351 1730 16360
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1504 15638 1532 15982
rect 1688 15706 1716 16351
rect 2148 16114 2176 16526
rect 2884 16522 2912 17070
rect 2976 16794 3004 17070
rect 3054 16824 3110 16833
rect 2964 16788 3016 16794
rect 3054 16759 3110 16768
rect 2964 16730 3016 16736
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2792 16046 2820 16390
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 1766 15872 1822 15881
rect 1766 15807 1822 15816
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1492 15632 1544 15638
rect 1492 15574 1544 15580
rect 1674 15464 1730 15473
rect 1674 15399 1730 15408
rect 572 15088 624 15094
rect 572 15030 624 15036
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1596 14414 1624 14894
rect 1688 14618 1716 15399
rect 1780 15162 1808 15807
rect 3068 15706 3096 16759
rect 3160 16114 3188 17682
rect 3252 17678 3280 18022
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3252 17066 3280 17614
rect 3436 17490 3464 19615
rect 3528 18034 3556 22063
rect 3790 22000 3846 22800
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 3606 21584 3662 21593
rect 3606 21519 3662 21528
rect 3620 20058 3648 21519
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3804 19360 3832 22000
rect 4080 21842 4108 22471
rect 4250 22000 4306 22800
rect 4710 22000 4766 22800
rect 5170 22000 5226 22800
rect 5630 22000 5686 22800
rect 6090 22000 6146 22800
rect 6550 22000 6606 22800
rect 7010 22000 7066 22800
rect 7470 22000 7526 22800
rect 7930 22000 7986 22800
rect 8390 22000 8446 22800
rect 8850 22000 8906 22800
rect 9310 22000 9366 22800
rect 9770 22000 9826 22800
rect 10230 22000 10286 22800
rect 10690 22000 10746 22800
rect 11150 22000 11206 22800
rect 11610 22000 11666 22800
rect 11978 22000 12034 22800
rect 12438 22000 12494 22800
rect 12898 22000 12954 22800
rect 13358 22000 13414 22800
rect 13818 22000 13874 22800
rect 14278 22000 14334 22800
rect 14738 22000 14794 22800
rect 15198 22000 15254 22800
rect 15658 22000 15714 22800
rect 16118 22000 16174 22800
rect 16578 22000 16634 22800
rect 17038 22000 17094 22800
rect 17498 22000 17554 22800
rect 17958 22000 18014 22800
rect 18418 22000 18474 22800
rect 18878 22000 18934 22800
rect 19338 22000 19394 22800
rect 19798 22000 19854 22800
rect 20258 22000 20314 22800
rect 20718 22000 20774 22800
rect 21178 22000 21234 22800
rect 21638 22000 21694 22800
rect 22098 22000 22154 22800
rect 22558 22000 22614 22800
rect 4264 21962 4292 22000
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4080 21814 4292 21842
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3804 19332 4016 19360
rect 3792 19236 3844 19242
rect 3792 19178 3844 19184
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3712 18426 3740 18702
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3804 18154 3832 19178
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3528 18006 3648 18034
rect 3620 17610 3648 18006
rect 3790 17640 3846 17649
rect 3608 17604 3660 17610
rect 3790 17575 3846 17584
rect 3608 17546 3660 17552
rect 3436 17462 3556 17490
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3252 15994 3280 16662
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 16114 3372 16594
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3436 16250 3464 16526
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3160 15966 3280 15994
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1872 15026 1900 15506
rect 3068 15026 3096 15506
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2976 14618 3004 14894
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2778 14512 2834 14521
rect 1860 14476 1912 14482
rect 2778 14447 2834 14456
rect 1860 14418 1912 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1582 13560 1638 13569
rect 1582 13495 1638 13504
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12782 1440 13262
rect 1596 12986 1624 13495
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1688 12374 1716 12854
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1492 11620 1544 11626
rect 1492 11562 1544 11568
rect 1504 11218 1532 11562
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1688 10810 1716 11630
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1872 8498 1900 14418
rect 2792 14074 2820 14447
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2778 13968 2834 13977
rect 2778 13903 2834 13912
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 12986 1992 13330
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1964 9518 1992 11086
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1964 9042 1992 9454
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1964 8378 1992 8978
rect 1872 8350 1992 8378
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6254 1440 7142
rect 1504 6458 1532 7890
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 6458 1808 7142
rect 1872 6798 1900 8350
rect 2056 8022 2084 13806
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12782 2360 13126
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2700 12102 2728 12786
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2516 11286 2544 12038
rect 2792 11354 2820 13903
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2504 11280 2556 11286
rect 2884 11234 2912 11630
rect 2504 11222 2556 11228
rect 2792 11206 2912 11234
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10198 2176 10406
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9110 2176 9998
rect 2240 9178 2268 10610
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2240 8022 2268 9114
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5166 1440 5646
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 204 4480 256 4486
rect 204 4422 256 4428
rect 216 800 244 4422
rect 1412 3602 1440 5102
rect 1872 4690 1900 6734
rect 1964 6662 1992 7346
rect 2240 6934 2268 7822
rect 2792 7206 2820 11206
rect 2872 10532 2924 10538
rect 2872 10474 2924 10480
rect 2884 8634 2912 10474
rect 3160 10266 3188 15966
rect 3238 14920 3294 14929
rect 3238 14855 3294 14864
rect 3252 13870 3280 14855
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 14074 3372 14418
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3344 11898 3372 13330
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3436 11558 3464 12038
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10674 3280 10950
rect 3436 10690 3464 11494
rect 3528 10810 3556 17462
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 3620 11898 3648 13398
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3712 12850 3740 13262
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3240 10668 3292 10674
rect 3436 10662 3556 10690
rect 3240 10610 3292 10616
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7410 2912 7686
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2228 6928 2280 6934
rect 2228 6870 2280 6876
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 5846 1992 6598
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5914 2084 6258
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1964 4146 1992 5170
rect 2056 4758 2084 5850
rect 2240 5166 2268 6870
rect 2792 6202 2820 7142
rect 2884 6866 2912 7346
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6322 2912 6802
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2792 6174 2912 6202
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 664 2100 716 2106
rect 664 2042 716 2048
rect 676 800 704 2042
rect 1124 1896 1176 1902
rect 1124 1838 1176 1844
rect 1136 800 1164 1838
rect 1596 800 1624 2790
rect 1780 2553 1808 4014
rect 1964 3602 1992 4082
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3194 1992 3538
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2148 2650 2176 4966
rect 2240 4282 2268 4966
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 2332 2922 2360 4150
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 1766 2544 1822 2553
rect 2700 2514 2728 4150
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 1766 2479 1822 2488
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2792 2378 2820 3878
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2884 2145 2912 6174
rect 2976 4078 3004 10202
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6254 3096 7142
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3160 3942 3188 10066
rect 3252 10062 3280 10610
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9518 3280 9998
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3344 8922 3372 10406
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9110 3464 9318
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3252 8894 3372 8922
rect 3252 7426 3280 8894
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8498 3372 8774
rect 3436 8498 3464 9046
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3252 7398 3464 7426
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3252 6361 3280 6666
rect 3238 6352 3294 6361
rect 3238 6287 3294 6296
rect 3344 5166 3372 7278
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4214 3280 4422
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3148 3936 3200 3942
rect 3200 3896 3280 3924
rect 3148 3878 3200 3884
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 3146 3496 3202 3505
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 2056 800 2084 1974
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 2516 800 2544 1906
rect 2976 800 3004 3470
rect 3146 3431 3202 3440
rect 3160 2582 3188 3431
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3252 1601 3280 3896
rect 3344 3738 3372 5102
rect 3436 3913 3464 7398
rect 3528 6118 3556 10662
rect 3620 7274 3648 11494
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3712 9586 3740 10474
rect 3804 10470 3832 17575
rect 3896 17542 3924 18770
rect 3988 18034 4016 19332
rect 4080 19310 4108 19790
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3988 18006 4108 18034
rect 4080 17762 4108 18006
rect 4172 17882 4200 19110
rect 4264 18698 4292 21814
rect 4632 19972 4660 21898
rect 4724 20074 4752 22000
rect 4724 20046 5120 20074
rect 4988 19984 5040 19990
rect 4632 19944 4752 19972
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4356 18612 4384 18702
rect 4325 18584 4384 18612
rect 4325 18578 4353 18584
rect 4264 18550 4353 18578
rect 4264 18222 4292 18550
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4724 18222 4752 19944
rect 4988 19926 5040 19932
rect 5000 19310 5028 19926
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4816 18766 4844 19246
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4080 17734 4200 17762
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3896 16726 3924 17478
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3988 16522 4016 17138
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3988 15570 4016 16458
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3988 14958 4016 15506
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3988 14346 4016 14894
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3896 12617 3924 13398
rect 3988 12764 4016 14282
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4080 12918 4108 12951
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4172 12850 4200 17734
rect 4264 17202 4292 18158
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16726 4292 16934
rect 4724 16794 4752 17002
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4264 16114 4292 16662
rect 4724 16658 4752 16730
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4724 14074 4752 15370
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 4620 14000 4672 14006
rect 4672 13948 4752 13954
rect 4620 13942 4752 13948
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3988 12736 4108 12764
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3974 12472 4030 12481
rect 3974 12407 4030 12416
rect 3988 11694 4016 12407
rect 4080 12374 4108 12736
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4066 12064 4122 12073
rect 4066 11999 4122 12008
rect 4080 11898 4108 11999
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11762 4200 12242
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3976 11688 4028 11694
rect 3882 11656 3938 11665
rect 3976 11630 4028 11636
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3882 11591 3938 11600
rect 3896 11286 3924 11591
rect 4080 11558 4108 11630
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 4080 11121 4108 11290
rect 4172 11218 4200 11494
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10713 4108 10950
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3988 9602 4016 10542
rect 4068 10192 4120 10198
rect 4066 10160 4068 10169
rect 4120 10160 4122 10169
rect 4066 10095 4122 10104
rect 4172 10062 4200 11154
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4066 9752 4122 9761
rect 4066 9687 4068 9696
rect 4120 9687 4122 9696
rect 4068 9658 4120 9664
rect 3700 9580 3752 9586
rect 3988 9574 4108 9602
rect 3700 9522 3752 9528
rect 4080 9450 4108 9574
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3882 9208 3938 9217
rect 3882 9143 3938 9152
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3804 8809 3832 9046
rect 3896 8906 3924 9143
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3422 3904 3478 3913
rect 3422 3839 3478 3848
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3238 1592 3294 1601
rect 3238 1527 3294 1536
rect 3436 800 3464 3674
rect 3528 3097 3556 6054
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2582 3556 2790
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3620 1193 3648 7210
rect 3712 3924 3740 8434
rect 3882 8256 3938 8265
rect 3882 8191 3938 8200
rect 3896 8090 3924 8191
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 5914 3832 7210
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3896 6458 3924 7142
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3790 5400 3846 5409
rect 3790 5335 3846 5344
rect 3804 4758 3832 5335
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3896 4457 3924 5102
rect 3882 4448 3938 4457
rect 3882 4383 3938 4392
rect 3988 4298 4016 8978
rect 4080 8498 4108 9386
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4080 8362 4108 8434
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4080 7313 4108 7958
rect 4264 7546 4292 13942
rect 4632 13926 4752 13942
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13530 4476 13670
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4724 10810 4752 13926
rect 4816 13870 4844 18022
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4908 15978 4936 16594
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4908 14006 4936 14554
rect 4896 14000 4948 14006
rect 4896 13942 4948 13948
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9602 4752 10610
rect 4816 10266 4844 13806
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4908 11370 4936 12718
rect 5000 12481 5028 15914
rect 5092 14906 5120 20046
rect 5184 16046 5212 22000
rect 5644 19718 5672 22000
rect 6104 21962 6132 22000
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5460 18612 5488 19178
rect 5552 18902 5580 19654
rect 5920 18970 5948 19858
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5816 18624 5868 18630
rect 5460 18584 5816 18612
rect 5460 17814 5488 18584
rect 5816 18566 5868 18572
rect 6012 18426 6040 19790
rect 6288 19446 6316 21898
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6092 19440 6144 19446
rect 6092 19382 6144 19388
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5276 16454 5304 17614
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5368 15978 5396 17682
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5828 16590 5856 17614
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5920 16794 5948 16934
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 6012 16726 6040 16934
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5092 14878 5212 14906
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14346 5120 14758
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5184 12986 5212 14878
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 4908 11342 5028 11370
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4724 9574 4844 9602
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 8974 4752 9454
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8498 4752 8910
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4816 8294 4844 9574
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4264 6474 4292 6802
rect 4632 6746 4660 7346
rect 4724 6934 4752 7822
rect 4816 7410 4844 8230
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4908 7290 4936 11154
rect 5000 10674 5028 11342
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 9466 5028 10474
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 9654 5120 10406
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5000 9438 5120 9466
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9178 5028 9318
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4908 7262 5028 7290
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4632 6718 4752 6746
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4172 6446 4292 6474
rect 4172 5370 4200 6446
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4068 5024 4120 5030
rect 4066 4992 4068 5001
rect 4120 4992 4122 5001
rect 4066 4927 4122 4936
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3896 4270 4016 4298
rect 3792 3936 3844 3942
rect 3712 3896 3792 3924
rect 3792 3878 3844 3884
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3712 2038 3740 3470
rect 3700 2032 3752 2038
rect 3700 1974 3752 1980
rect 3606 1184 3662 1193
rect 3606 1119 3662 1128
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3804 649 3832 3878
rect 3896 800 3924 4270
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 3988 2650 4016 3567
rect 4080 3058 4108 4558
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3790 640 3846 649
rect 3790 575 3846 584
rect 3882 0 3938 800
rect 4066 232 4122 241
rect 4172 218 4200 5170
rect 4264 1442 4292 6054
rect 4356 5642 4384 6054
rect 4632 5710 4660 6258
rect 4724 5914 4752 6718
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5234 4752 5850
rect 4816 5302 4844 7142
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 3738 4476 4082
rect 4908 4078 4936 7142
rect 5000 6118 5028 7262
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5092 5710 5120 9438
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5030 5120 5646
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4528 3936 4580 3942
rect 4526 3904 4528 3913
rect 4712 3936 4764 3942
rect 4580 3904 4582 3913
rect 4712 3878 4764 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4526 3839 4582 3848
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4724 2650 4752 3878
rect 5092 3738 5120 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3618 5212 12718
rect 5276 12102 5304 15846
rect 5552 15638 5580 16050
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5552 14958 5580 15574
rect 5644 15026 5672 15846
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5460 14618 5488 14826
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5644 14074 5672 14214
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5736 13802 5764 16118
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 14278 5948 14418
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5724 13320 5776 13326
rect 5828 13308 5856 14214
rect 5920 13938 5948 14214
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5776 13280 5856 13308
rect 5724 13262 5776 13268
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12782 5396 13126
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5460 12306 5488 12786
rect 5552 12442 5580 13262
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5736 12374 5764 13262
rect 6104 13172 6132 19382
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6196 16726 6224 17206
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 5828 13144 6132 13172
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 10674 5396 11562
rect 5460 11082 5488 12242
rect 5736 12238 5764 12310
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11218 5764 12174
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5368 10266 5396 10610
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5356 10260 5408 10266
rect 5460 10248 5488 10474
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5460 10220 5580 10248
rect 5356 10202 5408 10208
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5276 9586 5304 10066
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5262 9480 5318 9489
rect 5262 9415 5318 9424
rect 5276 8566 5304 9415
rect 5368 9178 5396 9862
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7750 5396 8230
rect 5460 8090 5488 10066
rect 5552 10062 5580 10220
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5644 9994 5672 10406
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5828 9654 5856 13144
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10606 6132 10950
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10266 6132 10406
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 6866 5304 7346
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5460 6474 5488 8026
rect 5552 7954 5580 8434
rect 5644 8430 5672 9318
rect 5736 8634 5764 9318
rect 6104 9042 6132 9522
rect 5908 9036 5960 9042
rect 6092 9036 6144 9042
rect 5960 8996 6040 9024
rect 5908 8978 5960 8984
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5828 8786 5856 8842
rect 5828 8758 5948 8786
rect 5920 8634 5948 8758
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7002 5580 7890
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5828 6746 5856 8502
rect 6012 8294 6040 8996
rect 6092 8978 6144 8984
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5920 7546 5948 8230
rect 6104 8090 6132 8978
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6196 7546 6224 11222
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 5998 6896 6054 6905
rect 6196 6866 6224 7482
rect 6288 7206 6316 11290
rect 6380 9602 6408 19654
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 13938 6500 15302
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11898 6500 12242
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6380 9574 6500 9602
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 8090 6408 9386
rect 6472 8634 6500 9574
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5998 6831 6054 6840
rect 6184 6860 6236 6866
rect 5828 6718 5948 6746
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5276 6446 5488 6474
rect 5276 5778 5304 6446
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5914 5396 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5552 5692 5580 6258
rect 5644 6254 5672 6598
rect 5828 6458 5856 6598
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5632 5704 5684 5710
rect 5552 5664 5632 5692
rect 5632 5646 5684 5652
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4146 5396 4490
rect 5644 4146 5672 4626
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 4816 3590 5212 3618
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4384 1442
rect 4356 800 4384 1414
rect 4816 800 4844 3590
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 2922 5304 3470
rect 5368 2990 5396 4082
rect 5538 3904 5594 3913
rect 5538 3839 5594 3848
rect 5552 3126 5580 3839
rect 5644 3534 5672 4082
rect 5736 3602 5764 5102
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5736 3058 5764 3538
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5356 2984 5408 2990
rect 5920 2938 5948 6718
rect 6012 6186 6040 6831
rect 6184 6802 6236 6808
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6288 5914 6316 6734
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 3194 6040 3538
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5356 2926 5408 2932
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5736 2910 5948 2938
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5276 800 5304 2450
rect 5736 800 5764 2910
rect 5908 2440 5960 2446
rect 6012 2428 6040 3130
rect 5960 2400 6040 2428
rect 5908 2382 5960 2388
rect 6196 800 6224 5782
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6380 5030 6408 5646
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6288 4078 6316 4422
rect 6380 4146 6408 4966
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6472 921 6500 7210
rect 6564 3641 6592 22000
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19310 6868 19654
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6932 18834 6960 19790
rect 7024 18902 7052 22000
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6840 18086 6868 18226
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6840 17814 6868 18022
rect 6932 17882 6960 18770
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 7116 17202 7144 20266
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 18358 7328 18566
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7288 18216 7340 18222
rect 7194 18184 7250 18193
rect 7288 18158 7340 18164
rect 7194 18119 7250 18128
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6932 16250 6960 17002
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 13870 6868 14758
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6932 12986 6960 14418
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 13870 7144 14350
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 13530 7144 13806
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 7116 12442 7144 13330
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6840 11354 6868 11494
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10470 6776 11086
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 10062 6776 10406
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9110 6684 9318
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6656 8430 6684 9046
rect 6840 8974 6868 10542
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 10266 6960 10474
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6932 8922 6960 9590
rect 7116 9518 7144 11494
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7324 6684 8230
rect 6748 8090 6776 8298
rect 6840 8294 6868 8910
rect 6932 8894 7052 8922
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6736 7336 6788 7342
rect 6656 7296 6736 7324
rect 6736 7278 6788 7284
rect 6748 6934 6776 7278
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 4826 6684 5510
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6748 4690 6776 5714
rect 6840 5030 6868 6326
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5914 6960 6054
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5574 7052 8894
rect 7208 8634 7236 18119
rect 7300 17746 7328 18158
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7484 17354 7512 22000
rect 7944 20330 7972 22000
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7300 17326 7512 17354
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7116 8514 7144 8570
rect 7116 8486 7236 8514
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 7018 7144 7210
rect 7208 7154 7236 8486
rect 7300 7274 7328 17326
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 9518 7420 17138
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7484 13258 7512 13330
rect 7576 13326 7604 19110
rect 7668 18902 7696 19246
rect 7760 18970 7788 19858
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7852 19514 7880 19790
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 8036 18630 8064 18838
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8116 18624 8168 18630
rect 8220 18612 8248 19790
rect 8168 18584 8248 18612
rect 8116 18566 8168 18572
rect 8128 18222 8156 18566
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16794 7696 16934
rect 7760 16794 7788 17478
rect 8220 17338 8248 17478
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 15978 8248 16526
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15434 8248 15914
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8312 15366 8340 15982
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14600 8248 14894
rect 8312 14822 8340 15302
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8300 14612 8352 14618
rect 8220 14572 8300 14600
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7668 13530 7696 14486
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7484 12850 7512 13194
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7576 12730 7604 13262
rect 8220 12918 8248 14572
rect 8300 14554 8352 14560
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 7484 12702 7604 12730
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7484 11694 7512 12702
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 12442 7604 12582
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7668 11558 7696 12718
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8404 12374 8432 22000
rect 8864 19802 8892 22000
rect 8772 19774 8892 19802
rect 9036 19780 9088 19786
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8496 18970 8524 19178
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8574 18864 8630 18873
rect 8574 18799 8630 18808
rect 8482 18728 8538 18737
rect 8482 18663 8538 18672
rect 8496 18290 8524 18663
rect 8588 18358 8616 18799
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8588 17649 8616 17818
rect 8772 17814 8800 19774
rect 9036 19722 9088 19728
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19310 8892 19654
rect 9048 19378 9076 19722
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9140 18222 9168 18702
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9324 18086 9352 22000
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9508 18902 9536 19246
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9508 18766 9536 18838
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8760 17672 8812 17678
rect 8574 17640 8630 17649
rect 8760 17614 8812 17620
rect 8574 17575 8630 17584
rect 8588 17338 8616 17575
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8772 17270 8800 17614
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 15706 8524 16594
rect 8588 16250 8616 17138
rect 9508 17134 9536 18702
rect 9692 17542 9720 18906
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9496 17128 9548 17134
rect 8942 17096 8998 17105
rect 9496 17070 9548 17076
rect 8942 17031 8998 17040
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8760 16516 8812 16522
rect 8760 16458 8812 16464
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8772 16046 8800 16458
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8864 15706 8892 16934
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8956 14958 8984 17031
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9324 16794 9352 16934
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9508 16522 9536 17070
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9692 15026 9720 16662
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 9416 14906 9444 14962
rect 9784 14906 9812 22000
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 19242 9904 19790
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 18970 9904 19178
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10152 18426 10180 19858
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9862 17776 9918 17785
rect 9862 17711 9918 17720
rect 9876 15706 9904 17711
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9416 14878 9812 14906
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8496 14074 8524 14486
rect 8680 14482 8708 14758
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8680 13870 8708 14418
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13530 9168 13738
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 8392 12368 8444 12374
rect 8576 12368 8628 12374
rect 8392 12310 8444 12316
rect 8496 12316 8576 12322
rect 8496 12310 8628 12316
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11898 8064 12174
rect 8312 11898 8340 12242
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8404 11778 8432 12310
rect 8496 12294 8616 12310
rect 8496 12238 8524 12294
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 8312 11750 8432 11778
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7760 11014 7788 11698
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7392 8498 7420 9114
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7208 7126 7328 7154
rect 7116 6990 7236 7018
rect 7208 6662 7236 6990
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 5710 7236 6598
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 3670 6776 4626
rect 6932 4622 6960 5034
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6736 3664 6788 3670
rect 6550 3632 6606 3641
rect 6736 3606 6788 3612
rect 6550 3567 6606 3576
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6458 912 6514 921
rect 6458 847 6514 856
rect 6656 800 6684 3130
rect 6748 1902 6776 3606
rect 6840 3602 6868 4558
rect 6932 4214 6960 4558
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 2106 6960 3470
rect 7208 2582 7236 4422
rect 7300 4185 7328 7126
rect 7392 5794 7420 8434
rect 7484 8090 7512 10950
rect 8220 10810 8248 11086
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7576 9722 7604 9998
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9110 7788 9522
rect 8220 9450 8248 9998
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 9178 8248 9386
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7484 5914 7512 6190
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7392 5766 7512 5794
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4758 7420 4966
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7286 4176 7342 4185
rect 7286 4111 7342 4120
rect 7300 4078 7328 4111
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 2990 7420 3334
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 6920 2100 6972 2106
rect 6920 2042 6972 2048
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 7102 912 7158 921
rect 7484 898 7512 5766
rect 7576 3738 7604 6190
rect 7668 6118 7696 7686
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 6866 8248 7822
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6322 8248 6802
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 4049 7696 6054
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8116 5840 8168 5846
rect 8114 5808 8116 5817
rect 8168 5808 8170 5817
rect 8114 5743 8170 5752
rect 8220 5710 8248 6258
rect 8312 6118 8340 11750
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8312 5642 8340 6054
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7840 4208 7892 4214
rect 7840 4150 7892 4156
rect 7654 4040 7710 4049
rect 7654 3975 7710 3984
rect 7852 3924 7880 4150
rect 7760 3896 7880 3924
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7760 3534 7788 3896
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 2650 7604 3334
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8116 2916 8168 2922
rect 8220 2904 8248 2994
rect 8168 2876 8248 2904
rect 8116 2858 8168 2864
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 2650 8248 2876
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8312 2446 8340 2790
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8404 2292 8432 9318
rect 8496 7478 8524 12174
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11286 8708 11494
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8588 10606 8616 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8588 10062 8616 10542
rect 8772 10266 8800 10950
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8680 8430 8708 8910
rect 8772 8430 8800 9454
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 7546 8800 8230
rect 8956 8090 8984 12174
rect 9140 11762 9168 13466
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8944 7812 8996 7818
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8496 3074 8524 7414
rect 8864 7342 8892 7783
rect 8944 7754 8996 7760
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8956 6866 8984 7754
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8864 6322 8892 6802
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8588 3194 8616 6151
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5098 8708 5510
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8772 4282 8800 4626
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 3738 8892 4558
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 4049 8984 4082
rect 8942 4040 8998 4049
rect 8942 3975 8998 3984
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8496 3046 8616 3074
rect 8128 2264 8432 2292
rect 7484 870 7604 898
rect 7102 847 7158 856
rect 7116 800 7144 847
rect 7576 800 7604 870
rect 8128 800 8156 2264
rect 8588 800 8616 3046
rect 8680 2990 8708 3130
rect 8772 3126 8800 3402
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8680 2514 8708 2926
rect 8772 2854 8800 3062
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8668 2508 8720 2514
rect 8668 2450 8720 2456
rect 8956 1970 8984 3402
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 9048 800 9076 10066
rect 9140 7886 9168 11698
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11354 9260 11494
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9416 8922 9444 14878
rect 9876 14600 9904 15506
rect 9968 14618 9996 18022
rect 10060 17814 10088 18294
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10244 16776 10272 22000
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10336 18630 10364 18770
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18290 10364 18566
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10152 16748 10272 16776
rect 10152 15706 10180 16748
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10244 16182 10272 16594
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10060 15473 10088 15506
rect 10046 15464 10102 15473
rect 10046 15399 10102 15408
rect 10152 15366 10180 15642
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 9692 14572 9904 14600
rect 9956 14612 10008 14618
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13326 9628 13670
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9600 12850 9628 13262
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9692 12764 9720 14572
rect 9956 14554 10008 14560
rect 10046 14512 10102 14521
rect 10046 14447 10048 14456
rect 10100 14447 10102 14456
rect 10048 14418 10100 14424
rect 10060 14226 10088 14418
rect 9876 14198 10088 14226
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 12918 9812 13670
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9692 12736 9812 12764
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9692 11082 9720 11766
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 9518 9720 10678
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9232 8894 9444 8922
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6934 9168 7278
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 6254 9168 6666
rect 9232 6474 9260 8894
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 6730 9352 8366
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9232 6446 9352 6474
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5710 9168 6190
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 3602 9168 5646
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9232 4146 9260 4626
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9140 2990 9168 3538
rect 9232 3534 9260 4082
rect 9324 3942 9352 6446
rect 9416 4758 9444 8774
rect 9692 7818 9720 9454
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7410 9720 7754
rect 9784 7750 9812 12736
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9586 6352 9642 6361
rect 9586 6287 9642 6296
rect 9600 6118 9628 6287
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9770 5808 9826 5817
rect 9770 5743 9772 5752
rect 9824 5743 9826 5752
rect 9772 5714 9824 5720
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9416 4010 9444 4694
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4214 9628 4558
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9232 2854 9260 3470
rect 9324 2961 9352 3878
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9310 2952 9366 2961
rect 9310 2887 9366 2896
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2446 9260 2790
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9508 800 9536 3674
rect 9600 3466 9628 4150
rect 9692 4078 9720 4966
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4146 9812 4422
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9876 3890 9904 14198
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9968 13394 9996 14010
rect 10152 14006 10180 14826
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10232 13728 10284 13734
rect 10336 13716 10364 18022
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10520 16250 10548 16934
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10612 15858 10640 18294
rect 10704 18154 10732 22000
rect 11164 18170 11192 22000
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 11072 18142 11192 18170
rect 11624 18154 11652 22000
rect 11992 19242 12020 22000
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11980 19236 12032 19242
rect 11980 19178 12032 19184
rect 11612 18148 11664 18154
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17746 10824 18022
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10520 15830 10640 15858
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10284 13688 10364 13716
rect 10232 13670 10284 13676
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 13274 9996 13330
rect 9968 13246 10088 13274
rect 10060 12238 10088 13246
rect 10140 12776 10192 12782
rect 10192 12736 10272 12764
rect 10140 12718 10192 12724
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9968 10674 9996 11698
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10810 10088 11154
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9968 10470 9996 10610
rect 10152 10577 10180 12582
rect 10244 12238 10272 12736
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10336 11694 10364 13398
rect 10428 12442 10456 14758
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10138 10568 10194 10577
rect 10138 10503 10194 10512
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9956 9512 10008 9518
rect 9954 9480 9956 9489
rect 10008 9480 10010 9489
rect 9954 9415 10010 9424
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9968 4826 9996 8978
rect 10152 8430 10180 9522
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7290 10088 7890
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7478 10180 7822
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10060 7262 10180 7290
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10060 7002 10088 7142
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10152 6798 10180 7262
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 10060 5846 10088 6015
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10152 5370 10180 6734
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10060 4690 10088 5238
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9784 3862 9904 3890
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9784 3738 9812 3862
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9600 2922 9628 3402
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9692 2582 9720 3606
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9876 1306 9904 3674
rect 9968 2650 9996 3878
rect 10060 3534 10088 3878
rect 10244 3738 10272 10746
rect 10428 10538 10456 12242
rect 10520 11286 10548 15830
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10612 13462 10640 14486
rect 10704 13546 10732 15506
rect 10796 14550 10824 17478
rect 11072 17184 11100 18142
rect 11612 18090 11664 18096
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10980 17156 11100 17184
rect 10980 16674 11008 17156
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16794 11100 17002
rect 11164 16794 11192 18022
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11808 17338 11836 17750
rect 11796 17332 11848 17338
rect 11900 17320 11928 19178
rect 12176 18358 12204 19314
rect 12452 19174 12480 22000
rect 12912 20058 12940 22000
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12636 19310 12664 19858
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12164 18352 12216 18358
rect 12070 18320 12126 18329
rect 12164 18294 12216 18300
rect 12070 18255 12126 18264
rect 11900 17292 12020 17320
rect 11796 17274 11848 17280
rect 11808 17218 11836 17274
rect 11808 17190 11928 17218
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10980 16646 11100 16674
rect 11716 16658 11744 16934
rect 11808 16794 11836 17070
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11072 16454 11100 16646
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11900 16590 11928 17190
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10874 16008 10930 16017
rect 10874 15943 10876 15952
rect 10928 15943 10930 15952
rect 10876 15914 10928 15920
rect 11072 15910 11100 16390
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11716 15706 11744 16458
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13734 10824 14214
rect 10888 13938 10916 14282
rect 10980 14074 11008 14962
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10704 13518 10916 13546
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10612 12889 10640 12922
rect 10598 12880 10654 12889
rect 10598 12815 10654 12824
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10600 12368 10652 12374
rect 10598 12336 10600 12345
rect 10652 12336 10654 12345
rect 10598 12271 10654 12280
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10428 10130 10456 10474
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10520 9518 10548 11018
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8566 10364 8842
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10336 6798 10364 7346
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 5778 10364 6734
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10152 2650 10180 3538
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3194 10272 3470
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9876 1278 9996 1306
rect 9968 800 9996 1278
rect 10428 800 10456 7686
rect 10520 6338 10548 9454
rect 10612 9382 10640 10406
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10704 7562 10732 12650
rect 10782 12608 10838 12617
rect 10782 12543 10838 12552
rect 10796 12306 10824 12543
rect 10888 12442 10916 13518
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12850 11008 13126
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10784 11756 10836 11762
rect 10888 11744 10916 12378
rect 10836 11716 10916 11744
rect 10968 11756 11020 11762
rect 10784 11698 10836 11704
rect 10968 11698 11020 11704
rect 10980 10742 11008 11698
rect 11072 11665 11100 14554
rect 11164 13258 11192 14758
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 14006 11652 14894
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11440 13462 11468 13670
rect 11716 13530 11744 14214
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11532 13326 11560 13466
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11164 12617 11192 12650
rect 11244 12640 11296 12646
rect 11150 12608 11206 12617
rect 11244 12582 11296 12588
rect 11150 12543 11206 12552
rect 11256 12374 11284 12582
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11624 11898 11652 12922
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11354 11100 11494
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 11072 10130 11100 11290
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10796 10010 10824 10066
rect 10796 9982 11100 10010
rect 11072 9586 11100 9982
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9178 10916 9318
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11072 8974 11100 9522
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11164 8498 11192 11766
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11082 11376 11494
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 9926 11652 10950
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11624 8362 11652 9454
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10704 7534 10916 7562
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10796 6390 10824 6802
rect 10784 6384 10836 6390
rect 10520 6310 10732 6338
rect 10784 6326 10836 6332
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10520 5234 10548 6054
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10612 5166 10640 6054
rect 10704 5302 10732 6310
rect 10782 5672 10838 5681
rect 10782 5607 10838 5616
rect 10796 5574 10824 5607
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10520 2553 10548 5034
rect 10796 4049 10824 5238
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10796 2582 10824 3878
rect 10784 2576 10836 2582
rect 10506 2544 10562 2553
rect 10784 2518 10836 2524
rect 10506 2479 10562 2488
rect 10888 800 10916 7534
rect 10980 7342 11008 8230
rect 11164 7886 11192 8298
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 8090 11376 8230
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11716 7954 11744 12786
rect 11808 12646 11836 15506
rect 11900 13734 11928 15642
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 12986 11928 13670
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11992 12288 12020 17292
rect 12084 15570 12112 18255
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12268 15502 12296 18158
rect 12360 17542 12388 18770
rect 12544 18290 12572 18838
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 17882 12572 18226
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17218 12388 17478
rect 12360 17190 12480 17218
rect 12348 17060 12400 17066
rect 12348 17002 12400 17008
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11900 12260 12020 12288
rect 11900 12102 11928 12260
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 6322 11008 6598
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11072 6254 11100 7482
rect 11164 7274 11192 7822
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11164 6730 11192 7210
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10980 5914 11008 6122
rect 11164 6118 11192 6394
rect 11716 6254 11744 7890
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10980 5234 11008 5850
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11072 4826 11100 5646
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5166 11192 5510
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11624 4690 11652 6054
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5302 11744 5714
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11704 5024 11756 5030
rect 11808 5012 11836 11834
rect 11886 11792 11942 11801
rect 11886 11727 11942 11736
rect 11900 11694 11928 11727
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11992 11354 12020 12106
rect 12084 11898 12112 15302
rect 12268 15042 12296 15438
rect 12176 15014 12296 15042
rect 12176 14550 12204 15014
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 13938 12204 14350
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 12850 12204 13874
rect 12268 13530 12296 14826
rect 12360 14618 12388 17002
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 14006 12480 17190
rect 12636 14618 12664 18906
rect 12728 18902 12756 19246
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12820 18766 12848 19178
rect 13280 18970 13308 19926
rect 13372 19174 13400 22000
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13648 18834 13676 19858
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17882 12848 18022
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12912 17746 12940 18158
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 13096 17814 13124 18090
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12452 13530 12480 13942
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12256 12776 12308 12782
rect 12360 12753 12388 13194
rect 12256 12718 12308 12724
rect 12346 12744 12402 12753
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12176 11830 12204 12582
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11992 9926 12020 10610
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 12084 9586 12112 11698
rect 12176 11218 12204 11766
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12162 11112 12218 11121
rect 12162 11047 12218 11056
rect 12176 10538 12204 11047
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 9042 12020 9318
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 6934 12112 7142
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 5840 11940 5846
rect 11886 5808 11888 5817
rect 11940 5808 11942 5817
rect 11886 5743 11942 5752
rect 11992 5114 12020 6258
rect 12084 5234 12112 6870
rect 12176 6746 12204 10474
rect 12268 10266 12296 12718
rect 12452 12714 12480 13466
rect 12544 13462 12572 13670
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12530 12744 12586 12753
rect 12346 12679 12402 12688
rect 12440 12708 12492 12714
rect 12530 12679 12532 12688
rect 12440 12650 12492 12656
rect 12584 12679 12586 12688
rect 12532 12650 12584 12656
rect 12636 12220 12664 14554
rect 12728 14521 12756 17478
rect 12912 17105 12940 17682
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12898 17096 12954 17105
rect 12898 17031 12954 17040
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 15706 12940 16934
rect 13004 16046 13032 17138
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13082 15464 13138 15473
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12820 14890 12848 15030
rect 13004 15026 13032 15438
rect 13082 15399 13138 15408
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12808 14884 12860 14890
rect 12860 14844 12940 14872
rect 12808 14826 12860 14832
rect 12714 14512 12770 14521
rect 12714 14447 12770 14456
rect 12728 13394 12756 14447
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12820 12986 12848 13806
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12912 12866 12940 14844
rect 13004 14414 13032 14962
rect 13096 14414 13124 15399
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13188 13530 13216 13942
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12820 12838 12940 12866
rect 12820 12458 12848 12838
rect 12811 12442 12848 12458
rect 12808 12436 12860 12442
rect 12544 12192 12664 12220
rect 12728 12396 12808 12424
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11354 12388 12038
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12268 8430 12296 10202
rect 12452 10130 12480 11698
rect 12544 11626 12572 12192
rect 12728 12152 12756 12396
rect 12808 12378 12860 12384
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12636 12124 12756 12152
rect 12636 11801 12664 12124
rect 12622 11792 12678 11801
rect 12622 11727 12678 11736
rect 12714 11656 12770 11665
rect 12532 11620 12584 11626
rect 12820 11626 12848 12174
rect 12714 11591 12770 11600
rect 12808 11620 12860 11626
rect 12532 11562 12584 11568
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12360 9489 12388 9930
rect 12544 9738 12572 11222
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10266 12664 10406
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12452 9710 12572 9738
rect 12452 9654 12480 9710
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12728 9568 12756 11591
rect 12808 11562 12860 11568
rect 12820 11150 12848 11562
rect 13004 11354 13032 12174
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11354 13308 11494
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12912 10674 12940 11018
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 9636 12848 10406
rect 12719 9540 12756 9568
rect 12811 9608 12848 9636
rect 12719 9500 12747 9540
rect 12811 9500 12839 9608
rect 12346 9480 12402 9489
rect 12719 9472 12756 9500
rect 12811 9472 12848 9500
rect 12346 9415 12348 9424
rect 12400 9415 12402 9424
rect 12348 9386 12400 9392
rect 12360 8974 12388 9386
rect 12728 9058 12756 9472
rect 12820 9178 12848 9472
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12532 9036 12584 9042
rect 12728 9030 12848 9058
rect 12532 8978 12584 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12544 8362 12572 8978
rect 12716 8968 12768 8974
rect 12714 8936 12716 8945
rect 12768 8936 12770 8945
rect 12714 8871 12770 8880
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8022 12664 8230
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7342 12664 7958
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12728 7188 12756 8871
rect 12636 7160 12756 7188
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12440 6792 12492 6798
rect 12176 6718 12296 6746
rect 12440 6734 12492 6740
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 5710 12204 6598
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12176 5166 12204 5646
rect 12164 5160 12216 5166
rect 11992 5086 12112 5114
rect 12164 5102 12216 5108
rect 11808 4984 12020 5012
rect 11704 4966 11756 4972
rect 11716 4826 11744 4966
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 4146 11008 4490
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11072 3194 11100 4558
rect 11164 4214 11192 4626
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11256 3670 11284 4082
rect 11244 3664 11296 3670
rect 11164 3624 11244 3652
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11072 2854 11100 2994
rect 11164 2922 11192 3624
rect 11244 3606 11296 3612
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 2446 11100 2790
rect 11164 2446 11192 2858
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2553 11376 2790
rect 11716 2650 11744 4082
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11334 2544 11390 2553
rect 11334 2479 11390 2488
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11334 2000 11390 2009
rect 11334 1935 11390 1944
rect 11348 800 11376 1935
rect 11808 800 11836 4422
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 2650 11928 3334
rect 11992 2922 12020 4984
rect 12084 4690 12112 5086
rect 12268 4808 12296 6718
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12360 5352 12388 6326
rect 12452 5914 12480 6734
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12360 5324 12480 5352
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12176 4780 12296 4808
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12084 4282 12112 4626
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12176 4026 12204 4780
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12268 4146 12296 4626
rect 12360 4622 12388 5170
rect 12452 4826 12480 5324
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12544 4026 12572 6870
rect 12636 4486 12664 7160
rect 12820 6610 12848 9030
rect 12728 6582 12848 6610
rect 12728 5012 12756 6582
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12820 5166 12848 5646
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12912 5098 12940 10503
rect 13004 9636 13032 10610
rect 13004 9625 13124 9636
rect 13280 9625 13308 11154
rect 13004 9616 13138 9625
rect 13004 9608 13082 9616
rect 13082 9551 13138 9560
rect 13266 9616 13322 9625
rect 13266 9551 13322 9560
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 8974 13124 9454
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13372 6746 13400 13738
rect 13464 11121 13492 18770
rect 13832 18426 13860 22000
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17882 13860 18090
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13648 15994 13676 17750
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13740 16726 13768 17002
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 16130 13768 16390
rect 13832 16250 13860 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13924 16130 13952 17070
rect 13740 16102 13952 16130
rect 13820 16040 13872 16046
rect 13648 15966 13768 15994
rect 13820 15982 13872 15988
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 15094 13676 15506
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13740 15042 13768 15966
rect 13832 15162 13860 15982
rect 13924 15978 13952 16102
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13924 15366 13952 15914
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13740 15014 13860 15042
rect 13832 13818 13860 15014
rect 13924 14006 13952 15302
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13832 13790 13952 13818
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13556 11898 13584 12310
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 11286 13584 11562
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13544 11144 13596 11150
rect 13450 11112 13506 11121
rect 13544 11086 13596 11092
rect 13450 11047 13506 11056
rect 13556 10674 13584 11086
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10198 13584 10406
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13556 9364 13584 10134
rect 13464 9336 13584 9364
rect 13464 7002 13492 9336
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 8430 13584 8910
rect 13648 8498 13676 12815
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13740 12170 13768 12650
rect 13832 12442 13860 12650
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11898 13768 12106
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10826 13860 11086
rect 13740 10798 13860 10826
rect 13740 10470 13768 10798
rect 13924 10690 13952 13790
rect 14016 13462 14044 18838
rect 14108 15706 14136 19246
rect 14292 19174 14320 22000
rect 14752 20346 14780 22000
rect 14568 20318 14780 20346
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14108 15026 14136 15506
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14200 14770 14228 18838
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14292 16250 14320 17614
rect 14384 17134 14412 17614
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16794 14412 17070
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14476 15994 14504 19246
rect 14568 18970 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 15120 18902 15148 19246
rect 15212 19174 15240 22000
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15108 18896 15160 18902
rect 15108 18838 15160 18844
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15016 18216 15068 18222
rect 15016 18158 15068 18164
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14476 15966 14596 15994
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 14816 14332 14822
rect 14108 14764 14280 14770
rect 14108 14758 14332 14764
rect 14108 14742 14320 14758
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14108 12866 14136 14742
rect 14384 14600 14412 15642
rect 14476 15638 14504 15846
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14568 15484 14596 15966
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14200 14572 14412 14600
rect 14476 15456 14596 15484
rect 14200 13802 14228 14572
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14200 12986 14228 13330
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14108 12838 14228 12866
rect 14200 11268 14228 12838
rect 14292 12374 14320 13942
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14384 11778 14412 14418
rect 14292 11750 14412 11778
rect 14292 11336 14320 11750
rect 14476 11642 14504 15456
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14414 14596 14962
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14568 12986 14596 13398
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 11898 14596 12582
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14384 11626 14504 11642
rect 14372 11620 14504 11626
rect 14424 11614 14504 11620
rect 14648 11620 14700 11626
rect 14372 11562 14424 11568
rect 14568 11580 14648 11608
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11354 14504 11494
rect 14464 11348 14516 11354
rect 14292 11308 14412 11336
rect 14200 11240 14320 11268
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13832 10662 13952 10690
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13832 10248 13860 10662
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13740 10220 13860 10248
rect 13740 9466 13768 10220
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9654 13860 10066
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13740 9438 13860 9466
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 7936 13584 8366
rect 13636 7948 13688 7954
rect 13556 7908 13636 7936
rect 13636 7890 13688 7896
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7206 13584 7686
rect 13648 7410 13676 7890
rect 13832 7478 13860 9438
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13280 6718 13400 6746
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12808 5024 12860 5030
rect 12728 4984 12808 5012
rect 12808 4966 12860 4972
rect 12716 4752 12768 4758
rect 12820 4729 12848 4966
rect 13280 4758 13308 6718
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6254 13400 6598
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13556 5166 13584 7142
rect 13648 6202 13676 7346
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6322 13768 6734
rect 13924 6730 13952 10542
rect 14016 10266 14044 11154
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14200 10674 14228 11086
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14292 9602 14320 11240
rect 14384 11234 14412 11308
rect 14464 11290 14516 11296
rect 14384 11206 14504 11234
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14016 9574 14320 9602
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13648 6174 13768 6202
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13268 4752 13320 4758
rect 12716 4694 12768 4700
rect 12806 4720 12862 4729
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12176 3998 12296 4026
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 3194 12112 3470
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11900 2310 11928 2450
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12268 800 12296 3998
rect 12452 3998 12572 4026
rect 12452 3942 12480 3998
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12530 3224 12586 3233
rect 12530 3159 12586 3168
rect 12544 3126 12572 3159
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12438 2952 12494 2961
rect 12438 2887 12494 2896
rect 12452 2854 12480 2887
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12636 2514 12664 3334
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12728 800 12756 4694
rect 13268 4694 13320 4700
rect 12806 4655 12862 4664
rect 13556 4622 13584 5102
rect 13740 5030 13768 6174
rect 14016 5914 14044 9574
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 6662 14136 8978
rect 14200 8906 14228 9318
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14292 8566 14320 9454
rect 14384 9178 14412 9658
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14476 9058 14504 11206
rect 14568 10810 14596 11580
rect 14648 11562 14700 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14568 9586 14596 10474
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 15028 9450 15056 18158
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15120 16046 15148 17274
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15212 15706 15240 16050
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15304 14822 15332 18362
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14362 15332 14758
rect 15396 14482 15424 14894
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15108 14340 15160 14346
rect 15304 14334 15424 14362
rect 15108 14282 15160 14288
rect 15120 13258 15148 14282
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15212 13274 15240 14010
rect 15304 13530 15332 14214
rect 15396 13734 15424 14334
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15396 13462 15424 13670
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15108 13252 15160 13258
rect 15212 13246 15332 13274
rect 15108 13194 15160 13200
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15120 11762 15148 12310
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15212 10418 15240 12718
rect 15304 10674 15332 13246
rect 15488 11286 15516 19246
rect 15672 19174 15700 22000
rect 16132 19174 16160 22000
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 15042 15608 16526
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15672 15162 15700 15914
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15580 15014 15700 15042
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14618 15608 14758
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15672 14498 15700 15014
rect 15580 14470 15700 14498
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15384 10464 15436 10470
rect 15212 10412 15384 10418
rect 15212 10406 15436 10412
rect 15120 10266 15148 10406
rect 15212 10390 15424 10406
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14384 9042 14504 9058
rect 14372 9036 14504 9042
rect 14424 9030 14504 9036
rect 14372 8978 14424 8984
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14292 6118 14320 8502
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14384 8090 14412 8298
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14568 7886 14596 8298
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 8090 15056 8570
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 7002 14504 7142
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6882 14596 7822
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14844 7342 14872 7414
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14568 6854 14688 6882
rect 14660 6798 14688 6854
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 15212 6662 15240 9318
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 14476 6322 14504 6598
rect 15304 6322 15332 10390
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15396 8430 15424 10066
rect 15384 8424 15436 8430
rect 15580 8378 15608 14470
rect 15764 12986 15792 15438
rect 15856 14414 15884 16934
rect 15948 16130 15976 18634
rect 16040 18290 16068 18770
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16132 16250 16160 17682
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 15948 16102 16160 16130
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15948 15026 15976 15438
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 13870 15884 14350
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15856 12782 15884 12815
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15672 11354 15700 11630
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15764 9722 15792 12650
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15384 8366 15436 8372
rect 15396 7342 15424 8366
rect 15488 8350 15608 8378
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 14280 6112 14332 6118
rect 14476 6089 14504 6258
rect 14280 6054 14332 6060
rect 14462 6080 14518 6089
rect 14462 6015 14518 6024
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 15120 5778 15148 6258
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 5574 15148 5714
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12898 4176 12954 4185
rect 12898 4111 12954 4120
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12820 2990 12848 3402
rect 12912 3398 12940 4111
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13004 3233 13032 3878
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12990 3224 13046 3233
rect 12990 3159 13046 3168
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 13096 2378 13124 3470
rect 13372 2514 13400 3946
rect 13464 2582 13492 4014
rect 13556 2990 13584 4558
rect 13740 4214 13768 4966
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13832 2378 13860 5034
rect 14016 3738 14044 5238
rect 14200 4758 14228 5510
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14188 4752 14240 4758
rect 15028 4706 15056 5034
rect 14188 4694 14240 4700
rect 14936 4678 15056 4706
rect 14936 4486 14964 4678
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 15120 4146 15148 5510
rect 15212 4826 15240 6054
rect 15396 5710 15424 7278
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 5166 15424 5646
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14568 3942 14596 4082
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13188 800 13216 2246
rect 13648 800 13676 2246
rect 14108 800 14136 3878
rect 14568 3670 14596 3878
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 15120 3602 15148 4082
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15212 3738 15240 3878
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14476 2922 14504 3402
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14568 800 14596 2586
rect 15028 800 15056 2858
rect 15120 2854 15148 3538
rect 15304 3534 15332 3878
rect 15488 3670 15516 8350
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 7342 15608 8230
rect 15764 8090 15792 8774
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15580 6866 15608 7278
rect 15672 7002 15700 7686
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15856 6746 15884 11154
rect 15948 11150 15976 13262
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12850 16068 13194
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10674 15976 11086
rect 16132 10742 16160 16102
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10198 15976 10610
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15948 9586 15976 10134
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 16224 9110 16252 19246
rect 16592 18970 16620 22000
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16684 18902 16712 19654
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 11354 16344 18702
rect 16408 17542 16436 18770
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 15706 16528 15846
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16868 15314 16896 18090
rect 16960 15858 16988 19246
rect 17052 19242 17080 22000
rect 17512 19428 17540 22000
rect 17420 19400 17540 19428
rect 17224 19304 17276 19310
rect 17144 19264 17224 19292
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16960 15830 17080 15858
rect 16868 15286 16988 15314
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 13326 16436 13670
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11626 16896 12038
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 11354 16804 11494
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16684 10810 16712 11154
rect 16868 11150 16896 11562
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16960 11014 16988 15286
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 9654 16344 10406
rect 16684 10266 16712 10610
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 15580 6718 15884 6746
rect 15580 6225 15608 6718
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15566 6216 15622 6225
rect 15566 6151 15622 6160
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15580 800 15608 3062
rect 15672 2990 15700 6598
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15764 4826 15792 6394
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15856 5574 15884 6258
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15948 5681 15976 5782
rect 15934 5672 15990 5681
rect 15934 5607 15990 5616
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5166 15976 5510
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4826 16436 4966
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 16684 4570 16712 7210
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16776 4690 16804 6054
rect 16868 5030 16896 10678
rect 17052 10130 17080 15830
rect 17144 12345 17172 19264
rect 17224 19246 17276 19252
rect 17420 19174 17448 19400
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17512 18290 17540 19246
rect 17972 19174 18000 22000
rect 18432 19802 18460 22000
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18432 19774 18552 19802
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19174 18552 19774
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 18420 18216 18472 18222
rect 18418 18184 18420 18193
rect 18472 18184 18474 18193
rect 18418 18119 18474 18128
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17958 17232 18014 17241
rect 17958 17167 18014 17176
rect 17972 17066 18000 17167
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 16017 17448 16390
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17406 16008 17462 16017
rect 17406 15943 17462 15952
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17130 12336 17186 12345
rect 17130 12271 17186 12280
rect 17236 11694 17264 13126
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11762 17356 12242
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17328 10674 17356 11698
rect 17420 11082 17448 15943
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18616 14074 18644 19858
rect 18892 18970 18920 22000
rect 19352 20058 19380 22000
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18984 14346 19012 18770
rect 19352 18290 19380 19858
rect 19812 18970 19840 22000
rect 20272 20058 20300 22000
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 20364 16454 20392 19246
rect 20732 19174 20760 22000
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 21192 18358 21220 22000
rect 21652 18902 21680 22000
rect 22112 19242 22140 22000
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 22572 18426 22600 22000
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6866 17080 7142
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5098 16988 6054
rect 17052 5778 17080 6802
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17144 5778 17172 6258
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17052 5234 17080 5714
rect 17144 5574 17172 5714
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 15856 4214 15884 4558
rect 16684 4542 16804 4570
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 16684 4010 16712 4422
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 15750 3632 15806 3641
rect 15750 3567 15752 3576
rect 15804 3567 15806 3576
rect 15752 3538 15804 3544
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 2990 15976 3334
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16316 2582 16344 3878
rect 16776 3602 16804 4542
rect 16764 3596 16816 3602
rect 16868 3584 16896 4966
rect 17144 4622 17172 5510
rect 17236 5166 17264 8298
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17314 6352 17370 6361
rect 17314 6287 17370 6296
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16948 3596 17000 3602
rect 16868 3556 16948 3584
rect 16764 3538 16816 3544
rect 16948 3538 17000 3544
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 16040 800 16068 2314
rect 16500 800 16528 3334
rect 17328 2990 17356 6287
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16684 2650 16712 2790
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16960 800 16988 2790
rect 17130 2544 17186 2553
rect 17696 2514 17724 7210
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 5574 17908 5714
rect 18892 5710 18920 6734
rect 19168 5817 19196 6802
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6390 20300 6598
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19154 5808 19210 5817
rect 19154 5743 19210 5752
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 4434 17908 5102
rect 17972 4622 18000 5510
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 19812 5166 19840 6122
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 18878 4720 18934 4729
rect 18878 4655 18934 4664
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 17880 4406 18000 4434
rect 17972 2514 18000 4406
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18524 4078 18552 4558
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 17130 2479 17132 2488
rect 17184 2479 17186 2488
rect 17684 2508 17736 2514
rect 17132 2450 17184 2456
rect 17684 2450 17736 2456
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17420 800 17448 2246
rect 17972 1442 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18524 1442 18552 2790
rect 17880 1414 18000 1442
rect 18340 1414 18552 1442
rect 17880 800 17908 1414
rect 18340 800 18368 1414
rect 18800 800 18828 3878
rect 18892 2514 18920 4655
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19444 2514 19472 3130
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 800 19288 2246
rect 19720 800 19748 2790
rect 20272 2514 20300 3470
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 800 20208 2246
rect 20640 800 20668 4966
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21100 800 21128 2246
rect 21560 800 21588 3402
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 800 22048 3334
rect 22480 800 22508 3674
rect 4122 190 4200 218
rect 4066 167 4122 176
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
<< via2 >>
rect 3514 22072 3570 22128
rect 202 17040 258 17096
rect 1950 19216 2006 19272
rect 1950 18828 2006 18864
rect 1950 18808 1952 18828
rect 1952 18808 2004 18828
rect 2004 18808 2006 18828
rect 1674 18692 1730 18728
rect 1674 18672 1676 18692
rect 1676 18672 1728 18692
rect 1728 18672 1730 18692
rect 2134 18672 2190 18728
rect 1490 18264 1546 18320
rect 2778 20168 2834 20224
rect 3054 21120 3110 21176
rect 1674 17720 1730 17776
rect 1582 17312 1638 17368
rect 2410 18128 2466 18184
rect 3330 20576 3386 20632
rect 3422 19624 3478 19680
rect 2502 17720 2558 17776
rect 1674 16360 1730 16416
rect 3054 16768 3110 16824
rect 1766 15816 1822 15872
rect 1674 15408 1730 15464
rect 4066 22480 4122 22536
rect 3606 21528 3662 21584
rect 3790 17584 3846 17640
rect 2778 14456 2834 14512
rect 1582 13504 1638 13560
rect 2778 13912 2834 13968
rect 3238 14864 3294 14920
rect 1766 2488 1822 2544
rect 3238 6296 3294 6352
rect 2870 2080 2926 2136
rect 3146 3440 3202 3496
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4066 12960 4122 13016
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3882 12552 3938 12608
rect 3974 12416 4030 12472
rect 4066 12008 4122 12064
rect 3882 11600 3938 11656
rect 4066 11056 4122 11112
rect 4066 10648 4122 10704
rect 4066 10140 4068 10160
rect 4068 10140 4120 10160
rect 4120 10140 4122 10160
rect 4066 10104 4122 10140
rect 4066 9716 4122 9752
rect 4066 9696 4068 9716
rect 4068 9696 4120 9716
rect 4120 9696 4122 9716
rect 3882 9152 3938 9208
rect 3790 8744 3846 8800
rect 3422 3848 3478 3904
rect 3238 1536 3294 1592
rect 3514 3032 3570 3088
rect 3882 8200 3938 8256
rect 3790 5344 3846 5400
rect 3882 4392 3938 4448
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4986 12416 5042 12472
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4066 7248 4122 7304
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 4972 4068 4992
rect 4068 4972 4120 4992
rect 4120 4972 4122 4992
rect 4066 4936 4122 4972
rect 3606 1128 3662 1184
rect 3974 3576 4030 3632
rect 3790 584 3846 640
rect 4066 176 4122 232
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4526 3884 4528 3904
rect 4528 3884 4580 3904
rect 4580 3884 4582 3904
rect 4526 3848 4582 3884
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 5262 9424 5318 9480
rect 5998 6840 6054 6896
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5538 3848 5594 3904
rect 7194 18128 7250 18184
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8574 18808 8630 18864
rect 8482 18672 8538 18728
rect 8574 17584 8630 17640
rect 8942 17040 8998 17096
rect 9862 17720 9918 17776
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 6550 3576 6606 3632
rect 6458 856 6514 912
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7286 4120 7342 4176
rect 7102 856 7158 912
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8114 5788 8116 5808
rect 8116 5788 8168 5808
rect 8168 5788 8170 5808
rect 8114 5752 8170 5788
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7654 3984 7710 4040
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8850 7792 8906 7848
rect 8574 6160 8630 6216
rect 8942 3984 8998 4040
rect 10046 15408 10102 15464
rect 10046 14476 10102 14512
rect 10046 14456 10048 14476
rect 10048 14456 10100 14476
rect 10100 14456 10102 14476
rect 9586 6296 9642 6352
rect 9770 5772 9826 5808
rect 9770 5752 9772 5772
rect 9772 5752 9824 5772
rect 9824 5752 9826 5772
rect 9310 2896 9366 2952
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 10138 10512 10194 10568
rect 9954 9460 9956 9480
rect 9956 9460 10008 9480
rect 10008 9460 10010 9480
rect 9954 9424 10010 9460
rect 10046 6024 10102 6080
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 12070 18264 12126 18320
rect 10874 15972 10930 16008
rect 10874 15952 10876 15972
rect 10876 15952 10928 15972
rect 10928 15952 10930 15972
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 10598 12824 10654 12880
rect 10598 12316 10600 12336
rect 10600 12316 10652 12336
rect 10652 12316 10654 12336
rect 10598 12280 10654 12316
rect 10782 12552 10838 12608
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11150 12552 11206 12608
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11058 11600 11114 11656
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 10782 5616 10838 5672
rect 10782 3984 10838 4040
rect 10506 2488 10562 2544
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11886 11736 11942 11792
rect 12162 11056 12218 11112
rect 11886 5788 11888 5808
rect 11888 5788 11940 5808
rect 11940 5788 11942 5808
rect 11886 5752 11942 5788
rect 12346 12688 12402 12744
rect 12530 12708 12586 12744
rect 12530 12688 12532 12708
rect 12532 12688 12584 12708
rect 12584 12688 12586 12708
rect 12898 17040 12954 17096
rect 13082 15408 13138 15464
rect 12714 14456 12770 14512
rect 12622 11736 12678 11792
rect 12714 11600 12770 11656
rect 12898 10512 12954 10568
rect 12346 9444 12402 9480
rect 12346 9424 12348 9444
rect 12348 9424 12400 9444
rect 12400 9424 12402 9444
rect 12714 8916 12716 8936
rect 12716 8916 12768 8936
rect 12768 8916 12770 8936
rect 12714 8880 12770 8916
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11334 2488 11390 2544
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11334 1944 11390 2000
rect 13082 9560 13138 9616
rect 13266 9560 13322 9616
rect 13634 12824 13690 12880
rect 13450 11056 13506 11112
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 12530 3168 12586 3224
rect 12438 2896 12494 2952
rect 12806 4664 12862 4720
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 15842 12824 15898 12880
rect 14462 6024 14518 6080
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 12898 4120 12954 4176
rect 12990 3168 13046 3224
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15566 6160 15622 6216
rect 15934 5616 15990 5672
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18418 18164 18420 18184
rect 18420 18164 18472 18184
rect 18472 18164 18474 18184
rect 18418 18128 18474 18164
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 17176 18014 17232
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17406 15952 17462 16008
rect 17130 12280 17186 12336
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 15750 3596 15806 3632
rect 15750 3576 15752 3596
rect 15752 3576 15804 3596
rect 15804 3576 15806 3596
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 17314 6296 17370 6352
rect 17130 2508 17186 2544
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 19154 5752 19210 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18878 4664 18934 4720
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17130 2488 17132 2508
rect 17132 2488 17184 2508
rect 17184 2488 17186 2508
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
<< metal3 >>
rect 0 22538 800 22568
rect 4061 22538 4127 22541
rect 0 22536 4127 22538
rect 0 22480 4066 22536
rect 4122 22480 4127 22536
rect 0 22478 4127 22480
rect 0 22448 800 22478
rect 4061 22475 4127 22478
rect 0 22130 800 22160
rect 3509 22130 3575 22133
rect 0 22128 3575 22130
rect 0 22072 3514 22128
rect 3570 22072 3575 22128
rect 0 22070 3575 22072
rect 0 22040 800 22070
rect 3509 22067 3575 22070
rect 0 21586 800 21616
rect 3601 21586 3667 21589
rect 0 21584 3667 21586
rect 0 21528 3606 21584
rect 3662 21528 3667 21584
rect 0 21526 3667 21528
rect 0 21496 800 21526
rect 3601 21523 3667 21526
rect 0 21178 800 21208
rect 3049 21178 3115 21181
rect 0 21176 3115 21178
rect 0 21120 3054 21176
rect 3110 21120 3115 21176
rect 0 21118 3115 21120
rect 0 21088 800 21118
rect 3049 21115 3115 21118
rect 0 20634 800 20664
rect 3325 20634 3391 20637
rect 0 20632 3391 20634
rect 0 20576 3330 20632
rect 3386 20576 3391 20632
rect 0 20574 3391 20576
rect 0 20544 800 20574
rect 3325 20571 3391 20574
rect 0 20226 800 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 800 20166
rect 2773 20163 2839 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19682 800 19712
rect 3417 19682 3483 19685
rect 0 19680 3483 19682
rect 0 19624 3422 19680
rect 3478 19624 3483 19680
rect 0 19622 3483 19624
rect 0 19592 800 19622
rect 3417 19619 3483 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 800 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 800 19214
rect 1945 19211 2011 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 1945 18866 2011 18869
rect 8569 18866 8635 18869
rect 1945 18864 8635 18866
rect 1945 18808 1950 18864
rect 2006 18808 8574 18864
rect 8630 18808 8635 18864
rect 1945 18806 8635 18808
rect 1945 18803 2011 18806
rect 8569 18803 8635 18806
rect 0 18730 800 18760
rect 1669 18730 1735 18733
rect 0 18728 1735 18730
rect 0 18672 1674 18728
rect 1730 18672 1735 18728
rect 0 18670 1735 18672
rect 0 18640 800 18670
rect 1669 18667 1735 18670
rect 2129 18730 2195 18733
rect 8477 18730 8543 18733
rect 2129 18728 8543 18730
rect 2129 18672 2134 18728
rect 2190 18672 8482 18728
rect 8538 18672 8543 18728
rect 2129 18670 8543 18672
rect 2129 18667 2195 18670
rect 8477 18667 8543 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 800 18352
rect 1485 18322 1551 18325
rect 12065 18322 12131 18325
rect 0 18320 1551 18322
rect 0 18264 1490 18320
rect 1546 18264 1551 18320
rect 0 18262 1551 18264
rect 0 18232 800 18262
rect 1485 18259 1551 18262
rect 7054 18320 12131 18322
rect 7054 18264 12070 18320
rect 12126 18264 12131 18320
rect 7054 18262 12131 18264
rect 2405 18186 2471 18189
rect 7054 18186 7114 18262
rect 12065 18259 12131 18262
rect 2405 18184 7114 18186
rect 2405 18128 2410 18184
rect 2466 18128 7114 18184
rect 2405 18126 7114 18128
rect 7189 18186 7255 18189
rect 18413 18186 18479 18189
rect 7189 18184 18479 18186
rect 7189 18128 7194 18184
rect 7250 18128 18418 18184
rect 18474 18128 18479 18184
rect 7189 18126 18479 18128
rect 2405 18123 2471 18126
rect 7189 18123 7255 18126
rect 18413 18123 18479 18126
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 0 17778 800 17808
rect 1669 17778 1735 17781
rect 0 17776 1735 17778
rect 0 17720 1674 17776
rect 1730 17720 1735 17776
rect 0 17718 1735 17720
rect 0 17688 800 17718
rect 1669 17715 1735 17718
rect 2497 17778 2563 17781
rect 9857 17778 9923 17781
rect 2497 17776 9923 17778
rect 2497 17720 2502 17776
rect 2558 17720 9862 17776
rect 9918 17720 9923 17776
rect 2497 17718 9923 17720
rect 2497 17715 2563 17718
rect 9857 17715 9923 17718
rect 3785 17642 3851 17645
rect 8569 17642 8635 17645
rect 3785 17640 8635 17642
rect 3785 17584 3790 17640
rect 3846 17584 8574 17640
rect 8630 17584 8635 17640
rect 3785 17582 8635 17584
rect 3785 17579 3851 17582
rect 8569 17579 8635 17582
rect 4376 17440 4696 17441
rect 0 17370 800 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 17953 17234 18019 17237
rect 22000 17234 22800 17264
rect 17953 17232 22800 17234
rect 17953 17176 17958 17232
rect 18014 17176 22800 17232
rect 17953 17174 22800 17176
rect 17953 17171 18019 17174
rect 22000 17144 22800 17174
rect 197 17098 263 17101
rect 8937 17098 9003 17101
rect 197 17096 9003 17098
rect 197 17040 202 17096
rect 258 17040 8942 17096
rect 8998 17040 9003 17096
rect 197 17038 9003 17040
rect 197 17035 263 17038
rect 8937 17035 9003 17038
rect 12750 17036 12756 17100
rect 12820 17098 12826 17100
rect 12893 17098 12959 17101
rect 12820 17096 12959 17098
rect 12820 17040 12898 17096
rect 12954 17040 12959 17096
rect 12820 17038 12959 17040
rect 12820 17036 12826 17038
rect 12893 17035 12959 17038
rect 7808 16896 8128 16897
rect 0 16826 800 16856
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 3049 16826 3115 16829
rect 0 16824 3115 16826
rect 0 16768 3054 16824
rect 3110 16768 3115 16824
rect 0 16766 3115 16768
rect 0 16736 800 16766
rect 3049 16763 3115 16766
rect 0 16418 800 16448
rect 1669 16418 1735 16421
rect 0 16416 1735 16418
rect 0 16360 1674 16416
rect 1730 16360 1735 16416
rect 0 16358 1735 16360
rect 0 16328 800 16358
rect 1669 16355 1735 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 10869 16010 10935 16013
rect 17401 16010 17467 16013
rect 10869 16008 17467 16010
rect 10869 15952 10874 16008
rect 10930 15952 17406 16008
rect 17462 15952 17467 16008
rect 10869 15950 17467 15952
rect 10869 15947 10935 15950
rect 17401 15947 17467 15950
rect 0 15874 800 15904
rect 1761 15874 1827 15877
rect 0 15872 1827 15874
rect 0 15816 1766 15872
rect 1822 15816 1827 15872
rect 0 15814 1827 15816
rect 0 15784 800 15814
rect 1761 15811 1827 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15466 800 15496
rect 1669 15466 1735 15469
rect 0 15464 1735 15466
rect 0 15408 1674 15464
rect 1730 15408 1735 15464
rect 0 15406 1735 15408
rect 0 15376 800 15406
rect 1669 15403 1735 15406
rect 10041 15466 10107 15469
rect 13077 15466 13143 15469
rect 10041 15464 13143 15466
rect 10041 15408 10046 15464
rect 10102 15408 13082 15464
rect 13138 15408 13143 15464
rect 10041 15406 13143 15408
rect 10041 15403 10107 15406
rect 13077 15403 13143 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 14922 800 14952
rect 3233 14922 3299 14925
rect 0 14920 3299 14922
rect 0 14864 3238 14920
rect 3294 14864 3299 14920
rect 0 14862 3299 14864
rect 0 14832 800 14862
rect 3233 14859 3299 14862
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 0 14514 800 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 800 14454
rect 2773 14451 2839 14454
rect 10041 14514 10107 14517
rect 12709 14514 12775 14517
rect 10041 14512 12775 14514
rect 10041 14456 10046 14512
rect 10102 14456 12714 14512
rect 12770 14456 12775 14512
rect 10041 14454 12775 14456
rect 10041 14451 10107 14454
rect 12709 14451 12775 14454
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 0 13970 800 14000
rect 2773 13970 2839 13973
rect 0 13968 2839 13970
rect 0 13912 2778 13968
rect 2834 13912 2839 13968
rect 0 13910 2839 13912
rect 0 13880 800 13910
rect 2773 13907 2839 13910
rect 7808 13632 8128 13633
rect 0 13562 800 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 4376 13088 4696 13089
rect 0 13018 800 13048
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 800 12958
rect 4061 12955 4127 12958
rect 10593 12882 10659 12885
rect 13629 12882 13695 12885
rect 15837 12882 15903 12885
rect 10593 12880 15903 12882
rect 10593 12824 10598 12880
rect 10654 12824 13634 12880
rect 13690 12824 15842 12880
rect 15898 12824 15903 12880
rect 10593 12822 15903 12824
rect 10593 12819 10659 12822
rect 13629 12819 13695 12822
rect 15837 12819 15903 12822
rect 12341 12746 12407 12749
rect 12525 12746 12591 12749
rect 12341 12744 12591 12746
rect 12341 12688 12346 12744
rect 12402 12688 12530 12744
rect 12586 12688 12591 12744
rect 12341 12686 12591 12688
rect 12341 12683 12407 12686
rect 12525 12683 12591 12686
rect 0 12610 800 12640
rect 3877 12610 3943 12613
rect 0 12608 3943 12610
rect 0 12552 3882 12608
rect 3938 12552 3943 12608
rect 0 12550 3943 12552
rect 0 12520 800 12550
rect 3877 12547 3943 12550
rect 10777 12610 10843 12613
rect 11145 12610 11211 12613
rect 10777 12608 11211 12610
rect 10777 12552 10782 12608
rect 10838 12552 11150 12608
rect 11206 12552 11211 12608
rect 10777 12550 11211 12552
rect 10777 12547 10843 12550
rect 11145 12547 11211 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 3969 12474 4035 12477
rect 4981 12474 5047 12477
rect 3969 12472 5047 12474
rect 3969 12416 3974 12472
rect 4030 12416 4986 12472
rect 5042 12416 5047 12472
rect 3969 12414 5047 12416
rect 3969 12411 4035 12414
rect 4981 12411 5047 12414
rect 10593 12338 10659 12341
rect 17125 12338 17191 12341
rect 10593 12336 17191 12338
rect 10593 12280 10598 12336
rect 10654 12280 17130 12336
rect 17186 12280 17191 12336
rect 10593 12278 17191 12280
rect 10593 12275 10659 12278
rect 17125 12275 17191 12278
rect 0 12066 800 12096
rect 4061 12066 4127 12069
rect 0 12064 4127 12066
rect 0 12008 4066 12064
rect 4122 12008 4127 12064
rect 0 12006 4127 12008
rect 0 11976 800 12006
rect 4061 12003 4127 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 11881 11794 11947 11797
rect 12617 11794 12683 11797
rect 11881 11792 12683 11794
rect 11881 11736 11886 11792
rect 11942 11736 12622 11792
rect 12678 11736 12683 11792
rect 11881 11734 12683 11736
rect 11881 11731 11947 11734
rect 12617 11731 12683 11734
rect 0 11658 800 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 800 11598
rect 3877 11595 3943 11598
rect 11053 11658 11119 11661
rect 12709 11658 12775 11661
rect 11053 11656 12775 11658
rect 11053 11600 11058 11656
rect 11114 11600 12714 11656
rect 12770 11600 12775 11656
rect 11053 11598 12775 11600
rect 11053 11595 11119 11598
rect 12709 11595 12775 11598
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 0 11114 800 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 800 11054
rect 4061 11051 4127 11054
rect 12157 11114 12223 11117
rect 13445 11114 13511 11117
rect 12157 11112 13511 11114
rect 12157 11056 12162 11112
rect 12218 11056 13450 11112
rect 13506 11056 13511 11112
rect 12157 11054 13511 11056
rect 12157 11051 12223 11054
rect 13445 11051 13511 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 0 10706 800 10736
rect 4061 10706 4127 10709
rect 0 10704 4127 10706
rect 0 10648 4066 10704
rect 4122 10648 4127 10704
rect 0 10646 4127 10648
rect 0 10616 800 10646
rect 4061 10643 4127 10646
rect 10133 10570 10199 10573
rect 12893 10570 12959 10573
rect 10133 10568 12959 10570
rect 10133 10512 10138 10568
rect 10194 10512 12898 10568
rect 12954 10512 12959 10568
rect 10133 10510 12959 10512
rect 10133 10507 10199 10510
rect 12893 10507 12959 10510
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10162 800 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 800 10102
rect 4061 10099 4127 10102
rect 4376 9824 4696 9825
rect 0 9754 800 9784
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 4061 9754 4127 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 800 9694
rect 4061 9691 4127 9694
rect 13077 9616 13143 9621
rect 13077 9560 13082 9616
rect 13138 9560 13143 9616
rect 13077 9555 13143 9560
rect 13261 9620 13327 9621
rect 13261 9616 13308 9620
rect 13372 9618 13378 9620
rect 13261 9560 13266 9616
rect 13261 9556 13308 9560
rect 13372 9558 13418 9618
rect 13372 9556 13378 9558
rect 13261 9555 13327 9556
rect 5257 9482 5323 9485
rect 9949 9482 10015 9485
rect 5257 9480 10015 9482
rect 5257 9424 5262 9480
rect 5318 9424 9954 9480
rect 10010 9424 10015 9480
rect 5257 9422 10015 9424
rect 5257 9419 5323 9422
rect 9949 9419 10015 9422
rect 12341 9482 12407 9485
rect 13080 9482 13140 9555
rect 12341 9480 13140 9482
rect 12341 9424 12346 9480
rect 12402 9424 13140 9480
rect 12341 9422 13140 9424
rect 12341 9419 12407 9422
rect 7808 9280 8128 9281
rect 0 9210 800 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 3877 9210 3943 9213
rect 0 9208 3943 9210
rect 0 9152 3882 9208
rect 3938 9152 3943 9208
rect 0 9150 3943 9152
rect 0 9120 800 9150
rect 3877 9147 3943 9150
rect 12709 8940 12775 8941
rect 12709 8936 12756 8940
rect 12820 8938 12826 8940
rect 12709 8880 12714 8936
rect 12709 8876 12756 8880
rect 12820 8878 12866 8938
rect 12820 8876 12826 8878
rect 12709 8875 12775 8876
rect 0 8802 800 8832
rect 3785 8802 3851 8805
rect 0 8800 3851 8802
rect 0 8744 3790 8800
rect 3846 8744 3851 8800
rect 0 8742 3851 8744
rect 0 8712 800 8742
rect 3785 8739 3851 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8258 800 8288
rect 3877 8258 3943 8261
rect 0 8256 3943 8258
rect 0 8200 3882 8256
rect 3938 8200 3943 8256
rect 0 8198 3943 8200
rect 0 8168 800 8198
rect 3877 8195 3943 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 0 7850 800 7880
rect 8845 7850 8911 7853
rect 0 7848 8911 7850
rect 0 7792 8850 7848
rect 8906 7792 8911 7848
rect 0 7790 8911 7792
rect 0 7760 800 7790
rect 8845 7787 8911 7790
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 0 7306 800 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 800 7246
rect 4061 7243 4127 7246
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6898 800 6928
rect 5993 6898 6059 6901
rect 0 6896 6059 6898
rect 0 6840 5998 6896
rect 6054 6840 6059 6896
rect 0 6838 6059 6840
rect 0 6808 800 6838
rect 5993 6835 6059 6838
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6354 800 6384
rect 3233 6354 3299 6357
rect 0 6352 3299 6354
rect 0 6296 3238 6352
rect 3294 6296 3299 6352
rect 0 6294 3299 6296
rect 0 6264 800 6294
rect 3233 6291 3299 6294
rect 9581 6354 9647 6357
rect 17309 6354 17375 6357
rect 9581 6352 17375 6354
rect 9581 6296 9586 6352
rect 9642 6296 17314 6352
rect 17370 6296 17375 6352
rect 9581 6294 17375 6296
rect 9581 6291 9647 6294
rect 17309 6291 17375 6294
rect 8569 6218 8635 6221
rect 15561 6218 15627 6221
rect 8569 6216 15627 6218
rect 8569 6160 8574 6216
rect 8630 6160 15566 6216
rect 15622 6160 15627 6216
rect 8569 6158 15627 6160
rect 8569 6155 8635 6158
rect 15561 6155 15627 6158
rect 10041 6082 10107 6085
rect 14457 6082 14523 6085
rect 10041 6080 14523 6082
rect 10041 6024 10046 6080
rect 10102 6024 14462 6080
rect 14518 6024 14523 6080
rect 10041 6022 14523 6024
rect 10041 6019 10107 6022
rect 14457 6019 14523 6022
rect 7808 6016 8128 6017
rect 0 5946 800 5976
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5886 4906 5946
rect 0 5856 800 5886
rect 4846 5810 4906 5886
rect 8109 5810 8175 5813
rect 4846 5808 8175 5810
rect 4846 5752 8114 5808
rect 8170 5752 8175 5808
rect 4846 5750 8175 5752
rect 8109 5747 8175 5750
rect 9765 5810 9831 5813
rect 11881 5810 11947 5813
rect 9765 5808 11947 5810
rect 9765 5752 9770 5808
rect 9826 5752 11886 5808
rect 11942 5752 11947 5808
rect 9765 5750 11947 5752
rect 9765 5747 9831 5750
rect 11881 5747 11947 5750
rect 19149 5810 19215 5813
rect 22000 5810 22800 5840
rect 19149 5808 22800 5810
rect 19149 5752 19154 5808
rect 19210 5752 22800 5808
rect 19149 5750 22800 5752
rect 19149 5747 19215 5750
rect 22000 5720 22800 5750
rect 10777 5674 10843 5677
rect 15929 5674 15995 5677
rect 10777 5672 15995 5674
rect 10777 5616 10782 5672
rect 10838 5616 15934 5672
rect 15990 5616 15995 5672
rect 10777 5614 15995 5616
rect 10777 5611 10843 5614
rect 15929 5611 15995 5614
rect 4376 5472 4696 5473
rect 0 5402 800 5432
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 3785 5402 3851 5405
rect 0 5400 3851 5402
rect 0 5344 3790 5400
rect 3846 5344 3851 5400
rect 0 5342 3851 5344
rect 0 5312 800 5342
rect 3785 5339 3851 5342
rect 0 4994 800 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 800 4934
rect 4061 4931 4127 4934
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 12801 4722 12867 4725
rect 18873 4722 18939 4725
rect 12801 4720 18939 4722
rect 12801 4664 12806 4720
rect 12862 4664 18878 4720
rect 18934 4664 18939 4720
rect 12801 4662 18939 4664
rect 12801 4659 12867 4662
rect 18873 4659 18939 4662
rect 0 4450 800 4480
rect 3877 4450 3943 4453
rect 0 4448 3943 4450
rect 0 4392 3882 4448
rect 3938 4392 3943 4448
rect 0 4390 3943 4392
rect 0 4360 800 4390
rect 3877 4387 3943 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 7281 4178 7347 4181
rect 12893 4178 12959 4181
rect 7281 4176 12959 4178
rect 7281 4120 7286 4176
rect 7342 4120 12898 4176
rect 12954 4120 12959 4176
rect 7281 4118 12959 4120
rect 7281 4115 7347 4118
rect 12893 4115 12959 4118
rect 0 4042 800 4072
rect 7649 4042 7715 4045
rect 0 4040 7715 4042
rect 0 3984 7654 4040
rect 7710 3984 7715 4040
rect 0 3982 7715 3984
rect 0 3952 800 3982
rect 7649 3979 7715 3982
rect 8937 4042 9003 4045
rect 10777 4042 10843 4045
rect 8937 4040 10843 4042
rect 8937 3984 8942 4040
rect 8998 3984 10782 4040
rect 10838 3984 10843 4040
rect 8937 3982 10843 3984
rect 8937 3979 9003 3982
rect 10777 3979 10843 3982
rect 3417 3906 3483 3909
rect 3190 3904 3483 3906
rect 3190 3848 3422 3904
rect 3478 3848 3483 3904
rect 3190 3846 3483 3848
rect 0 3498 800 3528
rect 3190 3501 3250 3846
rect 3417 3843 3483 3846
rect 4521 3906 4587 3909
rect 5533 3906 5599 3909
rect 4521 3904 5599 3906
rect 4521 3848 4526 3904
rect 4582 3848 5538 3904
rect 5594 3848 5599 3904
rect 4521 3846 5599 3848
rect 4521 3843 4587 3846
rect 5533 3843 5599 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 3969 3634 4035 3637
rect 6545 3634 6611 3637
rect 15745 3634 15811 3637
rect 3969 3632 15811 3634
rect 3969 3576 3974 3632
rect 4030 3576 6550 3632
rect 6606 3576 15750 3632
rect 15806 3576 15811 3632
rect 3969 3574 15811 3576
rect 3969 3571 4035 3574
rect 6545 3571 6611 3574
rect 15745 3571 15811 3574
rect 3141 3498 3250 3501
rect 0 3496 3250 3498
rect 0 3440 3146 3496
rect 3202 3440 3250 3496
rect 0 3438 3250 3440
rect 0 3408 800 3438
rect 3141 3435 3207 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 12525 3226 12591 3229
rect 12985 3226 13051 3229
rect 12525 3224 13051 3226
rect 12525 3168 12530 3224
rect 12586 3168 12990 3224
rect 13046 3168 13051 3224
rect 12525 3166 13051 3168
rect 12525 3163 12591 3166
rect 12985 3163 13051 3166
rect 0 3090 800 3120
rect 3509 3090 3575 3093
rect 0 3088 3575 3090
rect 0 3032 3514 3088
rect 3570 3032 3575 3088
rect 0 3030 3575 3032
rect 0 3000 800 3030
rect 3509 3027 3575 3030
rect 9305 2954 9371 2957
rect 12433 2954 12499 2957
rect 9305 2952 12499 2954
rect 9305 2896 9310 2952
rect 9366 2896 12438 2952
rect 12494 2896 12499 2952
rect 9305 2894 12499 2896
rect 9305 2891 9371 2894
rect 12433 2891 12499 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 800 2576
rect 1761 2546 1827 2549
rect 0 2544 1827 2546
rect 0 2488 1766 2544
rect 1822 2488 1827 2544
rect 0 2486 1827 2488
rect 0 2456 800 2486
rect 1761 2483 1827 2486
rect 10501 2546 10567 2549
rect 11329 2546 11395 2549
rect 17125 2546 17191 2549
rect 10501 2544 17191 2546
rect 10501 2488 10506 2544
rect 10562 2488 11334 2544
rect 11390 2488 17130 2544
rect 17186 2488 17191 2544
rect 10501 2486 17191 2488
rect 10501 2483 10567 2486
rect 11329 2483 11395 2486
rect 17125 2483 17191 2486
rect 4376 2208 4696 2209
rect 0 2138 800 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 800 2078
rect 2865 2075 2931 2078
rect 11329 2002 11395 2005
rect 13302 2002 13308 2004
rect 11329 2000 13308 2002
rect 11329 1944 11334 2000
rect 11390 1944 13308 2000
rect 11329 1942 13308 1944
rect 11329 1939 11395 1942
rect 13302 1940 13308 1942
rect 13372 1940 13378 2004
rect 0 1594 800 1624
rect 3233 1594 3299 1597
rect 0 1592 3299 1594
rect 0 1536 3238 1592
rect 3294 1536 3299 1592
rect 0 1534 3299 1536
rect 0 1504 800 1534
rect 3233 1531 3299 1534
rect 0 1186 800 1216
rect 3601 1186 3667 1189
rect 0 1184 3667 1186
rect 0 1128 3606 1184
rect 3662 1128 3667 1184
rect 0 1126 3667 1128
rect 0 1096 800 1126
rect 3601 1123 3667 1126
rect 6453 914 6519 917
rect 7097 914 7163 917
rect 6453 912 7163 914
rect 6453 856 6458 912
rect 6514 856 7102 912
rect 7158 856 7163 912
rect 6453 854 7163 856
rect 6453 851 6519 854
rect 7097 851 7163 854
rect 0 642 800 672
rect 3785 642 3851 645
rect 0 640 3851 642
rect 0 584 3790 640
rect 3846 584 3851 640
rect 0 582 3851 584
rect 0 552 800 582
rect 3785 579 3851 582
rect 0 234 800 264
rect 4061 234 4127 237
rect 0 232 4127 234
rect 0 176 4066 232
rect 4122 176 4127 232
rect 0 174 4127 176
rect 0 144 800 174
rect 4061 171 4127 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 12756 17036 12820 17100
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 13308 9616 13372 9620
rect 13308 9560 13322 9616
rect 13322 9560 13372 9616
rect 13308 9556 13372 9560
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 12756 8936 12820 8940
rect 12756 8880 12770 8936
rect 12770 8880 12820 8936
rect 12756 8876 12820 8880
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 13308 1940 13372 2004
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 12755 17100 12821 17101
rect 12755 17036 12756 17100
rect 12820 17036 12821 17100
rect 12755 17035 12821 17036
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 12758 8941 12818 17035
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 13307 9620 13373 9621
rect 13307 9556 13308 9620
rect 13372 9556 13373 9620
rect 13307 9555 13373 9556
rect 12755 8940 12821 8941
rect 12755 8876 12756 8940
rect 12820 8876 12821 8940
rect 12755 8875 12821 8876
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 13310 2005 13370 9555
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 13307 2004 13373 2005
rect 13307 1940 13308 2004
rect 13372 1940 13373 2004
rect 13307 1939 13373 1940
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608763155
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608763155
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_214
timestamp 1608763155
transform 1 0 20792 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608763155
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608763155
transform 1 0 18492 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608763155
transform 1 0 19320 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_193
timestamp 1608763155
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1608763155
transform 1 0 19228 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1608763155
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608763155
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1608763155
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1608763155
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1608763155
transform 1 0 18308 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608763155
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_147
timestamp 1608763155
transform 1 0 14628 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1608763155
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608763155
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1608763155
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_135
timestamp 1608763155
transform 1 0 13524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608763155
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608763155
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_115
timestamp 1608763155
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_123
timestamp 1608763155
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608763155
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608763155
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_89
timestamp 1608763155
transform 1 0 9292 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1608763155
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608763155
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1608763155
transform 1 0 6900 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_67
timestamp 1608763155
transform 1 0 7268 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_77
timestamp 1608763155
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608763155
transform 1 0 5520 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608763155
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_47
timestamp 1608763155
transform 1 0 5428 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1608763155
transform 1 0 6348 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1608763155
transform 1 0 6716 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608763155
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608763155
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608763155
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1608763155
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1608763155
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_35
timestamp 1608763155
transform 1 0 4324 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608763155
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608763155
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608763155
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608763155
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1608763155
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1608763155
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1608763155
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608763155
transform 1 0 20332 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608763155
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_213
timestamp 1608763155
transform 1 0 20700 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1608763155
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608763155
transform 1 0 19044 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_188
timestamp 1608763155
transform 1 0 18400 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_194
timestamp 1608763155
transform 1 0 18952 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1608763155
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608763155
transform 1 0 16744 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608763155
transform 1 0 17296 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608763155
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608763155
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_168
timestamp 1608763155
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 1608763155
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1608763155
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608763155
transform 1 0 14536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608763155
transform 1 0 15088 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608763155
transform 1 0 15640 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608763155
transform 1 0 16192 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 1608763155
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1608763155
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1608763155
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608763155
transform 1 0 13432 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608763155
transform 1 0 13984 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 12696 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1608763155
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1608763155
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1608763155
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 11500 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608763155
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1608763155
transform 1 0 11040 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_112
timestamp 1608763155
transform 1 0 11408 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1608763155
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1608763155
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 9568 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 8832 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1608763155
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608763155
transform 1 0 7820 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1608763155
transform 1 0 7360 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_72
timestamp 1608763155
transform 1 0 7728 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1608763155
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608763155
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1608763155
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608763155
transform 1 0 3128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 4876 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608763155
transform 1 0 3680 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1608763155
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_37
timestamp 1608763155
transform 1 0 4508 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2392 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1656 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608763155
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1608763155
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1608763155
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_20
timestamp 1608763155
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608763155
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608763155
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608763155
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608763155
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608763155
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608763155
transform 1 0 18952 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_188
timestamp 1608763155
transform 1 0 18400 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1608763155
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608763155
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_178
timestamp 1608763155
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608763155
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608763155
transform 1 0 16008 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608763155
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1608763155
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1608763155
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1608763155
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608763155
transform 1 0 13248 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_130
timestamp 1608763155
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1608763155
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1608763155
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 11592 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1608763155
transform 1 0 11132 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_113
timestamp 1608763155
transform 1 0 11500 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608763155
transform 1 0 9108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608763155
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_84
timestamp 1608763155
transform 1 0 8832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608763155
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608763155
transform 1 0 6900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 7360 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1608763155
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608763155
transform 1 0 6440 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_56
timestamp 1608763155
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 1608763155
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608763155
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 4784 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608763155
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1608763155
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_36
timestamp 1608763155
transform 1 0 4416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608763155
transform 1 0 1472 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2024 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608763155
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608763155
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1608763155
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_8
timestamp 1608763155
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1608763155
transform 1 0 2576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608763155
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1608763155
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 18400 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_194
timestamp 1608763155
transform 1 0 18952 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_206
timestamp 1608763155
transform 1 0 20056 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 16560 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608763155
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_174
timestamp 1608763155
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1608763155
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1608763155
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 14996 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_150
timestamp 1608763155
transform 1 0 14904 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1608763155
transform 1 0 15548 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1608763155
transform 1 0 16284 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608763155
transform 1 0 13984 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608763155
transform 1 0 12696 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 13248 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_130
timestamp 1608763155
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1608763155
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_144
timestamp 1608763155
transform 1 0 14352 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608763155
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608763155
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1608763155
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1608763155
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608763155
transform 1 0 9660 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_84
timestamp 1608763155
transform 1 0 8832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1608763155
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_102
timestamp 1608763155
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 7360 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608763155
transform 1 0 5704 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608763155
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_42
timestamp 1608763155
transform 1 0 4968 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608763155
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_62
timestamp 1608763155
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 3496 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1608763155
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608763155
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 1840 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608763155
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_6
timestamp 1608763155
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608763155
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608763155
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608763155
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608763155
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608763155
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1608763155
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608763155
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608763155
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1608763155
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608763155
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608763155
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608763155
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1608763155
transform 1 0 13800 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_136
timestamp 1608763155
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 11132 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_108
timestamp 1608763155
transform 1 0 11040 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1608763155
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 9752 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608763155
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_86
timestamp 1608763155
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1608763155
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_100
timestamp 1608763155
transform 1 0 10304 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608763155
transform 1 0 8188 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_75
timestamp 1608763155
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 6532 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608763155
transform 1 0 4968 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1608763155
transform 1 0 5796 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608763155
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608763155
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1608763155
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_36
timestamp 1608763155
transform 1 0 4416 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608763155
transform 1 0 1472 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608763155
transform 1 0 2852 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608763155
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1608763155
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_8
timestamp 1608763155
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_16
timestamp 1608763155
transform 1 0 2576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608763155
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608763155
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608763155
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608763155
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608763155
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1608763155
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1608763155
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1608763155
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1608763155
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608763155
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1608763155
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1608763155
transform 1 0 16652 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608763155
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608763155
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608763155
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_146
timestamp 1608763155
transform 1 0 14536 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608763155
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608763155
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608763155
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_157
timestamp 1608763155
transform 1 0 15548 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 13064 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 14076 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1608763155
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1608763155
transform 1 0 13248 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_140
timestamp 1608763155
transform 1 0 13984 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608763155
transform 1 0 11592 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1608763155
transform 1 0 11316 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608763155
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608763155
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1608763155
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_120
timestamp 1608763155
transform 1 0 12144 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1608763155
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1608763155
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1608763155
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 9936 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608763155
transform 1 0 8924 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608763155
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608763155
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1608763155
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1608763155
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608763155
transform 1 0 7544 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1608763155
transform 1 0 8556 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1608763155
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1608763155
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_79
timestamp 1608763155
transform 1 0 8372 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608763155
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 5888 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608763155
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_48
timestamp 1608763155
transform 1 0 5520 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1608763155
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1608763155
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1608763155
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 4508 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608763155
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1608763155
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1608763155
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 2852 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608763155
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1608763155
transform 1 0 2576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1608763155
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608763155
transform 1 0 1472 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608763155
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608763155
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608763155
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1608763155
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1608763155
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1608763155
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1608763155
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608763155
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1608763155
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1608763155
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608763155
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_172
timestamp 1608763155
transform 1 0 16928 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1608763155
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608763155
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608763155
transform 1 0 15088 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1608763155
transform 1 0 16100 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 1608763155
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1608763155
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608763155
transform 1 0 14076 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1608763155
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608763155
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_111
timestamp 1608763155
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1608763155
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 8832 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608763155
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1608763155
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 7176 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_82
timestamp 1608763155
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608763155
transform 1 0 5244 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608763155
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_44
timestamp 1608763155
transform 1 0 5152 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_54
timestamp 1608763155
transform 1 0 6072 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1608763155
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1608763155
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608763155
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608763155
transform 1 0 3956 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_24
timestamp 1608763155
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1608763155
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1608763155
transform 1 0 4784 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608763155
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2760 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608763155
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1608763155
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1608763155
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1608763155
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608763155
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608763155
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1608763155
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608763155
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608763155
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_199
timestamp 1608763155
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_175
timestamp 1608763155
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_187
timestamp 1608763155
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1608763155
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608763155
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608763155
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_163
timestamp 1608763155
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 13524 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_130
timestamp 1608763155
transform 1 0 13064 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_134
timestamp 1608763155
transform 1 0 13432 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608763155
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608763155
transform 1 0 12236 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1608763155
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608763155
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608763155
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608763155
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1608763155
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608763155
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1608763155
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1608763155
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 5152 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 6808 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1608763155
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608763155
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_23
timestamp 1608763155
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608763155
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608763155
transform 1 0 1564 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608763155
transform 1 0 2852 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2116 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608763155
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1608763155
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1608763155
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1608763155
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608763155
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1608763155
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1608763155
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608763155
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1608763155
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1608763155
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608763155
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1608763155
transform 1 0 15180 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1608763155
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_162
timestamp 1608763155
transform 1 0 16008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608763155
transform 1 0 13708 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1608763155
transform 1 0 14168 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1608763155
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_136
timestamp 1608763155
transform 1 0 13616 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_140
timestamp 1608763155
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608763155
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608763155
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1608763155
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608763155
transform 1 0 9660 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608763155
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1608763155
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1608763155
transform 1 0 9936 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1608763155
transform 1 0 10304 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 8096 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1608763155
transform 1 0 7636 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1608763155
transform 1 0 8004 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_79
timestamp 1608763155
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608763155
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608763155
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608763155
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_49
timestamp 1608763155
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_54
timestamp 1608763155
transform 1 0 6072 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608763155
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 4140 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_25
timestamp 1608763155
transform 1 0 3404 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608763155
transform 1 0 1564 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2116 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2852 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608763155
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1608763155
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1608763155
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_17
timestamp 1608763155
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608763155
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608763155
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1608763155
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608763155
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608763155
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1608763155
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1608763155
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1608763155
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608763155
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608763155
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1608763155
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1608763155
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1608763155
transform 1 0 13984 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1608763155
transform 1 0 13156 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1608763155
transform 1 0 13892 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608763155
transform 1 0 11316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1608763155
transform 1 0 12328 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_110
timestamp 1608763155
transform 1 0 11224 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1608763155
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608763155
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608763155
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608763155
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_102
timestamp 1608763155
transform 1 0 10488 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 7912 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_65
timestamp 1608763155
transform 1 0 7084 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1608763155
transform 1 0 7820 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1608763155
transform 1 0 6256 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_48
timestamp 1608763155
transform 1 0 5520 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp 1608763155
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608763155
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1608763155
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608763155
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 2208 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1608763155
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608763155
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1608763155
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1608763155
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1608763155
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608763155
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1608763155
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1608763155
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608763155
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_167
timestamp 1608763155
transform 1 0 16468 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1608763155
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608763155
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 14996 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608763155
transform 1 0 13156 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_128
timestamp 1608763155
transform 1 0 12880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1608763155
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_145
timestamp 1608763155
transform 1 0 14444 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608763155
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608763155
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 12604 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1608763155
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608763155
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1608763155
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608763155
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1608763155
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 6992 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_80
timestamp 1608763155
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608763155
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608763155
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_45
timestamp 1608763155
transform 1 0 5244 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1608763155
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1608763155
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608763155
transform 1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1608763155
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_26
timestamp 1608763155
transform 1 0 3496 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1608763155
transform 1 0 4876 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608763155
transform 1 0 2576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1840 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608763155
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1608763155
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1608763155
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1608763155
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1608763155
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608763155
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608763155
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608763155
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1608763155
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608763155
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608763155
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1608763155
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1608763155
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_199
timestamp 1608763155
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608763155
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1608763155
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1608763155
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_175
timestamp 1608763155
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1608763155
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1608763155
transform 1 0 15456 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608763155
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608763155
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_154
timestamp 1608763155
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_165
timestamp 1608763155
transform 1 0 16284 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1608763155
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_163
timestamp 1608763155
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 12788 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 13432 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1608763155
transform 1 0 14444 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1608763155
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_131
timestamp 1608763155
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608763155
transform 1 0 11316 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608763155
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608763155
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_111
timestamp 1608763155
transform 1 0 11316 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1608763155
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1608763155
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1608763155
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 9844 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608763155
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_89
timestamp 1608763155
transform 1 0 9292 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1608763155
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1608763155
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608763155
transform 1 0 8648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608763155
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1608763155
transform 1 0 7636 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1608763155
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_77
timestamp 1608763155
transform 1 0 8188 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1608763155
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_80
timestamp 1608763155
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 5980 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608763155
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608763155
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608763155
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608763155
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1608763155
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1608763155
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608763155
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608763155
transform 1 0 3956 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608763155
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_29
timestamp 1608763155
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1608763155
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608763155
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608763155
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1608763155
transform 1 0 4692 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608763155
transform 1 0 2944 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608763155
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1608763155
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_14
timestamp 1608763155
transform 1 0 2392 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608763155
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608763155
transform 1 0 1932 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1840 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608763155
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608763155
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1608763155
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1608763155
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1608763155
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608763155
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608763155
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608763155
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608763155
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_194
timestamp 1608763155
transform 1 0 18952 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1608763155
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_170
timestamp 1608763155
transform 1 0 16744 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_182
timestamp 1608763155
transform 1 0 17848 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608763155
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1608763155
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608763155
transform 1 0 13340 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1608763155
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_142
timestamp 1608763155
transform 1 0 14168 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608763155
transform 1 0 12328 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1608763155
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 10672 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608763155
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608763155
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1608763155
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1608763155
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608763155
transform 1 0 7452 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608763155
transform 1 0 8464 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1608763155
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1608763155
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 5704 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1608763155
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608763155
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_28
timestamp 1608763155
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 1472 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608763155
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608763155
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1608763155
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608763155
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1608763155
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1608763155
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608763155
transform 1 0 16744 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608763155
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_168
timestamp 1608763155
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1608763155
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1608763155
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 15088 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1608763155
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1608763155
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1608763155
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608763155
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608763155
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1608763155
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608763155
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608763155
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608763155
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1608763155
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1608763155
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608763155
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 7820 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_65
timestamp 1608763155
transform 1 0 7084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1608763155
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608763155
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608763155
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608763155
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608763155
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608763155
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1608763155
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1608763155
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1608763155
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1608763155
transform 1 0 2576 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1656 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608763155
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1608763155
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1608763155
transform 1 0 2208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608763155
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608763155
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1608763155
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608763155
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608763155
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_198
timestamp 1608763155
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_174
timestamp 1608763155
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_186
timestamp 1608763155
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608763155
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1608763155
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608763155
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1608763155
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608763155
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1608763155
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1608763155
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608763155
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608763155
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608763155
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 10120 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1608763155
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 7084 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608763155
transform 1 0 8740 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1608763155
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1608763155
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1608763155
transform 1 0 6072 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_48
timestamp 1608763155
transform 1 0 5520 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608763155
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1608763155
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608763155
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608763155
transform 1 0 1472 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 2024 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608763155
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1608763155
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_8
timestamp 1608763155
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608763155
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1608763155
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1608763155
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608763155
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1608763155
transform 1 0 16652 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608763155
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1608763155
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1608763155
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1608763155
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1608763155
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1608763155
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1608763155
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1608763155
transform 1 0 14260 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608763155
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608763155
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_107
timestamp 1608763155
transform 1 0 10948 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1608763155
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608763155
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1608763155
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1608763155
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608763155
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608763155
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1608763155
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608763155
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608763155
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1608763155
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1608763155
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_31
timestamp 1608763155
transform 1 0 3956 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1608763155
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608763155
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608763155
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1608763155
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1608763155
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608763155
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608763155
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608763155
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608763155
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608763155
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1608763155
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1608763155
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_194
timestamp 1608763155
transform 1 0 18952 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1608763155
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608763155
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1608763155
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608763155
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1608763155
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_170
timestamp 1608763155
transform 1 0 16744 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_182
timestamp 1608763155
transform 1 0 17848 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608763155
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1608763155
transform 1 0 15088 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608763155
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1608763155
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_161
timestamp 1608763155
transform 1 0 15916 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_146
timestamp 1608763155
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608763155
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608763155
transform 1 0 14260 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608763155
transform 1 0 14076 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1608763155
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1608763155
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 12604 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608763155
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608763155
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1608763155
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608763155
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1608763155
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1608763155
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1608763155
transform 1 0 10856 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 10488 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608763155
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_98
timestamp 1608763155
transform 1 0 10120 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1608763155
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608763155
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1608763155
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1608763155
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 8648 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608763155
transform 1 0 7452 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608763155
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608763155
transform 1 0 8096 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 6992 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_67
timestamp 1608763155
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1608763155
transform 1 0 8280 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1608763155
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1608763155
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608763155
transform 1 0 5612 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1608763155
transform 1 0 6072 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608763155
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1608763155
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1608763155
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608763155
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_52
timestamp 1608763155
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608763155
transform 1 0 3680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 4416 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1608763155
transform 1 0 4600 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608763155
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_26
timestamp 1608763155
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_31
timestamp 1608763155
transform 1 0 3956 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_37
timestamp 1608763155
transform 1 0 4508 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1608763155
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1608763155
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 2024 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1608763155
transform 1 0 2576 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608763155
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608763155
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608763155
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1608763155
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1608763155
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1608763155
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_14
timestamp 1608763155
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608763155
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608763155
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608763155
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608763155
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1608763155
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1608763155
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1608763155
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608763155
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1608763155
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608763155
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1608763155
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1608763155
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1608763155
transform 1 0 13892 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1608763155
transform 1 0 13340 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608763155
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608763155
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1608763155
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_119
timestamp 1608763155
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_123
timestamp 1608763155
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608763155
transform 1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1608763155
transform 1 0 10212 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608763155
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1608763155
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608763155
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1608763155
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1608763155
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 7452 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_67
timestamp 1608763155
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608763155
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 5520 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1608763155
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608763155
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608763155
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1608763155
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608763155
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1608763155
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608763155
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608763155
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1608763155
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608763155
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1608763155
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608763155
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1608763155
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 14260 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1608763155
transform 1 0 13248 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_128
timestamp 1608763155
transform 1 0 12880 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1608763155
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608763155
transform 1 0 10948 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608763155
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1608763155
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1608763155
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1608763155
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 9292 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_87
timestamp 1608763155
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608763155
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608763155
transform 1 0 7268 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1608763155
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1608763155
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608763155
transform 1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608763155
transform 1 0 5428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608763155
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1608763155
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_56
timestamp 1608763155
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1608763155
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608763155
transform 1 0 3864 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1608763155
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_39
timestamp 1608763155
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608763155
transform 1 0 2852 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1932 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608763155
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1608763155
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1608763155
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608763155
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608763155
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1608763155
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608763155
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608763155
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1608763155
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_175
timestamp 1608763155
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1608763155
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608763155
transform 1 0 14536 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608763155
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608763155
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1608763155
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_163
timestamp 1608763155
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 12788 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_143
timestamp 1608763155
transform 1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 10764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_108
timestamp 1608763155
transform 1 0 11040 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1608763155
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1608763155
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608763155
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608763155
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_102
timestamp 1608763155
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1608763155
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608763155
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1608763155
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1608763155
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608763155
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1608763155
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 4692 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608763155
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1608763155
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1608763155
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1608763155
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 2208 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 1472 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608763155
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608763155
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1608763155
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608763155
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1608763155
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1608763155
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608763155
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1608763155
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1608763155
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1608763155
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 15456 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1608763155
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608763155
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608763155
transform 1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp 1608763155
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1608763155
transform 1 0 14076 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608763155
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608763155
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608763155
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 10672 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1608763155
transform 1 0 9660 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1608763155
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1608763155
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1608763155
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1608763155
transform 1 0 8280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608763155
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608763155
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1608763155
transform 1 0 5244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1608763155
transform 1 0 5612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608763155
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608763155
transform 1 0 3404 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608763155
transform 1 0 4416 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1608763155
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1608763155
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608763155
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608763155
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608763155
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1608763155
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608763155
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608763155
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1608763155
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608763155
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608763155
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608763155
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 18860 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1608763155
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_187
timestamp 1608763155
transform 1 0 18308 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608763155
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608763155
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608763155
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1608763155
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608763155
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1608763155
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1608763155
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_139
timestamp 1608763155
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 11408 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1608763155
transform 1 0 10948 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1608763155
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608763155
transform 1 0 10672 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1608763155
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608763155
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1608763155
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1608763155
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1608763155
transform 1 0 8464 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1608763155
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 6808 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1608763155
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_49
timestamp 1608763155
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 1608763155
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 4140 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608763155
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_26
timestamp 1608763155
transform 1 0 3496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1608763155
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_32
timestamp 1608763155
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 2024 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608763155
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1608763155
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1608763155
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608763155
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608763155
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608763155
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1608763155
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1608763155
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608763155
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608763155
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_212
timestamp 1608763155
transform 1 0 20608 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 18860 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 18952 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1608763155
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1608763155
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_200
timestamp 1608763155
transform 1 0 19504 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 17204 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608763155
transform 1 0 16560 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608763155
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_173
timestamp 1608763155
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_177
timestamp 1608763155
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_184
timestamp 1608763155
transform 1 0 18032 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608763155
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 15548 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1608763155
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608763155
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1608763155
transform 1 0 14628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608763155
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1608763155
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1608763155
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1608763155
transform 1 0 16008 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 12788 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1608763155
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1608763155
transform 1 0 12696 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1608763155
transform 1 0 14260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_132
timestamp 1608763155
transform 1 0 13248 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1608763155
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608763155
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1608763155
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608763155
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608763155
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1608763155
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_120
timestamp 1608763155
transform 1 0 12144 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_114
timestamp 1608763155
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 9108 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608763155
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608763155
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1608763155
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608763155
transform 1 0 8464 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608763155
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608763155
transform 1 0 7452 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1608763155
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_79
timestamp 1608763155
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1608763155
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1608763155
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1608763155
transform 1 0 8740 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1608763155
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608763155
transform 1 0 6072 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608763155
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608763155
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_52
timestamp 1608763155
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1608763155
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608763155
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1608763155
transform 1 0 5060 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1608763155
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608763155
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608763155
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608763155
transform 1 0 3864 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608763155
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608763155
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1608763155
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1608763155
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_28
timestamp 1608763155
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_39
timestamp 1608763155
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 1380 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608763155
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608763155
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608763155
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608763155
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_19
timestamp 1608763155
transform 1 0 2852 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 1608763155
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608763155
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1608763155
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608763155
transform 1 0 19780 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1608763155
transform 1 0 19136 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1608763155
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1608763155
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608763155
transform 1 0 17388 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608763155
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1608763155
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1608763155
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1608763155
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608763155
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_160
timestamp 1608763155
transform 1 0 15824 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 14352 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_5_132
timestamp 1608763155
transform 1 0 13248 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608763155
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608763155
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608763155
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1608763155
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608763155
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608763155
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1608763155
transform 1 0 9292 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1608763155
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 7084 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1608763155
transform 1 0 8556 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 5060 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608763155
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_42
timestamp 1608763155
transform 1 0 4968 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608763155
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_62
timestamp 1608763155
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_34
timestamp 1608763155
transform 1 0 4232 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 2760 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608763155
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608763155
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608763155
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1608763155
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608763155
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608763155
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608763155
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608763155
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608763155
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_193
timestamp 1608763155
transform 1 0 18860 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_205
timestamp 1608763155
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608763155
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 18308 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1608763155
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_185
timestamp 1608763155
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608763155
transform 1 0 16284 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1608763155
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608763155
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608763155
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1608763155
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 13524 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1608763155
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608763155
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608763155
transform 1 0 10764 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1608763155
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_125
timestamp 1608763155
transform 1 0 12604 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1608763155
transform 1 0 9752 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608763155
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608763155
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1608763155
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1608763155
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1608763155
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1608763155
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1608763155
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1608763155
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608763155
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_48
timestamp 1608763155
transform 1 0 5520 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp 1608763155
transform 1 0 6256 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608763155
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_24
timestamp 1608763155
transform 1 0 3312 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608763155
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 1840 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608763155
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1608763155
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1608763155
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608763155
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_212
timestamp 1608763155
transform 1 0 20608 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_188
timestamp 1608763155
transform 1 0 18400 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_200
timestamp 1608763155
transform 1 0 19504 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608763155
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608763155
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_174
timestamp 1608763155
transform 1 0 17112 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608763155
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608763155
transform 1 0 15272 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1608763155
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_152
timestamp 1608763155
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1608763155
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608763155
transform 1 0 13432 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608763155
transform 1 0 14260 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1608763155
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1608763155
transform 1 0 13800 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1608763155
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 11592 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608763155
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608763155
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1608763155
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608763155
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1608763155
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1608763155
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1608763155
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1608763155
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1608763155
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_71
timestamp 1608763155
transform 1 0 7636 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1608763155
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608763155
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608763155
transform 1 0 5704 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608763155
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_48
timestamp 1608763155
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608763155
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608763155
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608763155
transform 1 0 3680 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1608763155
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1608763155
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1608763155
transform 1 0 2484 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608763155
transform 1 0 1472 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608763155
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608763155
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1608763155
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608763155
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608763155
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1608763155
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608763155
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608763155
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_193
timestamp 1608763155
transform 1 0 18860 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1608763155
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608763155
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608763155
transform 1 0 17388 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1608763155
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_175
timestamp 1608763155
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_181
timestamp 1608763155
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608763155
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608763155
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608763155
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1608763155
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608763155
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1608763155
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1608763155
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1608763155
transform 1 0 12604 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_123
timestamp 1608763155
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608763155
transform 1 0 9752 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608763155
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608763155
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1608763155
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1608763155
transform 1 0 10580 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608763155
transform 1 0 7544 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1608763155
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1608763155
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1608763155
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1608763155
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608763155
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608763155
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_22
timestamp 1608763155
transform 1 0 3128 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608763155
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1608763155
transform 1 0 4048 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1608763155
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 1656 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608763155
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1608763155
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608763155
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608763155
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608763155
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1608763155
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1608763155
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608763155
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_209
timestamp 1608763155
transform 1 0 20332 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp 1608763155
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_197
timestamp 1608763155
transform 1 0 19228 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608763155
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608763155
transform 1 0 20240 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_203
timestamp 1608763155
transform 1 0 19780 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_207
timestamp 1608763155
transform 1 0 20148 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608763155
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608763155
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1608763155
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1608763155
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1608763155
transform 1 0 18400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_192
timestamp 1608763155
transform 1 0 18768 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608763155
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608763155
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608763155
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608763155
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608763155
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1608763155
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608763155
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1608763155
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1608763155
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608763155
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608763155
transform 1 0 17112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1608763155
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1608763155
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608763155
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608763155
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608763155
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608763155
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 15824 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608763155
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608763155
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1608763155
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1608763155
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1608763155
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1608763155
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608763155
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 14168 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 14260 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1608763155
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_137
timestamp 1608763155
transform 1 0 13708 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1608763155
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608763155
transform 1 0 12512 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608763155
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608763155
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608763155
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1608763155
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608763155
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1608763155
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608763155
transform 1 0 10856 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608763155
transform 1 0 11408 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1608763155
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608763155
transform 1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608763155
transform 1 0 9200 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608763155
transform 1 0 10396 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608763155
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608763155
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1608763155
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp 1608763155
transform 1 0 10120 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1608763155
transform 1 0 9108 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1608763155
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 7084 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1608763155
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608763155
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1608763155
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83
timestamp 1608763155
transform 1 0 8740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp 1608763155
transform 1 0 8556 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1608763155
transform 1 0 4968 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608763155
transform 1 0 5980 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608763155
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608763155
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1608763155
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1608763155
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1608763155
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1608763155
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608763155
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608763155
transform 1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608763155
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1608763155
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1608763155
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1608763155
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1608763155
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_31
timestamp 1608763155
transform 1 0 3956 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608763155
transform 1 0 2024 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608763155
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1608763155
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608763155
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608763155
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 1608763155
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1608763155
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1608763155
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1608763155
transform 1 0 1932 0 1 2720
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 0 258 800 4 bottom_left_grid_pin_42_
port 1 nsew
rlabel metal2 s 662 0 718 800 4 bottom_left_grid_pin_43_
port 2 nsew
rlabel metal2 s 1122 0 1178 800 4 bottom_left_grid_pin_44_
port 3 nsew
rlabel metal2 s 1582 0 1638 800 4 bottom_left_grid_pin_45_
port 4 nsew
rlabel metal2 s 2042 0 2098 800 4 bottom_left_grid_pin_46_
port 5 nsew
rlabel metal2 s 2502 0 2558 800 4 bottom_left_grid_pin_47_
port 6 nsew
rlabel metal2 s 2962 0 3018 800 4 bottom_left_grid_pin_48_
port 7 nsew
rlabel metal2 s 3422 0 3478 800 4 bottom_left_grid_pin_49_
port 8 nsew
rlabel metal2 s 22466 0 22522 800 4 bottom_right_grid_pin_1_
port 9 nsew
rlabel metal3 s 22000 5720 22800 5840 4 ccff_head
port 10 nsew
rlabel metal3 s 22000 17144 22800 17264 4 ccff_tail
port 11 nsew
rlabel metal3 s 0 3952 800 4072 4 chanx_left_in[0]
port 12 nsew
rlabel metal3 s 0 8712 800 8832 4 chanx_left_in[10]
port 13 nsew
rlabel metal3 s 0 9120 800 9240 4 chanx_left_in[11]
port 14 nsew
rlabel metal3 s 0 9664 800 9784 4 chanx_left_in[12]
port 15 nsew
rlabel metal3 s 0 10072 800 10192 4 chanx_left_in[13]
port 16 nsew
rlabel metal3 s 0 10616 800 10736 4 chanx_left_in[14]
port 17 nsew
rlabel metal3 s 0 11024 800 11144 4 chanx_left_in[15]
port 18 nsew
rlabel metal3 s 0 11568 800 11688 4 chanx_left_in[16]
port 19 nsew
rlabel metal3 s 0 11976 800 12096 4 chanx_left_in[17]
port 20 nsew
rlabel metal3 s 0 12520 800 12640 4 chanx_left_in[18]
port 21 nsew
rlabel metal3 s 0 12928 800 13048 4 chanx_left_in[19]
port 22 nsew
rlabel metal3 s 0 4360 800 4480 4 chanx_left_in[1]
port 23 nsew
rlabel metal3 s 0 4904 800 5024 4 chanx_left_in[2]
port 24 nsew
rlabel metal3 s 0 5312 800 5432 4 chanx_left_in[3]
port 25 nsew
rlabel metal3 s 0 5856 800 5976 4 chanx_left_in[4]
port 26 nsew
rlabel metal3 s 0 6264 800 6384 4 chanx_left_in[5]
port 27 nsew
rlabel metal3 s 0 6808 800 6928 4 chanx_left_in[6]
port 28 nsew
rlabel metal3 s 0 7216 800 7336 4 chanx_left_in[7]
port 29 nsew
rlabel metal3 s 0 7760 800 7880 4 chanx_left_in[8]
port 30 nsew
rlabel metal3 s 0 8168 800 8288 4 chanx_left_in[9]
port 31 nsew
rlabel metal3 s 0 13472 800 13592 4 chanx_left_out[0]
port 32 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[10]
port 33 nsew
rlabel metal3 s 0 18640 800 18760 4 chanx_left_out[11]
port 34 nsew
rlabel metal3 s 0 19184 800 19304 4 chanx_left_out[12]
port 35 nsew
rlabel metal3 s 0 19592 800 19712 4 chanx_left_out[13]
port 36 nsew
rlabel metal3 s 0 20136 800 20256 4 chanx_left_out[14]
port 37 nsew
rlabel metal3 s 0 20544 800 20664 4 chanx_left_out[15]
port 38 nsew
rlabel metal3 s 0 21088 800 21208 4 chanx_left_out[16]
port 39 nsew
rlabel metal3 s 0 21496 800 21616 4 chanx_left_out[17]
port 40 nsew
rlabel metal3 s 0 22040 800 22160 4 chanx_left_out[18]
port 41 nsew
rlabel metal3 s 0 22448 800 22568 4 chanx_left_out[19]
port 42 nsew
rlabel metal3 s 0 13880 800 14000 4 chanx_left_out[1]
port 43 nsew
rlabel metal3 s 0 14424 800 14544 4 chanx_left_out[2]
port 44 nsew
rlabel metal3 s 0 14832 800 14952 4 chanx_left_out[3]
port 45 nsew
rlabel metal3 s 0 15376 800 15496 4 chanx_left_out[4]
port 46 nsew
rlabel metal3 s 0 15784 800 15904 4 chanx_left_out[5]
port 47 nsew
rlabel metal3 s 0 16328 800 16448 4 chanx_left_out[6]
port 48 nsew
rlabel metal3 s 0 16736 800 16856 4 chanx_left_out[7]
port 49 nsew
rlabel metal3 s 0 17280 800 17400 4 chanx_left_out[8]
port 50 nsew
rlabel metal3 s 0 17688 800 17808 4 chanx_left_out[9]
port 51 nsew
rlabel metal2 s 3882 0 3938 800 4 chany_bottom_in[0]
port 52 nsew
rlabel metal2 s 8574 0 8630 800 4 chany_bottom_in[10]
port 53 nsew
rlabel metal2 s 9034 0 9090 800 4 chany_bottom_in[11]
port 54 nsew
rlabel metal2 s 9494 0 9550 800 4 chany_bottom_in[12]
port 55 nsew
rlabel metal2 s 9954 0 10010 800 4 chany_bottom_in[13]
port 56 nsew
rlabel metal2 s 10414 0 10470 800 4 chany_bottom_in[14]
port 57 nsew
rlabel metal2 s 10874 0 10930 800 4 chany_bottom_in[15]
port 58 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_in[16]
port 59 nsew
rlabel metal2 s 11794 0 11850 800 4 chany_bottom_in[17]
port 60 nsew
rlabel metal2 s 12254 0 12310 800 4 chany_bottom_in[18]
port 61 nsew
rlabel metal2 s 12714 0 12770 800 4 chany_bottom_in[19]
port 62 nsew
rlabel metal2 s 4342 0 4398 800 4 chany_bottom_in[1]
port 63 nsew
rlabel metal2 s 4802 0 4858 800 4 chany_bottom_in[2]
port 64 nsew
rlabel metal2 s 5262 0 5318 800 4 chany_bottom_in[3]
port 65 nsew
rlabel metal2 s 5722 0 5778 800 4 chany_bottom_in[4]
port 66 nsew
rlabel metal2 s 6182 0 6238 800 4 chany_bottom_in[5]
port 67 nsew
rlabel metal2 s 6642 0 6698 800 4 chany_bottom_in[6]
port 68 nsew
rlabel metal2 s 7102 0 7158 800 4 chany_bottom_in[7]
port 69 nsew
rlabel metal2 s 7562 0 7618 800 4 chany_bottom_in[8]
port 70 nsew
rlabel metal2 s 8114 0 8170 800 4 chany_bottom_in[9]
port 71 nsew
rlabel metal2 s 13174 0 13230 800 4 chany_bottom_out[0]
port 72 nsew
rlabel metal2 s 17866 0 17922 800 4 chany_bottom_out[10]
port 73 nsew
rlabel metal2 s 18326 0 18382 800 4 chany_bottom_out[11]
port 74 nsew
rlabel metal2 s 18786 0 18842 800 4 chany_bottom_out[12]
port 75 nsew
rlabel metal2 s 19246 0 19302 800 4 chany_bottom_out[13]
port 76 nsew
rlabel metal2 s 19706 0 19762 800 4 chany_bottom_out[14]
port 77 nsew
rlabel metal2 s 20166 0 20222 800 4 chany_bottom_out[15]
port 78 nsew
rlabel metal2 s 20626 0 20682 800 4 chany_bottom_out[16]
port 79 nsew
rlabel metal2 s 21086 0 21142 800 4 chany_bottom_out[17]
port 80 nsew
rlabel metal2 s 21546 0 21602 800 4 chany_bottom_out[18]
port 81 nsew
rlabel metal2 s 22006 0 22062 800 4 chany_bottom_out[19]
port 82 nsew
rlabel metal2 s 13634 0 13690 800 4 chany_bottom_out[1]
port 83 nsew
rlabel metal2 s 14094 0 14150 800 4 chany_bottom_out[2]
port 84 nsew
rlabel metal2 s 14554 0 14610 800 4 chany_bottom_out[3]
port 85 nsew
rlabel metal2 s 15014 0 15070 800 4 chany_bottom_out[4]
port 86 nsew
rlabel metal2 s 15566 0 15622 800 4 chany_bottom_out[5]
port 87 nsew
rlabel metal2 s 16026 0 16082 800 4 chany_bottom_out[6]
port 88 nsew
rlabel metal2 s 16486 0 16542 800 4 chany_bottom_out[7]
port 89 nsew
rlabel metal2 s 16946 0 17002 800 4 chany_bottom_out[8]
port 90 nsew
rlabel metal2 s 17406 0 17462 800 4 chany_bottom_out[9]
port 91 nsew
rlabel metal2 s 3790 22000 3846 22800 4 chany_top_in[0]
port 92 nsew
rlabel metal2 s 8390 22000 8446 22800 4 chany_top_in[10]
port 93 nsew
rlabel metal2 s 8850 22000 8906 22800 4 chany_top_in[11]
port 94 nsew
rlabel metal2 s 9310 22000 9366 22800 4 chany_top_in[12]
port 95 nsew
rlabel metal2 s 9770 22000 9826 22800 4 chany_top_in[13]
port 96 nsew
rlabel metal2 s 10230 22000 10286 22800 4 chany_top_in[14]
port 97 nsew
rlabel metal2 s 10690 22000 10746 22800 4 chany_top_in[15]
port 98 nsew
rlabel metal2 s 11150 22000 11206 22800 4 chany_top_in[16]
port 99 nsew
rlabel metal2 s 11610 22000 11666 22800 4 chany_top_in[17]
port 100 nsew
rlabel metal2 s 11978 22000 12034 22800 4 chany_top_in[18]
port 101 nsew
rlabel metal2 s 12438 22000 12494 22800 4 chany_top_in[19]
port 102 nsew
rlabel metal2 s 4250 22000 4306 22800 4 chany_top_in[1]
port 103 nsew
rlabel metal2 s 4710 22000 4766 22800 4 chany_top_in[2]
port 104 nsew
rlabel metal2 s 5170 22000 5226 22800 4 chany_top_in[3]
port 105 nsew
rlabel metal2 s 5630 22000 5686 22800 4 chany_top_in[4]
port 106 nsew
rlabel metal2 s 6090 22000 6146 22800 4 chany_top_in[5]
port 107 nsew
rlabel metal2 s 6550 22000 6606 22800 4 chany_top_in[6]
port 108 nsew
rlabel metal2 s 7010 22000 7066 22800 4 chany_top_in[7]
port 109 nsew
rlabel metal2 s 7470 22000 7526 22800 4 chany_top_in[8]
port 110 nsew
rlabel metal2 s 7930 22000 7986 22800 4 chany_top_in[9]
port 111 nsew
rlabel metal2 s 12898 22000 12954 22800 4 chany_top_out[0]
port 112 nsew
rlabel metal2 s 17498 22000 17554 22800 4 chany_top_out[10]
port 113 nsew
rlabel metal2 s 17958 22000 18014 22800 4 chany_top_out[11]
port 114 nsew
rlabel metal2 s 18418 22000 18474 22800 4 chany_top_out[12]
port 115 nsew
rlabel metal2 s 18878 22000 18934 22800 4 chany_top_out[13]
port 116 nsew
rlabel metal2 s 19338 22000 19394 22800 4 chany_top_out[14]
port 117 nsew
rlabel metal2 s 19798 22000 19854 22800 4 chany_top_out[15]
port 118 nsew
rlabel metal2 s 20258 22000 20314 22800 4 chany_top_out[16]
port 119 nsew
rlabel metal2 s 20718 22000 20774 22800 4 chany_top_out[17]
port 120 nsew
rlabel metal2 s 21178 22000 21234 22800 4 chany_top_out[18]
port 121 nsew
rlabel metal2 s 21638 22000 21694 22800 4 chany_top_out[19]
port 122 nsew
rlabel metal2 s 13358 22000 13414 22800 4 chany_top_out[1]
port 123 nsew
rlabel metal2 s 13818 22000 13874 22800 4 chany_top_out[2]
port 124 nsew
rlabel metal2 s 14278 22000 14334 22800 4 chany_top_out[3]
port 125 nsew
rlabel metal2 s 14738 22000 14794 22800 4 chany_top_out[4]
port 126 nsew
rlabel metal2 s 15198 22000 15254 22800 4 chany_top_out[5]
port 127 nsew
rlabel metal2 s 15658 22000 15714 22800 4 chany_top_out[6]
port 128 nsew
rlabel metal2 s 16118 22000 16174 22800 4 chany_top_out[7]
port 129 nsew
rlabel metal2 s 16578 22000 16634 22800 4 chany_top_out[8]
port 130 nsew
rlabel metal2 s 17038 22000 17094 22800 4 chany_top_out[9]
port 131 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_34_
port 132 nsew
rlabel metal3 s 0 552 800 672 4 left_bottom_grid_pin_35_
port 133 nsew
rlabel metal3 s 0 1096 800 1216 4 left_bottom_grid_pin_36_
port 134 nsew
rlabel metal3 s 0 1504 800 1624 4 left_bottom_grid_pin_37_
port 135 nsew
rlabel metal3 s 0 2048 800 2168 4 left_bottom_grid_pin_38_
port 136 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_39_
port 137 nsew
rlabel metal3 s 0 3000 800 3120 4 left_bottom_grid_pin_40_
port 138 nsew
rlabel metal3 s 0 3408 800 3528 4 left_bottom_grid_pin_41_
port 139 nsew
rlabel metal2 s 22098 22000 22154 22800 4 prog_clk_0_N_in
port 140 nsew
rlabel metal2 s 202 22000 258 22800 4 top_left_grid_pin_42_
port 141 nsew
rlabel metal2 s 570 22000 626 22800 4 top_left_grid_pin_43_
port 142 nsew
rlabel metal2 s 1030 22000 1086 22800 4 top_left_grid_pin_44_
port 143 nsew
rlabel metal2 s 1490 22000 1546 22800 4 top_left_grid_pin_45_
port 144 nsew
rlabel metal2 s 1950 22000 2006 22800 4 top_left_grid_pin_46_
port 145 nsew
rlabel metal2 s 2410 22000 2466 22800 4 top_left_grid_pin_47_
port 146 nsew
rlabel metal2 s 2870 22000 2926 22800 4 top_left_grid_pin_48_
port 147 nsew
rlabel metal2 s 3330 22000 3386 22800 4 top_left_grid_pin_49_
port 148 nsew
rlabel metal2 s 22558 22000 22614 22800 4 top_right_grid_pin_1_
port 149 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 150 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 151 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_2__1_/results/magic/sb_2__1_.gds
string GDS_END 1232616
string GDS_START 78430
<< end >>
