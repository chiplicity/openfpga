* NGSPICE file created from cbx_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt cbx_1__1_ bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_11_ bottom_grid_pin_12_
+ bottom_grid_pin_13_ bottom_grid_pin_14_ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_
+ bottom_grid_pin_3_ bottom_grid_pin_4_ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_
+ bottom_grid_pin_8_ bottom_grid_pin_9_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ prog_clk VPWR VGND
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_8.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_13.mux_l3_in_0_ mux_top_ipin_13.mux_l2_in_1_/X mux_top_ipin_13.mux_l2_in_0_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_66_ chanx_left_in[5] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_6.mux_l1_in_0_/X mux_top_ipin_6.mux_l2_in_2_/S
+ mux_top_ipin_6.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_49_ chanx_right_in[2] chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_13.mux_l2_in_1_ chanx_left_in[9] chanx_right_in[3] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_1.mux_l1_in_0_/S
+ mux_top_ipin_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_65_ chanx_left_in[6] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_48_ chanx_right_in[3] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_13.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_13.mux_l1_in_0_/X mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_6.mux_l1_in_0_/S
+ mux_top_ipin_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_64_ chanx_left_in[7] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X bottom_grid_pin_4_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ chanx_right_in[4] chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_13.mux_l1_in_0_/S
+ mux_top_ipin_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ chanx_left_in[8] chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_46_ chanx_right_in[5] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_11.mux_l4_in_0_/X bottom_grid_pin_11_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l2_in_3_ _27_/HI chanx_right_in[14] mux_top_ipin_2.mux_l2_in_3_/S
+ mux_top_ipin_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_62_ chanx_left_in[9] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_45_ chanx_right_in[6] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_2.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_3_ _16_/HI chanx_right_in[17] mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_2.mux_l2_in_3_/S
+ mux_top_ipin_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S mux_top_ipin_7.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_61_ chanx_left_in[10] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ chanx_right_in[7] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_14.mux_l2_in_3_ _25_/HI chanx_right_in[18] mux_top_ipin_14.mux_l2_in_3_/S
+ mux_top_ipin_14.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_2.mux_l2_in_3_/S
+ mux_top_ipin_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_60_ chanx_left_in[11] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_14.mux_l4_in_0_ mux_top_ipin_14.mux_l3_in_1_/X mux_top_ipin_14.mux_l3_in_0_/X
+ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_14.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X bottom_grid_pin_7_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_43_ chanx_right_in[8] chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_14.mux_l3_in_1_ mux_top_ipin_14.mux_l2_in_3_/X mux_top_ipin_14.mux_l2_in_2_/X
+ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_1_/S
+ mux_top_ipin_7.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_14.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_14.mux_l2_in_3_/S
+ mux_top_ipin_14.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_2.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_2.mux_l1_in_0_/X mux_top_ipin_2.mux_l2_in_3_/S
+ mux_top_ipin_2.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_42_ chanx_right_in[9] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_14.mux_l3_in_0_ mux_top_ipin_14.mux_l2_in_1_/X mux_top_ipin_14.mux_l2_in_0_/X
+ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_1_/S mux_top_ipin_7.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_14.mux_l4_in_0_/X bottom_grid_pin_14_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_14.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_14.mux_l2_in_3_/S
+ mux_top_ipin_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_14.mux_l3_in_1_/S mux_top_ipin_14.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_1.mux_l2_in_2_/S mux_top_ipin_1.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_2.mux_l1_in_0_/S
+ mux_top_ipin_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_41_ chanx_right_in[10] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_11.mux_l2_in_3_/S mux_top_ipin_11.mux_l3_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_7.mux_l3_in_0_/S mux_top_ipin_7.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_14.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_14.mux_l1_in_0_/X mux_top_ipin_14.mux_l2_in_3_/S
+ mux_top_ipin_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X bottom_grid_pin_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_7.mux_l1_in_2_/S
+ mux_top_ipin_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_4.mux_l2_in_3_/S mux_top_ipin_4.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_14.mux_l2_in_3_/S mux_top_ipin_14.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_1.mux_l1_in_0_/S mux_top_ipin_1.mux_l2_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_40_ chanx_right_in[11] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_23_ _23_/HI _23_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_11.mux_l1_in_2_/S mux_top_ipin_11.mux_l2_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_7.mux_l2_in_1_/S mux_top_ipin_7.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_4.mux_l1_in_2_/S mux_top_ipin_4.mux_l2_in_3_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_14.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_14.mux_l1_in_0_/S
+ mux_top_ipin_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_14.mux_l1_in_0_/S mux_top_ipin_14.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_1_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_1.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_11.mux_l1_in_2_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_22_ _22_/HI _22_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_7.mux_l1_in_2_/S mux_top_ipin_7.mux_l2_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_4.mux_l1_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l2_in_3_ _28_/HI chanx_right_in[19] mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_21_ _21_/HI _21_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_7.mux_l1_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S mux_top_ipin_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_8.mux_l2_in_3_ _17_/HI chanx_right_in[18] mux_top_ipin_8.mux_l2_in_3_/S
+ mux_top_ipin_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_8.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_3_ _21_/HI chanx_right_in[14] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_20_ _20_/HI _20_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X bottom_grid_pin_3_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_10.mux_l4_in_0_ mux_top_ipin_10.mux_l3_in_1_/X mux_top_ipin_10.mux_l3_in_0_/X
+ mux_top_ipin_10.mux_l4_in_0_/S mux_top_ipin_10.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_8.mux_l2_in_3_/S
+ mux_top_ipin_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_3_ _26_/HI chanx_right_in[19] mux_top_ipin_15.mux_l2_in_2_/S
+ mux_top_ipin_15.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l3_in_1_ mux_top_ipin_10.mux_l2_in_3_/X mux_top_ipin_10.mux_l2_in_2_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_3_/S
+ mux_top_ipin_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_10.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_15.mux_l4_in_0_ mux_top_ipin_15.mux_l3_in_1_/X mux_top_ipin_15.mux_l3_in_0_/X
+ ccff_tail mux_top_ipin_15.mux_l4_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l3_in_1_ mux_top_ipin_15.mux_l2_in_3_/X mux_top_ipin_15.mux_l2_in_2_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_3_/S
+ mux_top_ipin_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_15.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[15] mux_top_ipin_15.mux_l2_in_2_/S
+ mux_top_ipin_15.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l3_in_0_ mux_top_ipin_10.mux_l2_in_1_/X mux_top_ipin_10.mux_l2_in_0_/X
+ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_3_/S mux_top_ipin_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_10.mux_l4_in_0_/X bottom_grid_pin_10_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_10.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_15.mux_l3_in_0_ mux_top_ipin_15.mux_l2_in_1_/X mux_top_ipin_15.mux_l2_in_0_/X
+ mux_top_ipin_15.mux_l3_in_1_/S mux_top_ipin_15.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_3_/S mux_top_ipin_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l2_in_1_ chanx_left_in[15] mux_top_ipin_15.mux_l1_in_2_/X mux_top_ipin_15.mux_l2_in_2_/S
+ mux_top_ipin_15.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_10.mux_l1_in_0_/X mux_top_ipin_10.mux_l2_in_3_/S
+ mux_top_ipin_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_3.mux_l1_in_0_/S
+ mux_top_ipin_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_15.mux_l2_in_0_ mux_top_ipin_15.mux_l1_in_1_/X mux_top_ipin_15.mux_l1_in_0_/X
+ mux_top_ipin_15.mux_l2_in_2_/S mux_top_ipin_15.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_8.mux_l1_in_0_/S
+ mux_top_ipin_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_15.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_10.mux_l1_in_0_/S
+ mux_top_ipin_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_59_ chanx_left_in[12] chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X bottom_grid_pin_6_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_15.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_15.mux_l1_in_2_/S
+ mux_top_ipin_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_58_ chanx_left_in[13] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_13.mux_l4_in_0_/X bottom_grid_pin_13_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_4.mux_l2_in_3_ _29_/HI chanx_right_in[14] mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ chanx_left_in[14] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_4.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_3_ _18_/HI chanx_right_in[13] mux_top_ipin_9.mux_l2_in_3_/S
+ mux_top_ipin_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_10.mux_l3_in_1_/S mux_top_ipin_10.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l4_in_0_ mux_top_ipin_9.mux_l3_in_1_/X mux_top_ipin_9.mux_l3_in_0_/X
+ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_3.mux_l3_in_1_/S mux_top_ipin_3.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ chanx_left_in[15] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_3_ _22_/HI chanx_right_in[15] mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_9.mux_l3_in_1_ mux_top_ipin_9.mux_l2_in_3_/X mux_top_ipin_9.mux_l2_in_2_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_39_ chanx_right_in[12] chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l4_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l4_in_0_ mux_top_ipin_11.mux_l3_in_1_/X mux_top_ipin_11.mux_l3_in_0_/X
+ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_11.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_9.mux_l2_in_2_ chanx_left_in[13] chanx_right_in[5] mux_top_ipin_9.mux_l2_in_3_/S
+ mux_top_ipin_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S mux_top_ipin_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_10.mux_l2_in_3_/S mux_top_ipin_10.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l3_in_1_ mux_top_ipin_11.mux_l2_in_3_/X mux_top_ipin_11.mux_l2_in_2_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_3_/S
+ mux_top_ipin_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_3.mux_l2_in_3_/S mux_top_ipin_3.mux_l3_in_1_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[11] mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_55_ chanx_left_in[16] chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_9.mux_l3_in_0_ mux_top_ipin_9.mux_l2_in_1_/X mux_top_ipin_9.mux_l2_in_0_/X
+ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_13.mux_l2_in_3_/S mux_top_ipin_13.mux_l3_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_38_ chanx_right_in[13] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_0.mux_l1_in_2_/S mux_top_ipin_0.mux_l2_in_2_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_9.mux_l4_in_0_/X bottom_grid_pin_9_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_9.mux_l3_in_1_/S mux_top_ipin_9.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_1_ chanx_left_in[5] chanx_right_in[3] mux_top_ipin_9.mux_l2_in_3_/S
+ mux_top_ipin_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_10.mux_l1_in_0_/S mux_top_ipin_10.mux_l2_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_6.mux_l2_in_2_/S mux_top_ipin_6.mux_l3_in_1_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_11.mux_l3_in_0_ mux_top_ipin_11.mux_l2_in_1_/X mux_top_ipin_11.mux_l2_in_0_/X
+ mux_top_ipin_11.mux_l3_in_1_/S mux_top_ipin_11.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_71_ chanx_left_in[0] chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_3_/S mux_top_ipin_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_3.mux_l1_in_0_/S mux_top_ipin_3.mux_l2_in_3_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_54_ chanx_left_in[17] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_11.mux_l1_in_2_/X mux_top_ipin_11.mux_l2_in_3_/S
+ mux_top_ipin_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_13.mux_l1_in_0_/S mux_top_ipin_13.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_37_ chanx_right_in[14] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_ipin_0.mux_l1_in_2_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_11.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_9.mux_l2_in_3_/S mux_top_ipin_9.mux_l3_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_9.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_9.mux_l1_in_0_/X mux_top_ipin_9.mux_l2_in_3_/S
+ mux_top_ipin_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_9.mux_l4_in_0_/S mux_top_ipin_10.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_6.mux_l1_in_0_/S mux_top_ipin_6.mux_l2_in_2_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ chanx_left_in[1] chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_2.mux_l4_in_0_/S mux_top_ipin_3.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_11.mux_l2_in_0_ mux_top_ipin_11.mux_l1_in_1_/X mux_top_ipin_11.mux_l1_in_0_/X
+ mux_top_ipin_11.mux_l2_in_3_/S mux_top_ipin_11.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_53_ chanx_left_in[18] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_4.mux_l1_in_2_/S
+ mux_top_ipin_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_13.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_36_ chanx_right_in[15] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_11.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19_ _19_/HI _19_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_9.mux_l1_in_0_/S mux_top_ipin_9.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_6.mux_l1_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_9.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_9.mux_l1_in_0_/S
+ mux_top_ipin_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X bottom_grid_pin_2_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ chanx_left_in[19] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_35_ chanx_right_in[16] chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_11.mux_l1_in_2_/S
+ mux_top_ipin_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18_ _18_/HI _18_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_8.mux_l4_in_0_/S mux_top_ipin_9.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_51_ chanx_right_in[0] chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_34_ chanx_right_in[17] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17_ _17_/HI _17_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l2_in_3_ _19_/HI chanx_right_in[16] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S mux_top_ipin_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_50_ chanx_right_in[1] chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_5.mux_l2_in_3_ _30_/HI chanx_right_in[17] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_33_ chanx_right_in[18] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_16_ _16_/HI _16_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S mux_top_ipin_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[9] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_32_ chanx_right_in[19] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S mux_top_ipin_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_12.mux_l2_in_3_ _23_/HI chanx_right_in[16] mux_top_ipin_12.mux_l2_in_3_/S
+ mux_top_ipin_12.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_2_/S
+ mux_top_ipin_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l4_in_0_ mux_top_ipin_12.mux_l3_in_1_/X mux_top_ipin_12.mux_l3_in_0_/X
+ mux_top_ipin_12.mux_l4_in_0_/S mux_top_ipin_12.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X bottom_grid_pin_5_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_12.mux_l3_in_1_ mux_top_ipin_12.mux_l2_in_3_/X mux_top_ipin_12.mux_l2_in_2_/X
+ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[9] chanx_right_in[3] mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_top_ipin_12.mux_l2_in_3_/S
+ mux_top_ipin_12.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_2_/S mux_top_ipin_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l3_in_0_ mux_top_ipin_12.mux_l2_in_1_/X mux_top_ipin_12.mux_l2_in_0_/X
+ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_5.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_5.mux_l1_in_0_/X mux_top_ipin_5.mux_l2_in_2_/S
+ mux_top_ipin_5.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_12.mux_l4_in_0_/X bottom_grid_pin_12_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_ipin_12.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_12.mux_l1_in_2_/X mux_top_ipin_12.mux_l2_in_3_/S
+ mux_top_ipin_12.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_12.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_0.mux_l1_in_2_/S
+ mux_top_ipin_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_12.mux_l2_in_0_ mux_top_ipin_12.mux_l1_in_1_/X mux_top_ipin_12.mux_l1_in_0_/X
+ mux_top_ipin_12.mux_l2_in_3_/S mux_top_ipin_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_5.mux_l1_in_0_/S
+ mux_top_ipin_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_12.mux_l1_in_2_/S
+ mux_top_ipin_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_2.mux_l3_in_1_/S mux_top_ipin_2.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_12.mux_l3_in_1_/S mux_top_ipin_12.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X bottom_grid_pin_8_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_5.mux_l3_in_0_/S mux_top_ipin_5.mux_l4_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_15.mux_l3_in_1_/S ccff_tail
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_2.mux_l2_in_3_/S mux_top_ipin_2.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _20_/HI chanx_right_in[13] mux_top_ipin_1.mux_l2_in_2_/S
+ mux_top_ipin_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_12.mux_l2_in_3_/S mux_top_ipin_12.mux_l3_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_ipin_8.mux_l3_in_0_/S mux_top_ipin_8.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_15.mux_l4_in_0_/X bottom_grid_pin_15_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_5.mux_l2_in_2_/S mux_top_ipin_5.mux_l3_in_0_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_69_ chanx_left_in[2] chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_3_ _31_/HI chanx_right_in[18] mux_top_ipin_6.mux_l2_in_2_/S
+ mux_top_ipin_6.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_15.mux_l2_in_2_/S mux_top_ipin_15.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_2.mux_l1_in_0_/S mux_top_ipin_2.mux_l2_in_3_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[13] chanx_right_in[5] mux_top_ipin_1.mux_l2_in_2_/S
+ mux_top_ipin_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S mux_top_ipin_6.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_12.mux_l1_in_2_/S mux_top_ipin_12.mux_l2_in_3_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_ipin_8.mux_l2_in_3_/S mux_top_ipin_8.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X bottom_grid_pin_1_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_5.mux_l1_in_0_/S mux_top_ipin_5.mux_l2_in_2_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_68_ chanx_left_in[3] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_6.mux_l2_in_2_/S
+ mux_top_ipin_6.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_0_/S mux_top_ipin_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_13.mux_l2_in_3_ _24_/HI chanx_right_in[17] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_15.mux_l1_in_2_/S mux_top_ipin_15.mux_l2_in_2_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_1.mux_l4_in_0_/S mux_top_ipin_2.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[5] chanx_right_in[3] mux_top_ipin_1.mux_l2_in_2_/S
+ mux_top_ipin_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_11.mux_l4_in_0_/S mux_top_ipin_12.mux_l1_in_2_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l4_in_0_ mux_top_ipin_13.mux_l3_in_1_/X mux_top_ipin_13.mux_l3_in_0_/X
+ mux_top_ipin_13.mux_l4_in_0_/S mux_top_ipin_13.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_ipin_8.mux_l1_in_0_/S mux_top_ipin_8.mux_l2_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S mux_top_ipin_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_13.mux_l3_in_1_ mux_top_ipin_13.mux_l2_in_3_/X mux_top_ipin_13.mux_l2_in_2_/X
+ mux_top_ipin_13.mux_l3_in_1_/S mux_top_ipin_13.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_4.mux_l4_in_0_/S mux_top_ipin_5.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_67_ chanx_left_in[4] chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_6.mux_l2_in_2_/S
+ mux_top_ipin_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_13.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[9] mux_top_ipin_13.mux_l2_in_3_/S
+ mux_top_ipin_13.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_ipin_14.mux_l4_in_0_/S mux_top_ipin_15.mux_l1_in_2_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_ipin_1.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_1.mux_l1_in_0_/X mux_top_ipin_1.mux_l2_in_2_/S
+ mux_top_ipin_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

