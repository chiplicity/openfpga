* NGSPICE file created from sb_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt sb_1__2_ bottom_left_grid_pin_34_ bottom_left_grid_pin_35_ bottom_left_grid_pin_36_
+ bottom_left_grid_pin_37_ bottom_left_grid_pin_38_ bottom_left_grid_pin_39_ bottom_left_grid_pin_40_
+ bottom_left_grid_pin_41_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_top_grid_pin_1_ prog_clk right_top_grid_pin_1_ VPWR VGND
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A0 bottom_left_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_3.mux_l1_in_3__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_7.mux_l2_in_1__S mux_bottom_track_7.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_114_ _114_/A chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l1_in_0_ bottom_left_grid_pin_38_ chanx_right_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_29.mux_l2_in_0_ _065_/HI mux_bottom_track_29.mux_l1_in_0_/X mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_1_/S mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__S mux_bottom_track_19.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_31.mux_l2_in_0_ _067_/HI mux_bottom_track_31.mux_l1_in_0_/X mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _126_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__127__A _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A1 chanx_right_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A mux_left_track_1.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l3_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l3_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ _113_/A chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_29.mux_l1_in_0_ bottom_left_grid_pin_36_ chanx_right_in[11] mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_31.mux_l1_in_0_ bottom_left_grid_pin_37_ chanx_right_in[7] mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_23.mux_l1_in_0__S mux_bottom_track_23.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_39.mux_l2_in_0__A1 mux_bottom_track_39.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l2_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_112_ _112_/A chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A0 _057_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_15.mux_l2_in_0__S mux_bottom_track_15.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A0 mux_bottom_track_13.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_11.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A0 bottom_left_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_1_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_111_ _111_/A chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A0 _061_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__072__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 mux_bottom_track_5.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A0 mux_bottom_track_21.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_1_ _054_/HI mux_right_track_8.mux_l1_in_2_/X mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_37.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A1 mux_bottom_track_13.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__080__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_2_ chanx_left_in[16] chanx_left_in[6] mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_110_ _110_/A chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l2_in_0_/S mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X
+ _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A1 mux_bottom_track_21.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_1_ chany_bottom_in[16] chany_bottom_in[9] mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0__S mux_bottom_track_11.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 bottom_left_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_11.mux_l3_in_0_/S
+ mux_bottom_track_13.mux_l1_in_1_/S mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 mux_right_track_8.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__094__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l2_in_0_/S mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S mux_bottom_track_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l1_in_0_ chany_bottom_in[2] right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_1_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__089__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chanx_right_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_13.mux_l1_in_1_ _057_/HI chanx_left_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_bottom_track_25.mux_l2_in_1_ _063_/HI chanx_left_in[18] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_099_ _099_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__097__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_1_ _040_/HI chanx_left_in[15] mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__S mux_bottom_track_37.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _091_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 bottom_left_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_1_/S mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A1 chanx_left_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_31.mux_l1_in_0_/S
+ mux_bottom_track_31.mux_l2_in_0_/S mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_13.mux_l1_in_0_ bottom_left_grid_pin_36_ chanx_right_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_35.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_25.mux_l2_in_0_ bottom_left_grid_pin_34_ mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__S mux_bottom_track_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_29.mux_l2_in_0__S mux_bottom_track_29.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_098_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ chanx_left_in[8] mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l3_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chanx_right_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A0 _060_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A0 mux_bottom_track_19.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_29.mux_l2_in_0_/S
+ mux_bottom_track_31.mux_l1_in_0_/S mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_2__S mux_right_track_8.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_097_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ chanx_right_in[19] chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/S mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_3.mux_l1_in_1_/S mux_left_track_3.mux_l2_in_1_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_37.mux_l2_in_0_ _036_/HI mux_bottom_track_37.mux_l1_in_0_/X mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A1 chanx_left_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A0 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[8] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _123_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l3_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A1 mux_bottom_track_19.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_1_ _044_/HI chany_bottom_in[14] mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A mux_left_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__100__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_096_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_7.mux_l1_in_1__S mux_bottom_track_7.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/S mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_3.mux_l1_in_1_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _079_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__S mux_bottom_track_19.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A1 mux_bottom_track_27.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_37.mux_l1_in_0_ bottom_left_grid_pin_40_ chanx_right_in[0] mux_bottom_track_37.mux_l1_in_0_/S
+ mux_bottom_track_37.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_1_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_31.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_1_ _049_/HI chanx_left_in[17] mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_4.mux_l2_in_1_ _053_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_1_/S
+ mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_095_ _095_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_right_track_0.mux_l1_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_35.mux_l2_in_0__A1 mux_bottom_track_35.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l3_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_33.mux_l2_in_1_/S ccff_tail
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_094_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2__A0 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_077_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__122__A _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_1_ chanx_left_in[8] chany_bottom_in[15] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_1_ chany_bottom_in[17] chany_bottom_in[10] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 bottom_left_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A0 chanx_left_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__S mux_bottom_track_21.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0__S mux_bottom_track_15.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/S mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_1_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 mux_bottom_track_1.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l3_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_3_ _038_/HI chanx_left_in[7] mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2__A1 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_076_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l1_in_0_ chany_bottom_in[8] chany_bottom_in[1] mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_bottom_in[3] right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_39.mux_l1_in_0__A1 bottom_left_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chanx_right_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 mux_left_track_9.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_35.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/S mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l2_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_092_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_29.mux_l1_in_0_/S
+ mux_bottom_track_29.mux_l2_in_0_/S mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A mux_left_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[5] bottom_left_grid_pin_40_ mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_075_ _075_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A0 bottom_left_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _099_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_127_ _127_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_7.mux_l2_in_1_/S
+ mux_bottom_track_7.mux_l3_in_0_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S mux_bottom_track_19.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S mux_bottom_track_21.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_39.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_39.mux_l2_in_0_/X
+ _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_bottom_track_19.mux_l1_in_1_ _060_/HI chanx_left_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A mux_left_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A0 _056_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_23.mux_l1_in_1__S mux_bottom_track_23.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_21.mux_l1_in_1_ _061_/HI chanx_left_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0__S mux_bottom_track_11.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_39.mux_l2_in_0__S mux_bottom_track_39.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X _087_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ _091_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_32.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l1_in_1_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A0 mux_bottom_track_11.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_29.mux_l1_in_0_/S mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A0 bottom_left_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_38_ bottom_left_grid_pin_36_
+ mux_bottom_track_5.mux_l1_in_1_/S mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A0 _066_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l2_in_1_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_126_ _126_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_7.mux_l3_in_0__S mux_bottom_track_7.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A mux_left_track_9.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _109_/A chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__070__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l1_in_0_ bottom_left_grid_pin_39_ chanx_right_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A1 chanx_left_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_21.mux_l1_in_0_ bottom_left_grid_pin_40_ chanx_right_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_33.mux_l2_in_0_ _034_/HI mux_bottom_track_33.mux_l1_in_0_/X mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_left_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A1 mux_bottom_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_090_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _125_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_1_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l3_in_0_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__073__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_39.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_125_ _125_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_7.mux_l1_in_2_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__068__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ _108_/A chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_7.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__081__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _071_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A0 _058_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__076__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_35.mux_l2_in_0__S mux_bottom_track_35.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_0_ bottom_left_grid_pin_38_ chanx_right_in[3] mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A0 mux_bottom_track_15.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_29.mux_l1_in_0__S mux_bottom_track_29.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_16.mux_l1_in_1_/S
+ mux_right_track_16.mux_l2_in_1_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_17.mux_l2_in_1_ _042_/HI chany_bottom_in[17] mux_left_track_17.mux_l2_in_1_/S
+ mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_124_ _124_/A chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__084__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_bottom_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l2_in_0_/S mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_107_ _107_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_1_ _047_/HI mux_left_track_9.mux_l1_in_2_/X mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__079__A _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_1_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__S mux_bottom_track_5.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_1_ _048_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A0 _062_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_1__S mux_bottom_track_11.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[16] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A1 chanx_left_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A0 mux_bottom_track_7.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_2_ chanx_left_in[12] chanx_left_in[2] mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A0 mux_bottom_track_23.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A1 mux_bottom_track_15.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A0 mux_bottom_track_7.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_8.mux_l3_in_0_/S mux_right_track_16.mux_l1_in_1_/S
+ mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__dfxbp_1
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _123_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_1_/S mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_106_ _106_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_1_ chany_bottom_in[10] chany_bottom_in[3] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A1 bottom_left_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_37.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A0 _067_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_31.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_1_ chany_bottom_in[9] chany_bottom_in[2] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A1 mux_bottom_track_7.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A1 mux_bottom_track_23.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_1_ chany_bottom_in[19] chany_bottom_in[12] mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_24.mux_l2_in_1_ _051_/HI chanx_left_in[18] mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_070_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A1 mux_bottom_track_7.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_31.mux_l2_in_0__S mux_bottom_track_31.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__098__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A0 bottom_left_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_122_ _122_/A chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_105_ _105_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chanx_right_in[17] chanx_right_in[8] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A mux_left_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_31.mux_l2_in_0__A1 mux_bottom_track_31.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _107_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_3_ _055_/HI chanx_left_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_3__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ chany_bottom_in[5] right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_29.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A0 bottom_left_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_33.mux_l1_in_0_/S
+ mux_bottom_track_33.mux_l2_in_0_/S mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_37.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_1_ chanx_left_in[9] chany_bottom_in[14] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_121_ _121_/A chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _063_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_40_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A0 bottom_left_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S mux_bottom_track_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_35.mux_l2_in_0_/X
+ _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_31.mux_l2_in_0_/S
+ mux_bottom_track_33.mux_l1_in_0_/S mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ chany_bottom_in[7] chany_bottom_in[0] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ _120_/A chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_15.mux_l1_in_1_ _058_/HI chanx_left_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_29.mux_l2_in_0_/X
+ _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_103_ _103_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_17.mux_l2_in_1_/S mux_left_track_17.mux_l3_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/S mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_5.mux_l1_in_2_/S mux_left_track_5.mux_l2_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__S mux_bottom_track_21.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_38_ bottom_left_grid_pin_36_
+ mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_35.mux_l1_in_0__A1 chanx_right_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__101__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_7.mux_l1_in_2__S mux_bottom_track_7.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_15.mux_l1_in_0_ bottom_left_grid_pin_37_ chanx_right_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.mux_l2_in_0_ _064_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0__S mux_bottom_track_13.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _127_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_102_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_1_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_37.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/S mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l1_in_1__S mux_bottom_track_19.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_2_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__104__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_34_ chanx_right_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A0 _065_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 mux_left_track_9.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_9.mux_l3_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__120__A _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[15] mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_39.mux_l2_in_0_ _037_/HI mux_bottom_track_39.mux_l1_in_0_/X mux_bottom_track_39.mux_l2_in_0_/S
+ mux_bottom_track_39.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_8.mux_l1_in_1_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_39.mux_l1_in_0__S mux_bottom_track_39.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_29.mux_l2_in_0__A1 mux_bottom_track_29.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_1_ _046_/HI mux_left_track_5.mux_l1_in_2_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_100_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_left_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__118__A _118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[15] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__S mux_bottom_track_7.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_1__S mux_bottom_track_15.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_37.mux_l2_in_0__A1 mux_bottom_track_37.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_1_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_39.mux_l1_in_0_ chanx_left_in[0] bottom_left_grid_pin_41_ mux_bottom_track_39.mux_l1_in_0_/S
+ mux_bottom_track_39.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__126__A _126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_1_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_29.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ _043_/HI chany_bottom_in[18] mux_left_track_25.mux_l2_in_1_/S
+ mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l3_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A0 chanx_left_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_35.mux_l1_in_0__S mux_bottom_track_35.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l2_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 mux_bottom_track_3.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S mux_bottom_track_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A mux_left_track_5.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_0_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l1_in_2_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l1_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_089_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A1 mux_bottom_track_11.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.mux_l2_in_1_ _056_/HI chanx_left_in[19] mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l3_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_27.mux_l2_in_0__S mux_bottom_track_27.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 bottom_left_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_1_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 mux_bottom_track_3.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_0_ chanx_right_in[18] chanx_right_in[9] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l3_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_088_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_31.mux_l2_in_0_/X
+ _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_7.mux_l1_in_3_ _039_/HI chanx_left_in[11] mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.mux_l2_in_0_ chanx_left_in[9] mux_bottom_track_11.mux_l1_in_0_/X
+ mux_bottom_track_11.mux_l2_in_0_/S mux_bottom_track_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_1_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A0 bottom_left_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_37.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_35.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ _118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_1_ _052_/HI chanx_left_in[10] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_31.mux_l1_in_0__S mux_bottom_track_31.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__074__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_087_ _087_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__069__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A0 bottom_left_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A0 bottom_left_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _095_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
Xmux_bottom_track_7.mux_l1_in_2_ chanx_left_in[6] bottom_left_grid_pin_41_ mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_7.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A1 chanx_right_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A0 mux_bottom_track_7.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__082__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_11.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[9] mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S mux_bottom_track_23.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__077__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_9.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_29.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[13] chany_bottom_in[6] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_23.mux_l2_in_0__S mux_bottom_track_23.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.mux_l1_in_1_ _062_/HI chanx_left_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A0 bottom_left_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__090__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _086_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A1 bottom_left_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_7.mux_l1_in_2_/S mux_bottom_track_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l2_in_0_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A1 mux_bottom_track_7.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__088__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l1_in_0_ bottom_left_grid_pin_41_ chanx_right_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_35.mux_l2_in_0_ _035_/HI mux_bottom_track_35.mux_l1_in_0_/X mux_bottom_track_35.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_31.mux_l1_in_0__A1 chanx_right_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_085_ _085_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 _059_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_35_ chanx_right_in[6] mux_bottom_track_7.mux_l1_in_2_/S
+ mux_bottom_track_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _124_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__096__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_39.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ _041_/HI left_top_grid_pin_1_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_39.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_33.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_084_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 bottom_left_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0__S mux_bottom_track_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/HI _067_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_35.mux_l1_in_0_ bottom_left_grid_pin_39_ chanx_right_in[1] mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_119_ _119_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_31.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_1_ _050_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_11.mux_l3_in_0__S mux_bottom_track_11.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 chanx_left_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_35.mux_l1_in_0_/S
+ mux_bottom_track_35.mux_l2_in_0_/S mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_1.mux_l1_in_1_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_39.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_39.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_066_ _066_/HI _066_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ _118_/A chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l1_in_1_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l2_in_1_ _045_/HI chany_bottom_in[19] mux_left_track_33.mux_l2_in_1_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_1_ chanx_left_in[4] chany_bottom_in[18] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_33.mux_l2_in_0_/S
+ mux_bottom_track_35.mux_l1_in_0_/S mem_bottom_track_35.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_39.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_1_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A0 bottom_left_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_1__S mux_bottom_track_21.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__S mux_bottom_track_7.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_117_ _117_/A chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_37.mux_l2_in_0__S mux_bottom_track_37.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l2_in_0_ chany_bottom_in[12] mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l1_in_3_ _066_/HI chanx_left_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _106_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__S mux_bottom_track_7.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_081_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l1_in_0_ chany_bottom_in[11] chany_bottom_in[4] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A0 bottom_left_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_29.mux_l1_in_0__A1 chanx_right_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l2_in_1_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_116_ _116_/A chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_41_ mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_0_ chany_bottom_in[5] chanx_right_in[10] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_37.mux_l1_in_0__A1 chanx_right_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__108__A _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_37.mux_l2_in_0_/X
+ _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_2_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_115_ _115_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l1_in_1_ _059_/HI chanx_left_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK prog_clk VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l2_in_0_/S mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S mux_bottom_track_33.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_27.mux_l1_in_0__S mux_bottom_track_27.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

