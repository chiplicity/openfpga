VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_top
  CLASS BLOCK ;
  FOREIGN grid_io_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2120.000 BY 50.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 47.600 132.850 50.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 10.920 2120.000 11.520 ;
    END
  END address[3]
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 15.680 2120.000 16.280 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 24.520 2120.000 25.120 ;
    END
  END bottom_width_0_height_0__pin_10_
  PIN bottom_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1192.410 47.600 1192.690 50.000 ;
    END
  END bottom_width_0_height_0__pin_11_
  PIN bottom_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END bottom_width_0_height_0__pin_12_
  PIN bottom_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 2.400 ;
    END
  END bottom_width_0_height_0__pin_13_
  PIN bottom_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 29.280 2120.000 29.880 ;
    END
  END bottom_width_0_height_0__pin_14_
  PIN bottom_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2117.600 34.040 2120.000 34.640 ;
    END
  END bottom_width_0_height_0__pin_15_
  PIN bottom_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 397.530 47.600 397.810 50.000 ;
    END
  END bottom_width_0_height_0__pin_1_
  PIN bottom_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 2.400 ;
    END
  END bottom_width_0_height_0__pin_2_
  PIN bottom_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2117.600 19.760 2120.000 20.360 ;
    END
  END bottom_width_0_height_0__pin_3_
  PIN bottom_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END bottom_width_0_height_0__pin_4_
  PIN bottom_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.400 21.040 ;
    END
  END bottom_width_0_height_0__pin_5_
  PIN bottom_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END bottom_width_0_height_0__pin_6_
  PIN bottom_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END bottom_width_0_height_0__pin_7_
  PIN bottom_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 47.600 662.770 50.000 ;
    END
  END bottom_width_0_height_0__pin_8_
  PIN bottom_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 927.450 47.600 927.730 50.000 ;
    END
  END bottom_width_0_height_0__pin_9_
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 6.160 2120.000 6.760 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 2.080 2120.000 2.680 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 38.120 2120.000 38.720 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1457.370 47.600 1457.650 50.000 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 42.880 2120.000 43.480 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1722.330 47.600 1722.610 50.000 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1483.590 0.000 1483.870 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 47.640 2120.000 48.240 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1907.710 0.000 1907.990 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1987.290 47.600 1987.570 50.000 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 358.055 10.640 359.655 38.320 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 711.385 10.640 712.985 38.320 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2114.160 38.165 ;
      LAYER met1 ;
        RECT 0.070 10.640 2118.690 41.440 ;
      LAYER met2 ;
        RECT 0.090 47.320 132.290 48.125 ;
        RECT 133.130 47.320 397.250 48.125 ;
        RECT 398.090 47.320 662.210 48.125 ;
        RECT 663.050 47.320 927.170 48.125 ;
        RECT 928.010 47.320 1192.130 48.125 ;
        RECT 1192.970 47.320 1457.090 48.125 ;
        RECT 1457.930 47.320 1722.050 48.125 ;
        RECT 1722.890 47.320 1987.010 48.125 ;
        RECT 1987.850 47.320 2118.670 48.125 ;
        RECT 0.090 2.680 2118.670 47.320 ;
        RECT 0.090 0.155 211.410 2.680 ;
        RECT 212.250 0.155 635.070 2.680 ;
        RECT 635.910 0.155 1059.190 2.680 ;
        RECT 1060.030 0.155 1483.310 2.680 ;
        RECT 1484.150 0.155 1907.430 2.680 ;
        RECT 1908.270 0.155 2118.670 2.680 ;
      LAYER met3 ;
        RECT 0.310 42.480 2117.200 43.330 ;
        RECT 0.310 39.120 2118.450 42.480 ;
        RECT 0.310 38.440 2117.200 39.120 ;
        RECT 2.800 37.720 2117.200 38.440 ;
        RECT 2.800 37.040 2118.450 37.720 ;
        RECT 0.310 35.040 2118.450 37.040 ;
        RECT 0.310 33.640 2117.200 35.040 ;
        RECT 0.310 30.280 2118.450 33.640 ;
        RECT 2.800 28.880 2117.200 30.280 ;
        RECT 0.310 25.520 2118.450 28.880 ;
        RECT 0.310 24.120 2117.200 25.520 ;
        RECT 0.310 21.440 2118.450 24.120 ;
        RECT 2.800 20.760 2118.450 21.440 ;
        RECT 2.800 20.040 2117.200 20.760 ;
        RECT 0.310 19.360 2117.200 20.040 ;
        RECT 0.310 16.680 2118.450 19.360 ;
        RECT 0.310 15.280 2117.200 16.680 ;
        RECT 0.310 13.280 2118.450 15.280 ;
        RECT 2.800 11.920 2118.450 13.280 ;
        RECT 2.800 11.880 2117.200 11.920 ;
        RECT 0.310 10.520 2117.200 11.880 ;
        RECT 0.310 7.160 2118.450 10.520 ;
        RECT 0.310 5.760 2117.200 7.160 ;
        RECT 0.310 5.120 2118.450 5.760 ;
        RECT 2.800 3.720 2118.450 5.120 ;
        RECT 0.310 3.080 2118.450 3.720 ;
        RECT 0.310 1.680 2117.200 3.080 ;
        RECT 0.310 0.175 2118.450 1.680 ;
      LAYER met4 ;
        RECT 358.050 38.720 2118.465 43.345 ;
        RECT 360.055 10.240 710.985 38.720 ;
        RECT 713.385 10.240 2118.465 38.720 ;
        RECT 358.050 0.175 2118.465 10.240 ;
      LAYER met5 ;
        RECT 635.380 11.100 1084.100 12.700 ;
  END
END grid_io_top
END LIBRARY

