magic
tech sky130A
magscale 1 2
timestamp 1604667938
<< viali >>
rect 3341 32521 3375 32555
rect 4997 32521 5031 32555
rect 7481 32521 7515 32555
rect 9321 32521 9355 32555
rect 13093 32521 13127 32555
rect 3157 32317 3191 32351
rect 3709 32317 3743 32351
rect 4813 32317 4847 32351
rect 5365 32317 5399 32351
rect 6837 32317 6871 32351
rect 8677 32317 8711 32351
rect 12449 32317 12483 32351
rect 7021 32181 7055 32215
rect 8861 32181 8895 32215
rect 12633 32181 12667 32215
rect 1777 31977 1811 32011
rect 2881 31977 2915 32011
rect 4261 31977 4295 32011
rect 5365 31977 5399 32011
rect 6837 31977 6871 32011
rect 8033 31977 8067 32011
rect 9873 31977 9907 32011
rect 12449 31977 12483 32011
rect 1593 31841 1627 31875
rect 2697 31841 2731 31875
rect 4077 31841 4111 31875
rect 5181 31841 5215 31875
rect 6653 31841 6687 31875
rect 7849 31841 7883 31875
rect 9689 31841 9723 31875
rect 12265 31841 12299 31875
rect 13369 31841 13403 31875
rect 13553 31637 13587 31671
rect 2881 31433 2915 31467
rect 7021 31433 7055 31467
rect 8861 31433 8895 31467
rect 9689 31433 9723 31467
rect 13369 31433 13403 31467
rect 3985 31365 4019 31399
rect 5825 31365 5859 31399
rect 12633 31365 12667 31399
rect 2697 31229 2731 31263
rect 3801 31229 3835 31263
rect 5641 31229 5675 31263
rect 6653 31229 6687 31263
rect 6837 31229 6871 31263
rect 8677 31229 8711 31263
rect 9781 31229 9815 31263
rect 12265 31229 12299 31263
rect 12449 31229 12483 31263
rect 1593 31093 1627 31127
rect 2513 31093 2547 31127
rect 3249 31093 3283 31127
rect 3617 31093 3651 31127
rect 4353 31093 4387 31127
rect 5181 31093 5215 31127
rect 6193 31093 6227 31127
rect 7389 31093 7423 31127
rect 7849 31093 7883 31127
rect 9321 31093 9355 31127
rect 9965 31093 9999 31127
rect 10425 31093 10459 31127
rect 13001 31093 13035 31127
rect 9965 30889 9999 30923
rect 11069 30889 11103 30923
rect 4353 30753 4387 30787
rect 9781 30753 9815 30787
rect 10885 30753 10919 30787
rect 4537 30549 4571 30583
rect 4353 30345 4387 30379
rect 9689 30277 9723 30311
rect 10793 30277 10827 30311
rect 9781 30141 9815 30175
rect 10885 30141 10919 30175
rect 9965 30005 9999 30039
rect 10425 30005 10459 30039
rect 11069 30005 11103 30039
rect 11437 30005 11471 30039
rect 10241 29665 10275 29699
rect 10425 29461 10459 29495
rect 10149 29257 10183 29291
rect 10425 29189 10459 29223
rect 10241 29053 10275 29087
rect 10793 29053 10827 29087
rect 1593 27081 1627 27115
rect 1409 26877 1443 26911
rect 1961 26741 1995 26775
rect 7113 26741 7147 26775
rect 7297 26537 7331 26571
rect 7205 26401 7239 26435
rect 7481 26333 7515 26367
rect 5089 26265 5123 26299
rect 6837 26265 6871 26299
rect 6285 25993 6319 26027
rect 6837 25925 6871 25959
rect 5457 25857 5491 25891
rect 5549 25857 5583 25891
rect 7297 25857 7331 25891
rect 7481 25857 7515 25891
rect 5365 25789 5399 25823
rect 4813 25721 4847 25755
rect 4997 25653 5031 25687
rect 6653 25653 6687 25687
rect 7205 25653 7239 25687
rect 7849 25653 7883 25687
rect 3157 25449 3191 25483
rect 5089 25449 5123 25483
rect 7205 25449 7239 25483
rect 12265 25449 12299 25483
rect 6929 25381 6963 25415
rect 12081 25313 12115 25347
rect 7573 25109 7607 25143
rect 3617 24769 3651 24803
rect 3433 24701 3467 24735
rect 2881 24565 2915 24599
rect 3065 24565 3099 24599
rect 3525 24565 3559 24599
rect 12081 24565 12115 24599
rect 3157 24021 3191 24055
rect 4537 21845 4571 21879
rect 4445 21641 4479 21675
rect 4353 21505 4387 21539
rect 5089 21505 5123 21539
rect 4813 21437 4847 21471
rect 4905 21301 4939 21335
rect 6009 21097 6043 21131
rect 6377 21029 6411 21063
rect 6469 20961 6503 20995
rect 6561 20893 6595 20927
rect 4537 20757 4571 20791
rect 6101 20553 6135 20587
rect 9689 20485 9723 20519
rect 6469 20417 6503 20451
rect 2973 20349 3007 20383
rect 3065 20349 3099 20383
rect 5733 20349 5767 20383
rect 8309 20349 8343 20383
rect 3332 20281 3366 20315
rect 8576 20281 8610 20315
rect 4445 20213 4479 20247
rect 8217 20213 8251 20247
rect 3157 20009 3191 20043
rect 5549 20009 5583 20043
rect 7113 20009 7147 20043
rect 7573 20009 7607 20043
rect 5917 19941 5951 19975
rect 7481 19941 7515 19975
rect 9956 19941 9990 19975
rect 6929 19873 6963 19907
rect 6009 19805 6043 19839
rect 6193 19805 6227 19839
rect 7757 19805 7791 19839
rect 9689 19805 9723 19839
rect 8401 19669 8435 19703
rect 11069 19669 11103 19703
rect 3893 19465 3927 19499
rect 7849 19465 7883 19499
rect 8309 19465 8343 19499
rect 6837 19397 6871 19431
rect 3985 19329 4019 19363
rect 7481 19329 7515 19363
rect 3525 19261 3559 19295
rect 4252 19261 4286 19295
rect 7205 19261 7239 19295
rect 6561 19193 6595 19227
rect 7297 19193 7331 19227
rect 5365 19125 5399 19159
rect 6193 19125 6227 19159
rect 9689 19125 9723 19159
rect 10057 19125 10091 19159
rect 5549 18921 5583 18955
rect 6009 18921 6043 18955
rect 6285 18921 6319 18955
rect 6469 18921 6503 18955
rect 7573 18921 7607 18955
rect 6837 18785 6871 18819
rect 6929 18717 6963 18751
rect 7021 18717 7055 18751
rect 6101 18377 6135 18411
rect 7021 18105 7055 18139
rect 6469 18037 6503 18071
rect 11529 13481 11563 13515
rect 10405 13345 10439 13379
rect 10149 13277 10183 13311
rect 10057 12937 10091 12971
rect 10609 12801 10643 12835
rect 10517 12733 10551 12767
rect 9229 12665 9263 12699
rect 9597 12597 9631 12631
rect 9873 12597 9907 12631
rect 10425 12597 10459 12631
rect 10057 12393 10091 12427
rect 8493 12053 8527 12087
rect 10425 12053 10459 12087
rect 8401 11849 8435 11883
rect 8309 11713 8343 11747
rect 9045 11713 9079 11747
rect 7941 11577 7975 11611
rect 8769 11577 8803 11611
rect 8861 11509 8895 11543
rect 6929 10965 6963 10999
rect 8493 10965 8527 10999
rect 6837 10761 6871 10795
rect 8309 10761 8343 10795
rect 8401 10761 8435 10795
rect 6653 10625 6687 10659
rect 7481 10625 7515 10659
rect 8953 10625 8987 10659
rect 7205 10557 7239 10591
rect 8769 10557 8803 10591
rect 7297 10421 7331 10455
rect 8861 10421 8895 10455
rect 5549 10217 5583 10251
rect 7113 10217 7147 10251
rect 5917 10149 5951 10183
rect 6009 10149 6043 10183
rect 6929 10149 6963 10183
rect 7481 10149 7515 10183
rect 6193 10013 6227 10047
rect 7573 10013 7607 10047
rect 7665 10013 7699 10047
rect 8493 9877 8527 9911
rect 5917 9673 5951 9707
rect 7481 9673 7515 9707
rect 5641 9605 5675 9639
rect 7849 9401 7883 9435
rect 6377 9333 6411 9367
rect 7113 9333 7147 9367
rect 5825 9129 5859 9163
rect 6285 9129 6319 9163
rect 6193 8993 6227 9027
rect 6469 8925 6503 8959
rect 5917 8585 5951 8619
rect 6193 8381 6227 8415
rect 6653 8313 6687 8347
rect 4333 6817 4367 6851
rect 4077 6749 4111 6783
rect 5457 6613 5491 6647
rect 10057 6613 10091 6647
rect 4169 6409 4203 6443
rect 9965 6409 9999 6443
rect 4445 6341 4479 6375
rect 9873 6273 9907 6307
rect 10609 6273 10643 6307
rect 9505 6137 9539 6171
rect 10333 6137 10367 6171
rect 10425 6069 10459 6103
rect 11069 5865 11103 5899
rect 9956 5729 9990 5763
rect 9689 5661 9723 5695
rect 6561 5321 6595 5355
rect 8217 5321 8251 5355
rect 8953 5321 8987 5355
rect 9873 5321 9907 5355
rect 6837 5185 6871 5219
rect 10425 5185 10459 5219
rect 10885 5185 10919 5219
rect 9321 5117 9355 5151
rect 10333 5117 10367 5151
rect 7082 5049 7116 5083
rect 9781 4981 9815 5015
rect 10241 4981 10275 5015
rect 6929 4777 6963 4811
rect 9965 4777 9999 4811
rect 10241 4777 10275 4811
rect 10701 4777 10735 4811
rect 10609 4641 10643 4675
rect 10793 4573 10827 4607
rect 9965 4233 9999 4267
rect 10333 4233 10367 4267
rect 10517 4097 10551 4131
rect 10977 4097 11011 4131
rect 4077 3553 4111 3587
rect 5181 3553 5215 3587
rect 4261 3417 4295 3451
rect 5365 3349 5399 3383
rect 3525 3145 3559 3179
rect 4169 3145 4203 3179
rect 4997 3145 5031 3179
rect 5733 3145 5767 3179
rect 7481 3145 7515 3179
rect 5273 3077 5307 3111
rect 6101 3009 6135 3043
rect 2881 2941 2915 2975
rect 3985 2941 4019 2975
rect 5089 2941 5123 2975
rect 6837 2941 6871 2975
rect 4629 2873 4663 2907
rect 3065 2805 3099 2839
rect 7021 2805 7055 2839
rect 2329 2601 2363 2635
rect 3065 2601 3099 2635
rect 4261 2601 4295 2635
rect 4721 2601 4755 2635
rect 5825 2601 5859 2635
rect 7389 2601 7423 2635
rect 7849 2601 7883 2635
rect 8953 2601 8987 2635
rect 3525 2533 3559 2567
rect 1685 2465 1719 2499
rect 2881 2465 2915 2499
rect 4077 2465 4111 2499
rect 5181 2465 5215 2499
rect 7205 2465 7239 2499
rect 8309 2465 8343 2499
rect 5365 2329 5399 2363
rect 8493 2329 8527 2363
rect 1869 2261 1903 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 2130 35640 2136 35692
rect 2188 35680 2194 35692
rect 2682 35680 2688 35692
rect 2188 35652 2688 35680
rect 2188 35640 2194 35652
rect 2682 35640 2688 35652
rect 2740 35640 2746 35692
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 198 34892 204 34944
rect 256 34932 262 34944
rect 1302 34932 1308 34944
rect 256 34904 1308 34932
rect 256 34892 262 34904
rect 1302 34892 1308 34904
rect 1360 34892 1366 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 4154 34688 4160 34740
rect 4212 34728 4218 34740
rect 5442 34728 5448 34740
rect 4212 34700 5448 34728
rect 4212 34688 4218 34700
rect 5442 34688 5448 34700
rect 5500 34688 5506 34740
rect 1394 34484 1400 34536
rect 1452 34524 1458 34536
rect 2774 34524 2780 34536
rect 1452 34496 2780 34524
rect 1452 34484 1458 34496
rect 2774 34484 2780 34496
rect 2832 34484 2838 34536
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 2774 32512 2780 32564
rect 2832 32552 2838 32564
rect 3329 32555 3387 32561
rect 3329 32552 3341 32555
rect 2832 32524 3341 32552
rect 2832 32512 2838 32524
rect 3329 32521 3341 32524
rect 3375 32521 3387 32555
rect 3329 32515 3387 32521
rect 4522 32512 4528 32564
rect 4580 32552 4586 32564
rect 4985 32555 5043 32561
rect 4985 32552 4997 32555
rect 4580 32524 4997 32552
rect 4580 32512 4586 32524
rect 4985 32521 4997 32524
rect 5031 32521 5043 32555
rect 7466 32552 7472 32564
rect 7427 32524 7472 32552
rect 4985 32515 5043 32521
rect 7466 32512 7472 32524
rect 7524 32512 7530 32564
rect 9306 32552 9312 32564
rect 9267 32524 9312 32552
rect 9306 32512 9312 32524
rect 9364 32512 9370 32564
rect 13078 32552 13084 32564
rect 13039 32524 13084 32552
rect 13078 32512 13084 32524
rect 13136 32512 13142 32564
rect 3142 32348 3148 32360
rect 3055 32320 3148 32348
rect 3142 32308 3148 32320
rect 3200 32348 3206 32360
rect 3697 32351 3755 32357
rect 3697 32348 3709 32351
rect 3200 32320 3709 32348
rect 3200 32308 3206 32320
rect 3697 32317 3709 32320
rect 3743 32317 3755 32351
rect 3697 32311 3755 32317
rect 4801 32351 4859 32357
rect 4801 32317 4813 32351
rect 4847 32348 4859 32351
rect 5074 32348 5080 32360
rect 4847 32320 5080 32348
rect 4847 32317 4859 32320
rect 4801 32311 4859 32317
rect 5074 32308 5080 32320
rect 5132 32348 5138 32360
rect 5353 32351 5411 32357
rect 5353 32348 5365 32351
rect 5132 32320 5365 32348
rect 5132 32308 5138 32320
rect 5353 32317 5365 32320
rect 5399 32317 5411 32351
rect 5353 32311 5411 32317
rect 6825 32351 6883 32357
rect 6825 32317 6837 32351
rect 6871 32348 6883 32351
rect 7466 32348 7472 32360
rect 6871 32320 7472 32348
rect 6871 32317 6883 32320
rect 6825 32311 6883 32317
rect 7466 32308 7472 32320
rect 7524 32308 7530 32360
rect 8665 32351 8723 32357
rect 8665 32317 8677 32351
rect 8711 32348 8723 32351
rect 9306 32348 9312 32360
rect 8711 32320 9312 32348
rect 8711 32317 8723 32320
rect 8665 32311 8723 32317
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 12437 32351 12495 32357
rect 12437 32317 12449 32351
rect 12483 32348 12495 32351
rect 13078 32348 13084 32360
rect 12483 32320 13084 32348
rect 12483 32317 12495 32320
rect 12437 32311 12495 32317
rect 13078 32308 13084 32320
rect 13136 32308 13142 32360
rect 7006 32212 7012 32224
rect 6967 32184 7012 32212
rect 7006 32172 7012 32184
rect 7064 32172 7070 32224
rect 7650 32172 7656 32224
rect 7708 32212 7714 32224
rect 8849 32215 8907 32221
rect 8849 32212 8861 32215
rect 7708 32184 8861 32212
rect 7708 32172 7714 32184
rect 8849 32181 8861 32184
rect 8895 32181 8907 32215
rect 12618 32212 12624 32224
rect 12579 32184 12624 32212
rect 8849 32175 8907 32181
rect 12618 32172 12624 32184
rect 12676 32172 12682 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1394 31968 1400 32020
rect 1452 32008 1458 32020
rect 1765 32011 1823 32017
rect 1765 32008 1777 32011
rect 1452 31980 1777 32008
rect 1452 31968 1458 31980
rect 1765 31977 1777 31980
rect 1811 31977 1823 32011
rect 2866 32008 2872 32020
rect 2827 31980 2872 32008
rect 1765 31971 1823 31977
rect 2866 31968 2872 31980
rect 2924 31968 2930 32020
rect 4246 32008 4252 32020
rect 4207 31980 4252 32008
rect 4246 31968 4252 31980
rect 4304 31968 4310 32020
rect 5166 31968 5172 32020
rect 5224 32008 5230 32020
rect 5353 32011 5411 32017
rect 5353 32008 5365 32011
rect 5224 31980 5365 32008
rect 5224 31968 5230 31980
rect 5353 31977 5365 31980
rect 5399 31977 5411 32011
rect 6822 32008 6828 32020
rect 6783 31980 6828 32008
rect 5353 31971 5411 31977
rect 6822 31968 6828 31980
rect 6880 31968 6886 32020
rect 6914 31968 6920 32020
rect 6972 32008 6978 32020
rect 8021 32011 8079 32017
rect 8021 32008 8033 32011
rect 6972 31980 8033 32008
rect 6972 31968 6978 31980
rect 8021 31977 8033 31980
rect 8067 31977 8079 32011
rect 9858 32008 9864 32020
rect 9819 31980 9864 32008
rect 8021 31971 8079 31977
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 12434 32008 12440 32020
rect 12395 31980 12440 32008
rect 12434 31968 12440 31980
rect 12492 31968 12498 32020
rect 1578 31872 1584 31884
rect 1539 31844 1584 31872
rect 1578 31832 1584 31844
rect 1636 31832 1642 31884
rect 2685 31875 2743 31881
rect 2685 31841 2697 31875
rect 2731 31841 2743 31875
rect 2685 31835 2743 31841
rect 4065 31875 4123 31881
rect 4065 31841 4077 31875
rect 4111 31872 4123 31875
rect 4154 31872 4160 31884
rect 4111 31844 4160 31872
rect 4111 31841 4123 31844
rect 4065 31835 4123 31841
rect 2700 31804 2728 31835
rect 4154 31832 4160 31844
rect 4212 31832 4218 31884
rect 5166 31872 5172 31884
rect 5127 31844 5172 31872
rect 5166 31832 5172 31844
rect 5224 31832 5230 31884
rect 6641 31875 6699 31881
rect 6641 31841 6653 31875
rect 6687 31841 6699 31875
rect 7834 31872 7840 31884
rect 7795 31844 7840 31872
rect 6641 31835 6699 31841
rect 6656 31804 6684 31835
rect 7834 31832 7840 31844
rect 7892 31832 7898 31884
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31872 9735 31875
rect 10318 31872 10324 31884
rect 9723 31844 10324 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 12253 31875 12311 31881
rect 12253 31841 12265 31875
rect 12299 31872 12311 31875
rect 13354 31872 13360 31884
rect 12299 31844 12388 31872
rect 13315 31844 13360 31872
rect 12299 31841 12311 31844
rect 12253 31835 12311 31841
rect 2700 31776 2820 31804
rect 6656 31776 6868 31804
rect 2792 31736 2820 31776
rect 3234 31736 3240 31748
rect 2792 31708 3240 31736
rect 3234 31696 3240 31708
rect 3292 31696 3298 31748
rect 6840 31736 6868 31776
rect 7374 31736 7380 31748
rect 6840 31708 7380 31736
rect 7374 31696 7380 31708
rect 7432 31696 7438 31748
rect 12360 31736 12388 31844
rect 13354 31832 13360 31844
rect 13412 31832 13418 31884
rect 12986 31736 12992 31748
rect 12360 31708 12992 31736
rect 12986 31696 12992 31708
rect 13044 31696 13050 31748
rect 13538 31668 13544 31680
rect 13499 31640 13544 31668
rect 13538 31628 13544 31640
rect 13596 31628 13602 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 2866 31464 2872 31476
rect 2827 31436 2872 31464
rect 2866 31424 2872 31436
rect 2924 31424 2930 31476
rect 7009 31467 7067 31473
rect 7009 31433 7021 31467
rect 7055 31464 7067 31467
rect 7098 31464 7104 31476
rect 7055 31436 7104 31464
rect 7055 31433 7067 31436
rect 7009 31427 7067 31433
rect 7098 31424 7104 31436
rect 7156 31424 7162 31476
rect 8294 31424 8300 31476
rect 8352 31464 8358 31476
rect 8849 31467 8907 31473
rect 8849 31464 8861 31467
rect 8352 31436 8861 31464
rect 8352 31424 8358 31436
rect 8849 31433 8861 31436
rect 8895 31433 8907 31467
rect 9674 31464 9680 31476
rect 9635 31436 9680 31464
rect 8849 31427 8907 31433
rect 9674 31424 9680 31436
rect 9732 31424 9738 31476
rect 13354 31464 13360 31476
rect 13315 31436 13360 31464
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 2774 31356 2780 31408
rect 2832 31396 2838 31408
rect 3973 31399 4031 31405
rect 3973 31396 3985 31399
rect 2832 31368 3985 31396
rect 2832 31356 2838 31368
rect 3973 31365 3985 31368
rect 4019 31365 4031 31399
rect 3973 31359 4031 31365
rect 5534 31356 5540 31408
rect 5592 31396 5598 31408
rect 5813 31399 5871 31405
rect 5813 31396 5825 31399
rect 5592 31368 5825 31396
rect 5592 31356 5598 31368
rect 5813 31365 5825 31368
rect 5859 31365 5871 31399
rect 5813 31359 5871 31365
rect 12526 31356 12532 31408
rect 12584 31396 12590 31408
rect 12621 31399 12679 31405
rect 12621 31396 12633 31399
rect 12584 31368 12633 31396
rect 12584 31356 12590 31368
rect 12621 31365 12633 31368
rect 12667 31365 12679 31399
rect 12621 31359 12679 31365
rect 2685 31263 2743 31269
rect 2685 31260 2697 31263
rect 2516 31232 2697 31260
rect 2516 31136 2544 31232
rect 2685 31229 2697 31232
rect 2731 31229 2743 31263
rect 3789 31263 3847 31269
rect 3789 31260 3801 31263
rect 2685 31223 2743 31229
rect 3620 31232 3801 31260
rect 1578 31124 1584 31136
rect 1539 31096 1584 31124
rect 1578 31084 1584 31096
rect 1636 31084 1642 31136
rect 2498 31124 2504 31136
rect 2459 31096 2504 31124
rect 2498 31084 2504 31096
rect 2556 31084 2562 31136
rect 3234 31124 3240 31136
rect 3195 31096 3240 31124
rect 3234 31084 3240 31096
rect 3292 31084 3298 31136
rect 3326 31084 3332 31136
rect 3384 31124 3390 31136
rect 3620 31133 3648 31232
rect 3789 31229 3801 31232
rect 3835 31229 3847 31263
rect 3789 31223 3847 31229
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31260 5687 31263
rect 6641 31263 6699 31269
rect 5675 31232 6224 31260
rect 5675 31229 5687 31232
rect 5629 31223 5687 31229
rect 6196 31136 6224 31232
rect 6641 31229 6653 31263
rect 6687 31260 6699 31263
rect 6822 31260 6828 31272
rect 6687 31232 6828 31260
rect 6687 31229 6699 31232
rect 6641 31223 6699 31229
rect 6822 31220 6828 31232
rect 6880 31220 6886 31272
rect 8665 31263 8723 31269
rect 8665 31229 8677 31263
rect 8711 31260 8723 31263
rect 8711 31232 9352 31260
rect 8711 31229 8723 31232
rect 8665 31223 8723 31229
rect 9324 31136 9352 31232
rect 9674 31220 9680 31272
rect 9732 31260 9738 31272
rect 9769 31263 9827 31269
rect 9769 31260 9781 31263
rect 9732 31232 9781 31260
rect 9732 31220 9738 31232
rect 9769 31229 9781 31232
rect 9815 31229 9827 31263
rect 9769 31223 9827 31229
rect 12253 31263 12311 31269
rect 12253 31229 12265 31263
rect 12299 31260 12311 31263
rect 12437 31263 12495 31269
rect 12437 31260 12449 31263
rect 12299 31232 12449 31260
rect 12299 31229 12311 31232
rect 12253 31223 12311 31229
rect 12437 31229 12449 31232
rect 12483 31260 12495 31263
rect 14182 31260 14188 31272
rect 12483 31232 14188 31260
rect 12483 31229 12495 31232
rect 12437 31223 12495 31229
rect 14182 31220 14188 31232
rect 14240 31220 14246 31272
rect 3605 31127 3663 31133
rect 3605 31124 3617 31127
rect 3384 31096 3617 31124
rect 3384 31084 3390 31096
rect 3605 31093 3617 31096
rect 3651 31093 3663 31127
rect 3605 31087 3663 31093
rect 4154 31084 4160 31136
rect 4212 31124 4218 31136
rect 4341 31127 4399 31133
rect 4341 31124 4353 31127
rect 4212 31096 4353 31124
rect 4212 31084 4218 31096
rect 4341 31093 4353 31096
rect 4387 31093 4399 31127
rect 4341 31087 4399 31093
rect 4982 31084 4988 31136
rect 5040 31124 5046 31136
rect 5166 31124 5172 31136
rect 5040 31096 5172 31124
rect 5040 31084 5046 31096
rect 5166 31084 5172 31096
rect 5224 31084 5230 31136
rect 6178 31124 6184 31136
rect 6139 31096 6184 31124
rect 6178 31084 6184 31096
rect 6236 31084 6242 31136
rect 7374 31124 7380 31136
rect 7335 31096 7380 31124
rect 7374 31084 7380 31096
rect 7432 31084 7438 31136
rect 7834 31124 7840 31136
rect 7795 31096 7840 31124
rect 7834 31084 7840 31096
rect 7892 31084 7898 31136
rect 9306 31124 9312 31136
rect 9267 31096 9312 31124
rect 9306 31084 9312 31096
rect 9364 31084 9370 31136
rect 9858 31084 9864 31136
rect 9916 31124 9922 31136
rect 9953 31127 10011 31133
rect 9953 31124 9965 31127
rect 9916 31096 9965 31124
rect 9916 31084 9922 31096
rect 9953 31093 9965 31096
rect 9999 31093 10011 31127
rect 9953 31087 10011 31093
rect 10318 31084 10324 31136
rect 10376 31124 10382 31136
rect 10413 31127 10471 31133
rect 10413 31124 10425 31127
rect 10376 31096 10425 31124
rect 10376 31084 10382 31096
rect 10413 31093 10425 31096
rect 10459 31124 10471 31127
rect 10686 31124 10692 31136
rect 10459 31096 10692 31124
rect 10459 31093 10471 31096
rect 10413 31087 10471 31093
rect 10686 31084 10692 31096
rect 10744 31084 10750 31136
rect 12986 31124 12992 31136
rect 12947 31096 12992 31124
rect 12986 31084 12992 31096
rect 13044 31084 13050 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 9950 30920 9956 30932
rect 9911 30892 9956 30920
rect 9950 30880 9956 30892
rect 10008 30880 10014 30932
rect 11054 30920 11060 30932
rect 11015 30892 11060 30920
rect 11054 30880 11060 30892
rect 11112 30880 11118 30932
rect 4338 30784 4344 30796
rect 4299 30756 4344 30784
rect 4338 30744 4344 30756
rect 4396 30744 4402 30796
rect 9769 30787 9827 30793
rect 9769 30753 9781 30787
rect 9815 30784 9827 30787
rect 10410 30784 10416 30796
rect 9815 30756 10416 30784
rect 9815 30753 9827 30756
rect 9769 30747 9827 30753
rect 10410 30744 10416 30756
rect 10468 30744 10474 30796
rect 10873 30787 10931 30793
rect 10873 30753 10885 30787
rect 10919 30784 10931 30787
rect 11422 30784 11428 30796
rect 10919 30756 11428 30784
rect 10919 30753 10931 30756
rect 10873 30747 10931 30753
rect 11422 30744 11428 30756
rect 11480 30744 11486 30796
rect 4062 30540 4068 30592
rect 4120 30580 4126 30592
rect 4525 30583 4583 30589
rect 4525 30580 4537 30583
rect 4120 30552 4537 30580
rect 4120 30540 4126 30552
rect 4525 30549 4537 30552
rect 4571 30549 4583 30583
rect 4525 30543 4583 30549
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 4338 30376 4344 30388
rect 4299 30348 4344 30376
rect 4338 30336 4344 30348
rect 4396 30336 4402 30388
rect 9677 30311 9735 30317
rect 9677 30277 9689 30311
rect 9723 30308 9735 30311
rect 10042 30308 10048 30320
rect 9723 30280 10048 30308
rect 9723 30277 9735 30280
rect 9677 30271 9735 30277
rect 9784 30181 9812 30280
rect 10042 30268 10048 30280
rect 10100 30268 10106 30320
rect 10781 30311 10839 30317
rect 10781 30277 10793 30311
rect 10827 30308 10839 30311
rect 10870 30308 10876 30320
rect 10827 30280 10876 30308
rect 10827 30277 10839 30280
rect 10781 30271 10839 30277
rect 10870 30268 10876 30280
rect 10928 30268 10934 30320
rect 10888 30181 10916 30268
rect 9769 30175 9827 30181
rect 9769 30141 9781 30175
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 10873 30175 10931 30181
rect 10873 30141 10885 30175
rect 10919 30141 10931 30175
rect 10873 30135 10931 30141
rect 9950 30036 9956 30048
rect 9911 30008 9956 30036
rect 9950 29996 9956 30008
rect 10008 29996 10014 30048
rect 10410 30036 10416 30048
rect 10371 30008 10416 30036
rect 10410 29996 10416 30008
rect 10468 29996 10474 30048
rect 11054 30036 11060 30048
rect 11015 30008 11060 30036
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 11422 30036 11428 30048
rect 11383 30008 11428 30036
rect 11422 29996 11428 30008
rect 11480 29996 11486 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 10226 29696 10232 29708
rect 10187 29668 10232 29696
rect 10226 29656 10232 29668
rect 10284 29656 10290 29708
rect 9674 29452 9680 29504
rect 9732 29492 9738 29504
rect 10413 29495 10471 29501
rect 10413 29492 10425 29495
rect 9732 29464 10425 29492
rect 9732 29452 9738 29464
rect 10413 29461 10425 29464
rect 10459 29461 10471 29495
rect 10413 29455 10471 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 10137 29291 10195 29297
rect 10137 29257 10149 29291
rect 10183 29288 10195 29291
rect 10226 29288 10232 29300
rect 10183 29260 10232 29288
rect 10183 29257 10195 29260
rect 10137 29251 10195 29257
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 9766 29180 9772 29232
rect 9824 29220 9830 29232
rect 10413 29223 10471 29229
rect 10413 29220 10425 29223
rect 9824 29192 10425 29220
rect 9824 29180 9830 29192
rect 10413 29189 10425 29192
rect 10459 29189 10471 29223
rect 10413 29183 10471 29189
rect 10226 29084 10232 29096
rect 10187 29056 10232 29084
rect 10226 29044 10232 29056
rect 10284 29084 10290 29096
rect 10781 29087 10839 29093
rect 10781 29084 10793 29087
rect 10284 29056 10793 29084
rect 10284 29044 10290 29056
rect 10781 29053 10793 29056
rect 10827 29053 10839 29087
rect 10781 29047 10839 29053
rect 4154 28908 4160 28960
rect 4212 28948 4218 28960
rect 4614 28948 4620 28960
rect 4212 28920 4620 28948
rect 4212 28908 4218 28920
rect 4614 28908 4620 28920
rect 4672 28908 4678 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1486 27072 1492 27124
rect 1544 27112 1550 27124
rect 1581 27115 1639 27121
rect 1581 27112 1593 27115
rect 1544 27084 1593 27112
rect 1544 27072 1550 27084
rect 1581 27081 1593 27084
rect 1627 27081 1639 27115
rect 1581 27075 1639 27081
rect 10318 27004 10324 27056
rect 10376 27044 10382 27056
rect 10594 27044 10600 27056
rect 10376 27016 10600 27044
rect 10376 27004 10382 27016
rect 10594 27004 10600 27016
rect 10652 27004 10658 27056
rect 1397 26911 1455 26917
rect 1397 26877 1409 26911
rect 1443 26908 1455 26911
rect 1443 26880 1992 26908
rect 1443 26877 1455 26880
rect 1397 26871 1455 26877
rect 1964 26781 1992 26880
rect 7466 26868 7472 26920
rect 7524 26908 7530 26920
rect 8018 26908 8024 26920
rect 7524 26880 8024 26908
rect 7524 26868 7530 26880
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 8386 26868 8392 26920
rect 8444 26908 8450 26920
rect 9398 26908 9404 26920
rect 8444 26880 9404 26908
rect 8444 26868 8450 26880
rect 9398 26868 9404 26880
rect 9456 26868 9462 26920
rect 10134 26868 10140 26920
rect 10192 26908 10198 26920
rect 10594 26908 10600 26920
rect 10192 26880 10600 26908
rect 10192 26868 10198 26880
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 1949 26775 2007 26781
rect 1949 26741 1961 26775
rect 1995 26772 2007 26775
rect 2682 26772 2688 26784
rect 1995 26744 2688 26772
rect 1995 26741 2007 26744
rect 1949 26735 2007 26741
rect 2682 26732 2688 26744
rect 2740 26732 2746 26784
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26772 7159 26775
rect 7190 26772 7196 26784
rect 7147 26744 7196 26772
rect 7147 26741 7159 26744
rect 7101 26735 7159 26741
rect 7190 26732 7196 26744
rect 7248 26732 7254 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7285 26571 7343 26577
rect 7285 26568 7297 26571
rect 6972 26540 7297 26568
rect 6972 26528 6978 26540
rect 7285 26537 7297 26540
rect 7331 26568 7343 26571
rect 7926 26568 7932 26580
rect 7331 26540 7932 26568
rect 7331 26537 7343 26540
rect 7285 26531 7343 26537
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 7190 26432 7196 26444
rect 7151 26404 7196 26432
rect 7190 26392 7196 26404
rect 7248 26392 7254 26444
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26364 7527 26367
rect 7558 26364 7564 26376
rect 7515 26336 7564 26364
rect 7515 26333 7527 26336
rect 7469 26327 7527 26333
rect 7558 26324 7564 26336
rect 7616 26324 7622 26376
rect 2406 26256 2412 26308
rect 2464 26296 2470 26308
rect 2590 26296 2596 26308
rect 2464 26268 2596 26296
rect 2464 26256 2470 26268
rect 2590 26256 2596 26268
rect 2648 26256 2654 26308
rect 5077 26299 5135 26305
rect 5077 26265 5089 26299
rect 5123 26296 5135 26299
rect 5350 26296 5356 26308
rect 5123 26268 5356 26296
rect 5123 26265 5135 26268
rect 5077 26259 5135 26265
rect 5350 26256 5356 26268
rect 5408 26296 5414 26308
rect 6825 26299 6883 26305
rect 6825 26296 6837 26299
rect 5408 26268 6837 26296
rect 5408 26256 5414 26268
rect 6825 26265 6837 26268
rect 6871 26265 6883 26299
rect 6825 26259 6883 26265
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 6273 26027 6331 26033
rect 6273 25993 6285 26027
rect 6319 26024 6331 26027
rect 6914 26024 6920 26036
rect 6319 25996 6920 26024
rect 6319 25993 6331 25996
rect 6273 25987 6331 25993
rect 6914 25984 6920 25996
rect 6972 25984 6978 26036
rect 6825 25959 6883 25965
rect 6825 25956 6837 25959
rect 5460 25928 6837 25956
rect 5074 25848 5080 25900
rect 5132 25888 5138 25900
rect 5460 25897 5488 25928
rect 6825 25925 6837 25928
rect 6871 25925 6883 25959
rect 6825 25919 6883 25925
rect 5445 25891 5503 25897
rect 5445 25888 5457 25891
rect 5132 25860 5457 25888
rect 5132 25848 5138 25860
rect 5445 25857 5457 25860
rect 5491 25857 5503 25891
rect 5445 25851 5503 25857
rect 5537 25891 5595 25897
rect 5537 25857 5549 25891
rect 5583 25857 5595 25891
rect 7282 25888 7288 25900
rect 7243 25860 7288 25888
rect 5537 25851 5595 25857
rect 5350 25820 5356 25832
rect 5311 25792 5356 25820
rect 5350 25780 5356 25792
rect 5408 25780 5414 25832
rect 5552 25820 5580 25851
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7558 25888 7564 25900
rect 7515 25860 7564 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7558 25848 7564 25860
rect 7616 25848 7622 25900
rect 5460 25792 5580 25820
rect 4801 25755 4859 25761
rect 4801 25721 4813 25755
rect 4847 25752 4859 25755
rect 5258 25752 5264 25764
rect 4847 25724 5264 25752
rect 4847 25721 4859 25724
rect 4801 25715 4859 25721
rect 5258 25712 5264 25724
rect 5316 25752 5322 25764
rect 5460 25752 5488 25792
rect 5316 25724 5488 25752
rect 5316 25712 5322 25724
rect 4890 25644 4896 25696
rect 4948 25684 4954 25696
rect 4985 25687 5043 25693
rect 4985 25684 4997 25687
rect 4948 25656 4997 25684
rect 4948 25644 4954 25656
rect 4985 25653 4997 25656
rect 5031 25653 5043 25687
rect 4985 25647 5043 25653
rect 6641 25687 6699 25693
rect 6641 25653 6653 25687
rect 6687 25684 6699 25687
rect 7193 25687 7251 25693
rect 7193 25684 7205 25687
rect 6687 25656 7205 25684
rect 6687 25653 6699 25656
rect 6641 25647 6699 25653
rect 7193 25653 7205 25656
rect 7239 25684 7251 25687
rect 7374 25684 7380 25696
rect 7239 25656 7380 25684
rect 7239 25653 7251 25656
rect 7193 25647 7251 25653
rect 7374 25644 7380 25656
rect 7432 25644 7438 25696
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 7837 25687 7895 25693
rect 7837 25684 7849 25687
rect 7616 25656 7849 25684
rect 7616 25644 7622 25656
rect 7837 25653 7849 25656
rect 7883 25653 7895 25687
rect 7837 25647 7895 25653
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 3145 25483 3203 25489
rect 3145 25449 3157 25483
rect 3191 25480 3203 25483
rect 3418 25480 3424 25492
rect 3191 25452 3424 25480
rect 3191 25449 3203 25452
rect 3145 25443 3203 25449
rect 3418 25440 3424 25452
rect 3476 25480 3482 25492
rect 4890 25480 4896 25492
rect 3476 25452 4896 25480
rect 3476 25440 3482 25452
rect 4890 25440 4896 25452
rect 4948 25440 4954 25492
rect 5074 25480 5080 25492
rect 5035 25452 5080 25480
rect 5074 25440 5080 25452
rect 5132 25440 5138 25492
rect 7190 25480 7196 25492
rect 7151 25452 7196 25480
rect 7190 25440 7196 25452
rect 7248 25440 7254 25492
rect 12250 25480 12256 25492
rect 12211 25452 12256 25480
rect 12250 25440 12256 25452
rect 12308 25440 12314 25492
rect 6917 25415 6975 25421
rect 6917 25381 6929 25415
rect 6963 25412 6975 25415
rect 7282 25412 7288 25424
rect 6963 25384 7288 25412
rect 6963 25381 6975 25384
rect 6917 25375 6975 25381
rect 7282 25372 7288 25384
rect 7340 25372 7346 25424
rect 12066 25344 12072 25356
rect 12027 25316 12072 25344
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 7558 25140 7564 25152
rect 7519 25112 7564 25140
rect 7558 25100 7564 25112
rect 7616 25100 7622 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 2866 24760 2872 24812
rect 2924 24800 2930 24812
rect 3605 24803 3663 24809
rect 3605 24800 3617 24803
rect 2924 24772 3617 24800
rect 2924 24760 2930 24772
rect 3605 24769 3617 24772
rect 3651 24769 3663 24803
rect 3605 24763 3663 24769
rect 3418 24732 3424 24744
rect 3379 24704 3424 24732
rect 3418 24692 3424 24704
rect 3476 24692 3482 24744
rect 2774 24624 2780 24676
rect 2832 24664 2838 24676
rect 2832 24636 3096 24664
rect 2832 24624 2838 24636
rect 2866 24596 2872 24608
rect 2827 24568 2872 24596
rect 2866 24556 2872 24568
rect 2924 24556 2930 24608
rect 3068 24605 3096 24636
rect 3053 24599 3111 24605
rect 3053 24565 3065 24599
rect 3099 24565 3111 24599
rect 3510 24596 3516 24608
rect 3471 24568 3516 24596
rect 3053 24559 3111 24565
rect 3510 24556 3516 24568
rect 3568 24556 3574 24608
rect 11054 24556 11060 24608
rect 11112 24596 11118 24608
rect 12066 24596 12072 24608
rect 11112 24568 12072 24596
rect 11112 24556 11118 24568
rect 12066 24556 12072 24568
rect 12124 24556 12130 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 3145 24055 3203 24061
rect 3145 24021 3157 24055
rect 3191 24052 3203 24055
rect 3510 24052 3516 24064
rect 3191 24024 3516 24052
rect 3191 24021 3203 24024
rect 3145 24015 3203 24021
rect 3510 24012 3516 24024
rect 3568 24052 3574 24064
rect 3970 24052 3976 24064
rect 3568 24024 3976 24052
rect 3568 24012 3574 24024
rect 3970 24012 3976 24024
rect 4028 24012 4034 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 11330 22108 11336 22160
rect 11388 22148 11394 22160
rect 12158 22148 12164 22160
rect 11388 22120 12164 22148
rect 11388 22108 11394 22120
rect 12158 22108 12164 22120
rect 12216 22108 12222 22160
rect 4522 21876 4528 21888
rect 4483 21848 4528 21876
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 4433 21675 4491 21681
rect 4433 21672 4445 21675
rect 4028 21644 4445 21672
rect 4028 21632 4034 21644
rect 4433 21641 4445 21644
rect 4479 21641 4491 21675
rect 4433 21635 4491 21641
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21536 4399 21539
rect 5077 21539 5135 21545
rect 5077 21536 5089 21539
rect 4387 21508 5089 21536
rect 4387 21505 4399 21508
rect 4341 21499 4399 21505
rect 5077 21505 5089 21508
rect 5123 21536 5135 21539
rect 5258 21536 5264 21548
rect 5123 21508 5264 21536
rect 5123 21505 5135 21508
rect 5077 21499 5135 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 4522 21428 4528 21480
rect 4580 21468 4586 21480
rect 4801 21471 4859 21477
rect 4801 21468 4813 21471
rect 4580 21440 4813 21468
rect 4580 21428 4586 21440
rect 4801 21437 4813 21440
rect 4847 21437 4859 21471
rect 4801 21431 4859 21437
rect 4890 21292 4896 21344
rect 4948 21332 4954 21344
rect 4948 21304 4993 21332
rect 4948 21292 4954 21304
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 4522 21088 4528 21140
rect 4580 21128 4586 21140
rect 5997 21131 6055 21137
rect 5997 21128 6009 21131
rect 4580 21100 6009 21128
rect 4580 21088 4586 21100
rect 5997 21097 6009 21100
rect 6043 21097 6055 21131
rect 5997 21091 6055 21097
rect 5534 21020 5540 21072
rect 5592 21060 5598 21072
rect 6086 21060 6092 21072
rect 5592 21032 6092 21060
rect 5592 21020 5598 21032
rect 6086 21020 6092 21032
rect 6144 21060 6150 21072
rect 6365 21063 6423 21069
rect 6365 21060 6377 21063
rect 6144 21032 6377 21060
rect 6144 21020 6150 21032
rect 6365 21029 6377 21032
rect 6411 21029 6423 21063
rect 6365 21023 6423 21029
rect 6457 20995 6515 21001
rect 6457 20961 6469 20995
rect 6503 20992 6515 20995
rect 6730 20992 6736 21004
rect 6503 20964 6736 20992
rect 6503 20961 6515 20964
rect 6457 20955 6515 20961
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6454 20816 6460 20868
rect 6512 20856 6518 20868
rect 6564 20856 6592 20887
rect 6512 20828 6592 20856
rect 6512 20816 6518 20828
rect 4525 20791 4583 20797
rect 4525 20757 4537 20791
rect 4571 20788 4583 20791
rect 4890 20788 4896 20800
rect 4571 20760 4896 20788
rect 4571 20757 4583 20760
rect 4525 20751 4583 20757
rect 4890 20748 4896 20760
rect 4948 20788 4954 20800
rect 5442 20788 5448 20800
rect 4948 20760 5448 20788
rect 4948 20748 4954 20760
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 6086 20584 6092 20596
rect 6047 20556 6092 20584
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 9674 20516 9680 20528
rect 9635 20488 9680 20516
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 6454 20448 6460 20460
rect 6415 20420 6460 20448
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 3007 20352 3065 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 3053 20349 3065 20352
rect 3099 20380 3111 20383
rect 5721 20383 5779 20389
rect 3099 20352 4016 20380
rect 3099 20349 3111 20352
rect 3053 20343 3111 20349
rect 3988 20324 4016 20352
rect 5721 20349 5733 20383
rect 5767 20380 5779 20383
rect 6730 20380 6736 20392
rect 5767 20352 6736 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 6730 20340 6736 20352
rect 6788 20340 6794 20392
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 3326 20321 3332 20324
rect 3320 20312 3332 20321
rect 3287 20284 3332 20312
rect 3320 20275 3332 20284
rect 3326 20272 3332 20275
rect 3384 20272 3390 20324
rect 3970 20272 3976 20324
rect 4028 20272 4034 20324
rect 4430 20244 4436 20256
rect 4391 20216 4436 20244
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 8202 20244 8208 20256
rect 8115 20216 8208 20244
rect 8202 20204 8208 20216
rect 8260 20244 8266 20256
rect 8312 20244 8340 20343
rect 8570 20321 8576 20324
rect 8564 20312 8576 20321
rect 8531 20284 8576 20312
rect 8564 20275 8576 20284
rect 8570 20272 8576 20275
rect 8628 20272 8634 20324
rect 9674 20244 9680 20256
rect 8260 20216 9680 20244
rect 8260 20204 8266 20216
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3326 20040 3332 20052
rect 3191 20012 3332 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 5534 20040 5540 20052
rect 5495 20012 5540 20040
rect 5534 20000 5540 20012
rect 5592 20000 5598 20052
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 7101 20043 7159 20049
rect 7101 20040 7113 20043
rect 6788 20012 7113 20040
rect 6788 20000 6794 20012
rect 7101 20009 7113 20012
rect 7147 20009 7159 20043
rect 7101 20003 7159 20009
rect 7374 20000 7380 20052
rect 7432 20040 7438 20052
rect 7561 20043 7619 20049
rect 7561 20040 7573 20043
rect 7432 20012 7573 20040
rect 7432 20000 7438 20012
rect 7561 20009 7573 20012
rect 7607 20009 7619 20043
rect 7561 20003 7619 20009
rect 4430 19932 4436 19984
rect 4488 19972 4494 19984
rect 4614 19972 4620 19984
rect 4488 19944 4620 19972
rect 4488 19932 4494 19944
rect 4614 19932 4620 19944
rect 4672 19932 4678 19984
rect 5905 19975 5963 19981
rect 5905 19941 5917 19975
rect 5951 19972 5963 19975
rect 6086 19972 6092 19984
rect 5951 19944 6092 19972
rect 5951 19941 5963 19944
rect 5905 19935 5963 19941
rect 6086 19932 6092 19944
rect 6144 19932 6150 19984
rect 7469 19975 7527 19981
rect 7469 19941 7481 19975
rect 7515 19972 7527 19975
rect 7742 19972 7748 19984
rect 7515 19944 7748 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 7742 19932 7748 19944
rect 7800 19932 7806 19984
rect 9944 19975 10002 19981
rect 9944 19941 9956 19975
rect 9990 19972 10002 19975
rect 10042 19972 10048 19984
rect 9990 19944 10048 19972
rect 9990 19941 10002 19944
rect 9944 19935 10002 19941
rect 10042 19932 10048 19944
rect 10100 19932 10106 19984
rect 6917 19907 6975 19913
rect 6917 19873 6929 19907
rect 6963 19904 6975 19907
rect 7098 19904 7104 19916
rect 6963 19876 7104 19904
rect 6963 19873 6975 19876
rect 6917 19867 6975 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 5994 19836 6000 19848
rect 5955 19808 6000 19836
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19836 6239 19839
rect 6822 19836 6828 19848
rect 6227 19808 6828 19836
rect 6227 19805 6239 19808
rect 6181 19799 6239 19805
rect 5534 19728 5540 19780
rect 5592 19768 5598 19780
rect 6196 19768 6224 19799
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 9674 19836 9680 19848
rect 7791 19808 8432 19836
rect 9635 19808 9680 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 5592 19740 6224 19768
rect 5592 19728 5598 19740
rect 8404 19709 8432 19808
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 8389 19703 8447 19709
rect 8389 19669 8401 19703
rect 8435 19700 8447 19703
rect 8570 19700 8576 19712
rect 8435 19672 8576 19700
rect 8435 19669 8447 19672
rect 8389 19663 8447 19669
rect 8570 19660 8576 19672
rect 8628 19700 8634 19712
rect 11057 19703 11115 19709
rect 11057 19700 11069 19703
rect 8628 19672 11069 19700
rect 8628 19660 8634 19672
rect 11057 19669 11069 19672
rect 11103 19669 11115 19703
rect 11057 19663 11115 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 3970 19496 3976 19508
rect 3927 19468 3976 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 7374 19456 7380 19508
rect 7432 19496 7438 19508
rect 7558 19496 7564 19508
rect 7432 19468 7564 19496
rect 7432 19456 7438 19468
rect 7558 19456 7564 19468
rect 7616 19496 7622 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7616 19468 7849 19496
rect 7616 19456 7622 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 7837 19459 7895 19465
rect 8297 19499 8355 19505
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 8570 19496 8576 19508
rect 8343 19468 8576 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 3988 19369 4016 19456
rect 5994 19388 6000 19440
rect 6052 19428 6058 19440
rect 6825 19431 6883 19437
rect 6825 19428 6837 19431
rect 6052 19400 6837 19428
rect 6052 19388 6058 19400
rect 6825 19397 6837 19400
rect 6871 19397 6883 19431
rect 6825 19391 6883 19397
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19329 4031 19363
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 3973 19323 4031 19329
rect 6748 19332 7481 19360
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 4240 19295 4298 19301
rect 4240 19292 4252 19295
rect 3559 19264 4252 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 4240 19261 4252 19264
rect 4286 19292 4298 19295
rect 5534 19292 5540 19304
rect 4286 19264 5540 19292
rect 4286 19261 4298 19264
rect 4240 19255 4298 19261
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6748 19292 6776 19332
rect 7469 19329 7481 19332
rect 7515 19360 7527 19363
rect 8312 19360 8340 19459
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 7515 19332 8340 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 10502 19360 10508 19372
rect 10376 19332 10508 19360
rect 10376 19320 10382 19332
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 6380 19264 6776 19292
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5316 19128 5365 19156
rect 5316 19116 5322 19128
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 5353 19119 5411 19125
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 5776 19128 6193 19156
rect 5776 19116 5782 19128
rect 6181 19125 6193 19128
rect 6227 19156 6239 19159
rect 6380 19156 6408 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 6546 19224 6552 19236
rect 6507 19196 6552 19224
rect 6546 19184 6552 19196
rect 6604 19224 6610 19236
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 6604 19196 7297 19224
rect 6604 19184 6610 19196
rect 7285 19193 7297 19196
rect 7331 19224 7343 19227
rect 8662 19224 8668 19236
rect 7331 19196 8668 19224
rect 7331 19193 7343 19196
rect 7285 19187 7343 19193
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 9674 19156 9680 19168
rect 6227 19128 6408 19156
rect 9635 19128 9680 19156
rect 6227 19125 6239 19128
rect 6181 19119 6239 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 5534 18952 5540 18964
rect 5495 18924 5540 18952
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 5994 18952 6000 18964
rect 5955 18924 6000 18952
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 6086 18912 6092 18964
rect 6144 18952 6150 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 6144 18924 6285 18952
rect 6144 18912 6150 18924
rect 6273 18921 6285 18924
rect 6319 18952 6331 18955
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 6319 18924 6469 18952
rect 6319 18921 6331 18924
rect 6273 18915 6331 18921
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6822 18952 6828 18964
rect 6457 18915 6515 18921
rect 6656 18924 6828 18952
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 6086 18816 6092 18828
rect 5868 18788 6092 18816
rect 5868 18776 5874 18788
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 5994 18748 6000 18760
rect 5684 18720 6000 18748
rect 5684 18708 5690 18720
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 6656 18748 6684 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7374 18912 7380 18964
rect 7432 18952 7438 18964
rect 7561 18955 7619 18961
rect 7561 18952 7573 18955
rect 7432 18924 7573 18952
rect 7432 18912 7438 18924
rect 7561 18921 7573 18924
rect 7607 18952 7619 18955
rect 7742 18952 7748 18964
rect 7607 18924 7748 18952
rect 7607 18921 7619 18924
rect 7561 18915 7619 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6788 18788 6837 18816
rect 6788 18776 6794 18788
rect 6825 18785 6837 18788
rect 6871 18816 6883 18819
rect 8386 18816 8392 18828
rect 6871 18788 8392 18816
rect 6871 18785 6883 18788
rect 6825 18779 6883 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6656 18720 6929 18748
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 5718 18640 5724 18692
rect 5776 18680 5782 18692
rect 7024 18680 7052 18711
rect 5776 18652 7052 18680
rect 5776 18640 5782 18652
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 6089 18411 6147 18417
rect 6089 18408 6101 18411
rect 5776 18380 6101 18408
rect 5776 18368 5782 18380
rect 6089 18377 6101 18380
rect 6135 18377 6147 18411
rect 6089 18371 6147 18377
rect 5718 18096 5724 18148
rect 5776 18136 5782 18148
rect 6730 18136 6736 18148
rect 5776 18108 6736 18136
rect 5776 18096 5782 18108
rect 6730 18096 6736 18108
rect 6788 18136 6794 18148
rect 7009 18139 7067 18145
rect 7009 18136 7021 18139
rect 6788 18108 7021 18136
rect 6788 18096 6794 18108
rect 7009 18105 7021 18108
rect 7055 18105 7067 18139
rect 7009 18099 7067 18105
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 5684 18040 6469 18068
rect 5684 18028 5690 18040
rect 6457 18037 6469 18040
rect 6503 18068 6515 18071
rect 6822 18068 6828 18080
rect 6503 18040 6828 18068
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 11517 13515 11575 13521
rect 11517 13512 11529 13515
rect 10100 13484 11529 13512
rect 10100 13472 10106 13484
rect 11517 13481 11529 13484
rect 11563 13481 11575 13515
rect 11517 13475 11575 13481
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 10393 13379 10451 13385
rect 10393 13376 10405 13379
rect 9640 13348 10405 13376
rect 9640 13336 9646 13348
rect 10393 13345 10405 13348
rect 10439 13345 10451 13379
rect 10393 13339 10451 13345
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9858 13308 9864 13320
rect 9732 13280 9864 13308
rect 9732 13268 9738 13280
rect 9858 13268 9864 13280
rect 9916 13308 9922 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9916 13280 10149 13308
rect 9916 13268 9922 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10778 12968 10784 12980
rect 10091 12940 10784 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10100 12804 10609 12832
rect 10100 12792 10106 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10468 12736 10517 12764
rect 10468 12724 10474 12736
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 9217 12699 9275 12705
rect 9217 12665 9229 12699
rect 9263 12696 9275 12699
rect 9263 12668 9996 12696
rect 9263 12665 9275 12668
rect 9217 12659 9275 12665
rect 9968 12640 9996 12668
rect 9582 12628 9588 12640
rect 9543 12600 9588 12628
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9858 12628 9864 12640
rect 9819 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10008 12600 10425 12628
rect 10008 12588 10014 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 10042 12424 10048 12436
rect 10003 12396 10048 12424
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6730 12220 6736 12232
rect 6052 12192 6736 12220
rect 6052 12180 6058 12192
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8846 12084 8852 12096
rect 8527 12056 8852 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 10410 12084 10416 12096
rect 10371 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 10410 11880 10416 11892
rect 8435 11852 10416 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7374 11744 7380 11756
rect 7248 11716 7380 11744
rect 7248 11704 7254 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 9030 11744 9036 11756
rect 8343 11716 9036 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 7374 11608 7380 11620
rect 7156 11580 7380 11608
rect 7156 11568 7162 11580
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 7929 11611 7987 11617
rect 7929 11577 7941 11611
rect 7975 11608 7987 11611
rect 8478 11608 8484 11620
rect 7975 11580 8484 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 8478 11568 8484 11580
rect 8536 11608 8542 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8536 11580 8769 11608
rect 8536 11568 8542 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 8846 11540 8852 11552
rect 8807 11512 8852 11540
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 8481 10999 8539 11005
rect 6972 10968 7017 10996
rect 6972 10956 6978 10968
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 8846 10996 8852 11008
rect 8527 10968 8852 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 6822 10792 6828 10804
rect 6783 10764 6828 10792
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 8389 10795 8447 10801
rect 8389 10761 8401 10795
rect 8435 10792 8447 10795
rect 8478 10792 8484 10804
rect 8435 10764 8484 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 6687 10628 7481 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7469 10625 7481 10628
rect 7515 10656 7527 10659
rect 8938 10656 8944 10668
rect 7515 10628 8944 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 6972 10560 7205 10588
rect 6972 10548 6978 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8478 10588 8484 10600
rect 8352 10560 8484 10588
rect 8352 10548 8358 10560
rect 8478 10548 8484 10560
rect 8536 10588 8542 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8536 10560 8769 10588
rect 8536 10548 8542 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 6972 10424 7297 10452
rect 6972 10412 6978 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 8846 10452 8852 10464
rect 8807 10424 8852 10452
rect 7285 10415 7343 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 5537 10251 5595 10257
rect 5537 10217 5549 10251
rect 5583 10248 5595 10251
rect 7101 10251 7159 10257
rect 5583 10220 6224 10248
rect 5583 10217 5595 10220
rect 5537 10211 5595 10217
rect 5902 10180 5908 10192
rect 5863 10152 5908 10180
rect 5902 10140 5908 10152
rect 5960 10140 5966 10192
rect 5994 10140 6000 10192
rect 6052 10180 6058 10192
rect 6196 10180 6224 10220
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 8846 10248 8852 10260
rect 7147 10220 8852 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 6914 10180 6920 10192
rect 6052 10152 6097 10180
rect 6196 10152 6920 10180
rect 6052 10140 6058 10152
rect 6914 10140 6920 10152
rect 6972 10180 6978 10192
rect 7466 10180 7472 10192
rect 6972 10152 7017 10180
rect 7427 10152 7472 10180
rect 6972 10140 6978 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6196 9976 6224 10007
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7064 10016 7573 10044
rect 7064 10004 7070 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 6840 9976 6868 10004
rect 7668 9976 7696 10007
rect 6196 9948 7696 9976
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 8846 9908 8852 9920
rect 8527 9880 8852 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 5902 9704 5908 9716
rect 5863 9676 5908 9704
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7466 9704 7472 9716
rect 7156 9676 7472 9704
rect 7156 9664 7162 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5629 9639 5687 9645
rect 5629 9636 5641 9639
rect 5592 9608 5641 9636
rect 5592 9596 5598 9608
rect 5629 9605 5641 9608
rect 5675 9636 5687 9639
rect 5994 9636 6000 9648
rect 5675 9608 6000 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 6932 9404 7849 9432
rect 6932 9376 6960 9404
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6914 9364 6920 9376
rect 6411 9336 6920 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 7064 9336 7113 9364
rect 7064 9324 7070 9336
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 7101 9327 7159 9333
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 5810 9160 5816 9172
rect 5771 9132 5816 9160
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6052 9132 6285 9160
rect 6052 9120 6058 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 6178 9024 6184 9036
rect 6139 8996 6184 9024
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6914 8956 6920 8968
rect 6503 8928 6920 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 5905 8619 5963 8625
rect 5905 8585 5917 8619
rect 5951 8616 5963 8619
rect 5994 8616 6000 8628
rect 5951 8588 6000 8616
rect 5951 8585 5963 8588
rect 5905 8579 5963 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6178 8412 6184 8424
rect 6139 8384 6184 8412
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6914 8344 6920 8356
rect 6687 8316 6920 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 13354 7936 13360 7948
rect 12492 7908 13360 7936
rect 12492 7896 12498 7908
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 14918 7732 14924 7744
rect 14056 7704 14924 7732
rect 14056 7692 14062 7704
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 15746 7528 15752 7540
rect 13872 7500 15752 7528
rect 13872 7488 13878 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4321 6851 4379 6857
rect 4321 6848 4333 6851
rect 4212 6820 4333 6848
rect 4212 6808 4218 6820
rect 4321 6817 4333 6820
rect 4367 6817 4379 6851
rect 4321 6811 4379 6817
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5316 6616 5457 6644
rect 5316 6604 5322 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10410 6644 10416 6656
rect 10091 6616 10416 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 9950 6440 9956 6452
rect 9911 6412 9956 6440
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4433 6375 4491 6381
rect 4433 6372 4445 6375
rect 4120 6344 4445 6372
rect 4120 6332 4126 6344
rect 4433 6341 4445 6344
rect 4479 6372 4491 6375
rect 5534 6372 5540 6384
rect 4479 6344 5540 6372
rect 4479 6341 4491 6344
rect 4433 6335 4491 6341
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 9907 6276 10609 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10597 6273 10609 6276
rect 10643 6304 10655 6307
rect 10962 6304 10968 6316
rect 10643 6276 10968 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 10226 6168 10232 6180
rect 9539 6140 10232 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 10226 6128 10232 6140
rect 10284 6168 10290 6180
rect 10321 6171 10379 6177
rect 10321 6168 10333 6171
rect 10284 6140 10333 6168
rect 10284 6128 10290 6140
rect 10321 6137 10333 6140
rect 10367 6137 10379 6171
rect 10321 6131 10379 6137
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 10468 6072 10513 6100
rect 10468 6060 10474 6072
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 9950 5769 9956 5772
rect 9944 5760 9956 5769
rect 9911 5732 9956 5760
rect 9944 5723 9956 5732
rect 9950 5720 9956 5723
rect 10008 5720 10014 5772
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 5592 5324 6561 5352
rect 5592 5312 5598 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8846 5352 8852 5364
rect 8251 5324 8852 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 6564 5216 6592 5315
rect 8846 5312 8852 5324
rect 8904 5352 8910 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8904 5324 8953 5352
rect 8904 5312 8910 5324
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 8941 5315 8999 5321
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10410 5352 10416 5364
rect 9907 5324 10416 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6564 5188 6837 5216
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 8956 5216 8984 5315
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 9950 5216 9956 5228
rect 8956 5188 9956 5216
rect 6825 5179 6883 5185
rect 6840 5148 6868 5179
rect 9950 5176 9956 5188
rect 10008 5216 10014 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10008 5188 10425 5216
rect 10008 5176 10014 5188
rect 10413 5185 10425 5188
rect 10459 5216 10471 5219
rect 10778 5216 10784 5228
rect 10459 5188 10784 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10778 5176 10784 5188
rect 10836 5216 10842 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10836 5188 10885 5216
rect 10836 5176 10842 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 6840 5120 9321 5148
rect 9309 5117 9321 5120
rect 9355 5148 9367 5151
rect 9582 5148 9588 5160
rect 9355 5120 9588 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10100 5120 10333 5148
rect 10100 5108 10106 5120
rect 10321 5117 10333 5120
rect 10367 5148 10379 5151
rect 11330 5148 11336 5160
rect 10367 5120 11336 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7070 5083 7128 5089
rect 7070 5080 7082 5083
rect 6972 5052 7082 5080
rect 6972 5040 6978 5052
rect 7070 5049 7082 5052
rect 7116 5049 7128 5083
rect 7070 5043 7128 5049
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 9815 4984 10241 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10229 4981 10241 4984
rect 10275 5012 10287 5015
rect 10318 5012 10324 5024
rect 10275 4984 10324 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 10318 4972 10324 4984
rect 10376 5012 10382 5024
rect 10594 5012 10600 5024
rect 10376 4984 10600 5012
rect 10376 4972 10382 4984
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 9953 4811 10011 4817
rect 6972 4780 7017 4808
rect 6972 4768 6978 4780
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10042 4808 10048 4820
rect 9999 4780 10048 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10226 4808 10232 4820
rect 10187 4780 10232 4808
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 10686 4808 10692 4820
rect 10647 4780 10692 4808
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 10836 4576 10881 4604
rect 10836 4564 10842 4576
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 9950 4264 9956 4276
rect 9911 4236 9956 4264
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10321 4267 10379 4273
rect 10321 4233 10333 4267
rect 10367 4264 10379 4267
rect 10686 4264 10692 4276
rect 10367 4236 10692 4264
rect 10367 4233 10379 4236
rect 10321 4227 10379 4233
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 10336 4196 10364 4227
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 9640 4168 10364 4196
rect 9640 4156 9646 4168
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5442 4128 5448 4140
rect 5040 4100 5448 4128
rect 5040 4088 5046 4100
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6638 4128 6644 4140
rect 5776 4100 6644 4128
rect 5776 4088 5782 4100
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10594 4088 10600 4100
rect 10652 4128 10658 4140
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10652 4100 10977 4128
rect 10652 4088 10658 4100
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3553 4123 3587
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 4065 3547 4123 3553
rect 4080 3516 4108 3547
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5074 3516 5080 3528
rect 4080 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 10962 3516 10968 3528
rect 9824 3488 10968 3516
rect 9824 3476 9830 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4249 3451 4307 3457
rect 4249 3448 4261 3451
rect 4212 3420 4261 3448
rect 4212 3408 4218 3420
rect 4249 3417 4261 3420
rect 4295 3417 4307 3451
rect 4249 3411 4307 3417
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 5353 3383 5411 3389
rect 5353 3380 5365 3383
rect 4580 3352 5365 3380
rect 4580 3340 4586 3352
rect 5353 3349 5365 3352
rect 5399 3349 5411 3383
rect 5353 3343 5411 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4246 3176 4252 3188
rect 4203 3148 4252 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5074 3176 5080 3188
rect 5031 3148 5080 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5224 3148 5733 3176
rect 5224 3136 5230 3148
rect 5721 3145 5733 3148
rect 5767 3176 5779 3179
rect 7282 3176 7288 3188
rect 5767 3148 7288 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3176 7527 3179
rect 7926 3176 7932 3188
rect 7515 3148 7932 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 5261 3111 5319 3117
rect 5261 3108 5273 3111
rect 2648 3080 5273 3108
rect 2648 3068 2654 3080
rect 5261 3077 5273 3080
rect 5307 3077 5319 3111
rect 5261 3071 5319 3077
rect 6086 3040 6092 3052
rect 5092 3012 6092 3040
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3510 2972 3516 2984
rect 2915 2944 3516 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 5092 2981 5120 3012
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 7484 2972 7512 3139
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 6871 2944 7512 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 3988 2904 4016 2935
rect 4614 2904 4620 2916
rect 3988 2876 4620 2904
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2832 2808 3065 2836
rect 2832 2796 2838 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 3053 2799 3111 2805
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7009 2839 7067 2845
rect 7009 2836 7021 2839
rect 6972 2808 7021 2836
rect 6972 2796 6978 2808
rect 7009 2805 7021 2808
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5442 2632 5448 2644
rect 4755 2604 5448 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2332 2496 2360 2592
rect 3510 2564 3516 2576
rect 2884 2536 3516 2564
rect 2884 2505 2912 2536
rect 3510 2524 3516 2536
rect 3568 2524 3574 2576
rect 1719 2468 2360 2496
rect 2869 2499 2927 2505
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4724 2496 4752 2595
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 7098 2632 7104 2644
rect 5859 2604 7104 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 4111 2468 4752 2496
rect 5169 2499 5227 2505
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5828 2496 5856 2595
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7834 2632 7840 2644
rect 7795 2604 7840 2632
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8941 2635 8999 2641
rect 8941 2601 8953 2635
rect 8987 2632 8999 2635
rect 9582 2632 9588 2644
rect 8987 2604 9588 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 5215 2468 5856 2496
rect 7193 2499 7251 2505
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7852 2496 7880 2592
rect 7239 2468 7880 2496
rect 8297 2499 8355 2505
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 8297 2465 8309 2499
rect 8343 2496 8355 2499
rect 8956 2496 8984 2595
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 8343 2468 8984 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 1762 2320 1768 2372
rect 1820 2360 1826 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 1820 2332 5365 2360
rect 1820 2320 1826 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 8481 2363 8539 2369
rect 8481 2360 8493 2363
rect 6604 2332 8493 2360
rect 6604 2320 6610 2332
rect 8481 2329 8493 2332
rect 8527 2329 8539 2363
rect 8481 2323 8539 2329
rect 1854 2292 1860 2304
rect 1815 2264 1860 2292
rect 1854 2252 1860 2264
rect 1912 2252 1918 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 2136 35640 2188 35692
rect 2688 35640 2740 35692
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 204 34892 256 34944
rect 1308 34892 1360 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 4160 34688 4212 34740
rect 5448 34688 5500 34740
rect 1400 34484 1452 34536
rect 2780 34484 2832 34536
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 2780 32512 2832 32564
rect 4528 32512 4580 32564
rect 7472 32555 7524 32564
rect 7472 32521 7481 32555
rect 7481 32521 7515 32555
rect 7515 32521 7524 32555
rect 7472 32512 7524 32521
rect 9312 32555 9364 32564
rect 9312 32521 9321 32555
rect 9321 32521 9355 32555
rect 9355 32521 9364 32555
rect 9312 32512 9364 32521
rect 13084 32555 13136 32564
rect 13084 32521 13093 32555
rect 13093 32521 13127 32555
rect 13127 32521 13136 32555
rect 13084 32512 13136 32521
rect 3148 32351 3200 32360
rect 3148 32317 3157 32351
rect 3157 32317 3191 32351
rect 3191 32317 3200 32351
rect 3148 32308 3200 32317
rect 5080 32308 5132 32360
rect 7472 32308 7524 32360
rect 9312 32308 9364 32360
rect 13084 32308 13136 32360
rect 7012 32215 7064 32224
rect 7012 32181 7021 32215
rect 7021 32181 7055 32215
rect 7055 32181 7064 32215
rect 7012 32172 7064 32181
rect 7656 32172 7708 32224
rect 12624 32215 12676 32224
rect 12624 32181 12633 32215
rect 12633 32181 12667 32215
rect 12667 32181 12676 32215
rect 12624 32172 12676 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 1400 31968 1452 32020
rect 2872 32011 2924 32020
rect 2872 31977 2881 32011
rect 2881 31977 2915 32011
rect 2915 31977 2924 32011
rect 2872 31968 2924 31977
rect 4252 32011 4304 32020
rect 4252 31977 4261 32011
rect 4261 31977 4295 32011
rect 4295 31977 4304 32011
rect 4252 31968 4304 31977
rect 5172 31968 5224 32020
rect 6828 32011 6880 32020
rect 6828 31977 6837 32011
rect 6837 31977 6871 32011
rect 6871 31977 6880 32011
rect 6828 31968 6880 31977
rect 6920 31968 6972 32020
rect 9864 32011 9916 32020
rect 9864 31977 9873 32011
rect 9873 31977 9907 32011
rect 9907 31977 9916 32011
rect 9864 31968 9916 31977
rect 12440 32011 12492 32020
rect 12440 31977 12449 32011
rect 12449 31977 12483 32011
rect 12483 31977 12492 32011
rect 12440 31968 12492 31977
rect 1584 31875 1636 31884
rect 1584 31841 1593 31875
rect 1593 31841 1627 31875
rect 1627 31841 1636 31875
rect 1584 31832 1636 31841
rect 4160 31832 4212 31884
rect 5172 31875 5224 31884
rect 5172 31841 5181 31875
rect 5181 31841 5215 31875
rect 5215 31841 5224 31875
rect 5172 31832 5224 31841
rect 7840 31875 7892 31884
rect 7840 31841 7849 31875
rect 7849 31841 7883 31875
rect 7883 31841 7892 31875
rect 7840 31832 7892 31841
rect 10324 31832 10376 31884
rect 13360 31875 13412 31884
rect 3240 31696 3292 31748
rect 7380 31696 7432 31748
rect 13360 31841 13369 31875
rect 13369 31841 13403 31875
rect 13403 31841 13412 31875
rect 13360 31832 13412 31841
rect 12992 31696 13044 31748
rect 13544 31671 13596 31680
rect 13544 31637 13553 31671
rect 13553 31637 13587 31671
rect 13587 31637 13596 31671
rect 13544 31628 13596 31637
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 2872 31467 2924 31476
rect 2872 31433 2881 31467
rect 2881 31433 2915 31467
rect 2915 31433 2924 31467
rect 2872 31424 2924 31433
rect 7104 31424 7156 31476
rect 8300 31424 8352 31476
rect 9680 31467 9732 31476
rect 9680 31433 9689 31467
rect 9689 31433 9723 31467
rect 9723 31433 9732 31467
rect 9680 31424 9732 31433
rect 13360 31467 13412 31476
rect 13360 31433 13369 31467
rect 13369 31433 13403 31467
rect 13403 31433 13412 31467
rect 13360 31424 13412 31433
rect 2780 31356 2832 31408
rect 5540 31356 5592 31408
rect 12532 31356 12584 31408
rect 1584 31127 1636 31136
rect 1584 31093 1593 31127
rect 1593 31093 1627 31127
rect 1627 31093 1636 31127
rect 1584 31084 1636 31093
rect 2504 31127 2556 31136
rect 2504 31093 2513 31127
rect 2513 31093 2547 31127
rect 2547 31093 2556 31127
rect 2504 31084 2556 31093
rect 3240 31127 3292 31136
rect 3240 31093 3249 31127
rect 3249 31093 3283 31127
rect 3283 31093 3292 31127
rect 3240 31084 3292 31093
rect 3332 31084 3384 31136
rect 6828 31263 6880 31272
rect 6828 31229 6837 31263
rect 6837 31229 6871 31263
rect 6871 31229 6880 31263
rect 6828 31220 6880 31229
rect 9680 31220 9732 31272
rect 14188 31220 14240 31272
rect 4160 31084 4212 31136
rect 4988 31084 5040 31136
rect 5172 31127 5224 31136
rect 5172 31093 5181 31127
rect 5181 31093 5215 31127
rect 5215 31093 5224 31127
rect 5172 31084 5224 31093
rect 6184 31127 6236 31136
rect 6184 31093 6193 31127
rect 6193 31093 6227 31127
rect 6227 31093 6236 31127
rect 6184 31084 6236 31093
rect 7380 31127 7432 31136
rect 7380 31093 7389 31127
rect 7389 31093 7423 31127
rect 7423 31093 7432 31127
rect 7380 31084 7432 31093
rect 7840 31127 7892 31136
rect 7840 31093 7849 31127
rect 7849 31093 7883 31127
rect 7883 31093 7892 31127
rect 7840 31084 7892 31093
rect 9312 31127 9364 31136
rect 9312 31093 9321 31127
rect 9321 31093 9355 31127
rect 9355 31093 9364 31127
rect 9312 31084 9364 31093
rect 9864 31084 9916 31136
rect 10324 31084 10376 31136
rect 10692 31084 10744 31136
rect 12992 31127 13044 31136
rect 12992 31093 13001 31127
rect 13001 31093 13035 31127
rect 13035 31093 13044 31127
rect 12992 31084 13044 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 9956 30923 10008 30932
rect 9956 30889 9965 30923
rect 9965 30889 9999 30923
rect 9999 30889 10008 30923
rect 9956 30880 10008 30889
rect 11060 30923 11112 30932
rect 11060 30889 11069 30923
rect 11069 30889 11103 30923
rect 11103 30889 11112 30923
rect 11060 30880 11112 30889
rect 4344 30787 4396 30796
rect 4344 30753 4353 30787
rect 4353 30753 4387 30787
rect 4387 30753 4396 30787
rect 4344 30744 4396 30753
rect 10416 30744 10468 30796
rect 11428 30744 11480 30796
rect 4068 30540 4120 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 4344 30379 4396 30388
rect 4344 30345 4353 30379
rect 4353 30345 4387 30379
rect 4387 30345 4396 30379
rect 4344 30336 4396 30345
rect 10048 30268 10100 30320
rect 10876 30268 10928 30320
rect 9956 30039 10008 30048
rect 9956 30005 9965 30039
rect 9965 30005 9999 30039
rect 9999 30005 10008 30039
rect 9956 29996 10008 30005
rect 10416 30039 10468 30048
rect 10416 30005 10425 30039
rect 10425 30005 10459 30039
rect 10459 30005 10468 30039
rect 10416 29996 10468 30005
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 11428 30039 11480 30048
rect 11428 30005 11437 30039
rect 11437 30005 11471 30039
rect 11471 30005 11480 30039
rect 11428 29996 11480 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 10232 29699 10284 29708
rect 10232 29665 10241 29699
rect 10241 29665 10275 29699
rect 10275 29665 10284 29699
rect 10232 29656 10284 29665
rect 9680 29452 9732 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 10232 29248 10284 29300
rect 9772 29180 9824 29232
rect 10232 29087 10284 29096
rect 10232 29053 10241 29087
rect 10241 29053 10275 29087
rect 10275 29053 10284 29087
rect 10232 29044 10284 29053
rect 4160 28908 4212 28960
rect 4620 28908 4672 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 1492 27072 1544 27124
rect 10324 27004 10376 27056
rect 10600 27004 10652 27056
rect 7472 26868 7524 26920
rect 8024 26868 8076 26920
rect 8392 26868 8444 26920
rect 9404 26868 9456 26920
rect 10140 26868 10192 26920
rect 10600 26868 10652 26920
rect 2688 26732 2740 26784
rect 7196 26732 7248 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 6920 26528 6972 26580
rect 7932 26528 7984 26580
rect 7196 26435 7248 26444
rect 7196 26401 7205 26435
rect 7205 26401 7239 26435
rect 7239 26401 7248 26435
rect 7196 26392 7248 26401
rect 7564 26324 7616 26376
rect 2412 26256 2464 26308
rect 2596 26256 2648 26308
rect 5356 26256 5408 26308
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 6920 25984 6972 26036
rect 5080 25848 5132 25900
rect 7288 25891 7340 25900
rect 5356 25823 5408 25832
rect 5356 25789 5365 25823
rect 5365 25789 5399 25823
rect 5399 25789 5408 25823
rect 5356 25780 5408 25789
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 7564 25848 7616 25900
rect 5264 25712 5316 25764
rect 4896 25644 4948 25696
rect 7380 25644 7432 25696
rect 7564 25644 7616 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 3424 25440 3476 25492
rect 4896 25440 4948 25492
rect 5080 25483 5132 25492
rect 5080 25449 5089 25483
rect 5089 25449 5123 25483
rect 5123 25449 5132 25483
rect 5080 25440 5132 25449
rect 7196 25483 7248 25492
rect 7196 25449 7205 25483
rect 7205 25449 7239 25483
rect 7239 25449 7248 25483
rect 7196 25440 7248 25449
rect 12256 25483 12308 25492
rect 12256 25449 12265 25483
rect 12265 25449 12299 25483
rect 12299 25449 12308 25483
rect 12256 25440 12308 25449
rect 7288 25372 7340 25424
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2872 24760 2924 24812
rect 3424 24735 3476 24744
rect 3424 24701 3433 24735
rect 3433 24701 3467 24735
rect 3467 24701 3476 24735
rect 3424 24692 3476 24701
rect 2780 24624 2832 24676
rect 2872 24599 2924 24608
rect 2872 24565 2881 24599
rect 2881 24565 2915 24599
rect 2915 24565 2924 24599
rect 2872 24556 2924 24565
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 11060 24556 11112 24608
rect 12072 24599 12124 24608
rect 12072 24565 12081 24599
rect 12081 24565 12115 24599
rect 12115 24565 12124 24599
rect 12072 24556 12124 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 3516 24012 3568 24064
rect 3976 24012 4028 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 11336 22108 11388 22160
rect 12164 22108 12216 22160
rect 4528 21879 4580 21888
rect 4528 21845 4537 21879
rect 4537 21845 4571 21879
rect 4571 21845 4580 21879
rect 4528 21836 4580 21845
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 3976 21632 4028 21684
rect 5264 21496 5316 21548
rect 4528 21428 4580 21480
rect 4896 21335 4948 21344
rect 4896 21301 4905 21335
rect 4905 21301 4939 21335
rect 4939 21301 4948 21335
rect 4896 21292 4948 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 4528 21088 4580 21140
rect 5540 21020 5592 21072
rect 6092 21020 6144 21072
rect 6736 20952 6788 21004
rect 6460 20816 6512 20868
rect 4896 20748 4948 20800
rect 5448 20748 5500 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 6092 20587 6144 20596
rect 6092 20553 6101 20587
rect 6101 20553 6135 20587
rect 6135 20553 6144 20587
rect 6092 20544 6144 20553
rect 9680 20519 9732 20528
rect 9680 20485 9689 20519
rect 9689 20485 9723 20519
rect 9723 20485 9732 20519
rect 9680 20476 9732 20485
rect 6460 20451 6512 20460
rect 6460 20417 6469 20451
rect 6469 20417 6503 20451
rect 6503 20417 6512 20451
rect 6460 20408 6512 20417
rect 6736 20340 6788 20392
rect 3332 20315 3384 20324
rect 3332 20281 3366 20315
rect 3366 20281 3384 20315
rect 3332 20272 3384 20281
rect 3976 20272 4028 20324
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 8208 20247 8260 20256
rect 8208 20213 8217 20247
rect 8217 20213 8251 20247
rect 8251 20213 8260 20247
rect 8576 20315 8628 20324
rect 8576 20281 8610 20315
rect 8610 20281 8628 20315
rect 8576 20272 8628 20281
rect 8208 20204 8260 20213
rect 9680 20204 9732 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 3332 20000 3384 20052
rect 5540 20043 5592 20052
rect 5540 20009 5549 20043
rect 5549 20009 5583 20043
rect 5583 20009 5592 20043
rect 5540 20000 5592 20009
rect 6736 20000 6788 20052
rect 7380 20000 7432 20052
rect 4436 19932 4488 19984
rect 4620 19932 4672 19984
rect 6092 19932 6144 19984
rect 7748 19932 7800 19984
rect 10048 19932 10100 19984
rect 7104 19864 7156 19916
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 5540 19728 5592 19780
rect 6828 19796 6880 19848
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 8576 19660 8628 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 3976 19456 4028 19508
rect 7380 19456 7432 19508
rect 7564 19456 7616 19508
rect 6000 19388 6052 19440
rect 5540 19252 5592 19304
rect 8576 19456 8628 19508
rect 10324 19320 10376 19372
rect 10508 19320 10560 19372
rect 5264 19116 5316 19168
rect 5724 19116 5776 19168
rect 7104 19252 7156 19304
rect 6552 19227 6604 19236
rect 6552 19193 6561 19227
rect 6561 19193 6595 19227
rect 6595 19193 6604 19227
rect 6552 19184 6604 19193
rect 8668 19184 8720 19236
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 9680 19116 9732 19125
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 5540 18955 5592 18964
rect 5540 18921 5549 18955
rect 5549 18921 5583 18955
rect 5583 18921 5592 18955
rect 5540 18912 5592 18921
rect 6000 18955 6052 18964
rect 6000 18921 6009 18955
rect 6009 18921 6043 18955
rect 6043 18921 6052 18955
rect 6000 18912 6052 18921
rect 6092 18912 6144 18964
rect 5816 18776 5868 18828
rect 6092 18776 6144 18828
rect 5632 18708 5684 18760
rect 6000 18708 6052 18760
rect 6828 18912 6880 18964
rect 7380 18912 7432 18964
rect 7748 18912 7800 18964
rect 6736 18776 6788 18828
rect 8392 18776 8444 18828
rect 5724 18640 5776 18692
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 5724 18368 5776 18420
rect 5724 18096 5776 18148
rect 6736 18096 6788 18148
rect 5632 18028 5684 18080
rect 6828 18028 6880 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 10048 13472 10100 13524
rect 9588 13336 9640 13388
rect 9680 13268 9732 13320
rect 9864 13268 9916 13320
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 10784 12928 10836 12980
rect 10048 12792 10100 12844
rect 10416 12724 10468 12776
rect 9588 12631 9640 12640
rect 9588 12597 9597 12631
rect 9597 12597 9631 12631
rect 9631 12597 9640 12631
rect 9588 12588 9640 12597
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 9956 12588 10008 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 6000 12180 6052 12232
rect 6736 12180 6788 12232
rect 8852 12044 8904 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 10416 11840 10468 11892
rect 7196 11704 7248 11756
rect 7380 11704 7432 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 7104 11568 7156 11620
rect 7380 11568 7432 11620
rect 8484 11568 8536 11620
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 8852 10956 8904 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 6828 10795 6880 10804
rect 6828 10761 6837 10795
rect 6837 10761 6871 10795
rect 6871 10761 6880 10795
rect 6828 10752 6880 10761
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 8484 10752 8536 10804
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 6920 10548 6972 10600
rect 8300 10548 8352 10600
rect 8484 10548 8536 10600
rect 6920 10412 6972 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 5908 10183 5960 10192
rect 5908 10149 5917 10183
rect 5917 10149 5951 10183
rect 5951 10149 5960 10183
rect 5908 10140 5960 10149
rect 6000 10183 6052 10192
rect 6000 10149 6009 10183
rect 6009 10149 6043 10183
rect 6043 10149 6052 10183
rect 8852 10208 8904 10260
rect 6920 10183 6972 10192
rect 6000 10140 6052 10149
rect 6920 10149 6929 10183
rect 6929 10149 6963 10183
rect 6963 10149 6972 10183
rect 7472 10183 7524 10192
rect 6920 10140 6972 10149
rect 7472 10149 7481 10183
rect 7481 10149 7515 10183
rect 7515 10149 7524 10183
rect 7472 10140 7524 10149
rect 6828 10004 6880 10056
rect 7012 10004 7064 10056
rect 8852 9868 8904 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 5908 9707 5960 9716
rect 5908 9673 5917 9707
rect 5917 9673 5951 9707
rect 5951 9673 5960 9707
rect 5908 9664 5960 9673
rect 7104 9664 7156 9716
rect 7472 9707 7524 9716
rect 7472 9673 7481 9707
rect 7481 9673 7515 9707
rect 7515 9673 7524 9707
rect 7472 9664 7524 9673
rect 5540 9596 5592 9648
rect 6000 9596 6052 9648
rect 6920 9324 6972 9376
rect 7012 9324 7064 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 6000 9120 6052 9172
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6920 8916 6972 8968
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 6000 8576 6052 8628
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 6920 8304 6972 8356
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 12440 7896 12492 7948
rect 13360 7896 13412 7948
rect 14004 7692 14056 7744
rect 14924 7692 14976 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 13820 7488 13872 7540
rect 15752 7488 15804 7540
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 4160 6808 4212 6860
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 5264 6604 5316 6656
rect 10416 6604 10468 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 4068 6332 4120 6384
rect 5540 6332 5592 6384
rect 10968 6264 11020 6316
rect 10232 6128 10284 6180
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 10968 5856 11020 5908
rect 9956 5763 10008 5772
rect 9956 5729 9990 5763
rect 9990 5729 10008 5763
rect 9956 5720 10008 5729
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 5540 5312 5592 5364
rect 8852 5312 8904 5364
rect 10416 5312 10468 5364
rect 9956 5176 10008 5228
rect 10784 5176 10836 5228
rect 9588 5108 9640 5160
rect 10048 5108 10100 5160
rect 11336 5108 11388 5160
rect 6920 5040 6972 5092
rect 10324 4972 10376 5024
rect 10600 4972 10652 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 10048 4768 10100 4820
rect 10232 4811 10284 4820
rect 10232 4777 10241 4811
rect 10241 4777 10275 4811
rect 10275 4777 10284 4811
rect 10232 4768 10284 4777
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 9956 4267 10008 4276
rect 9956 4233 9965 4267
rect 9965 4233 9999 4267
rect 9999 4233 10008 4267
rect 9956 4224 10008 4233
rect 9588 4156 9640 4208
rect 10692 4224 10744 4276
rect 4988 4088 5040 4140
rect 5448 4088 5500 4140
rect 5724 4088 5776 4140
rect 6644 4088 6696 4140
rect 10600 4088 10652 4140
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5080 3476 5132 3528
rect 9772 3476 9824 3528
rect 10968 3476 11020 3528
rect 4160 3408 4212 3460
rect 4528 3340 4580 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 4252 3136 4304 3188
rect 5080 3136 5132 3188
rect 5172 3136 5224 3188
rect 7288 3136 7340 3188
rect 2596 3068 2648 3120
rect 6092 3043 6144 3052
rect 3516 2932 3568 2984
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 7932 3136 7984 3188
rect 4620 2907 4672 2916
rect 4620 2873 4629 2907
rect 4629 2873 4663 2907
rect 4663 2873 4672 2907
rect 4620 2864 4672 2873
rect 2780 2796 2832 2848
rect 6920 2796 6972 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 3516 2567 3568 2576
rect 3516 2533 3525 2567
rect 3525 2533 3559 2567
rect 3559 2533 3568 2567
rect 3516 2524 3568 2533
rect 5448 2592 5500 2644
rect 7104 2592 7156 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 9588 2592 9640 2644
rect 1768 2320 1820 2372
rect 6552 2320 6604 2372
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39522 5410 40000
rect 5276 39520 5410 39522
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39522 10654 40000
rect 10598 39520 10732 39522
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39520 14242 40000
rect 14554 39520 14610 40000
rect 14922 39520 14978 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34950 244 39520
rect 204 34944 256 34950
rect 204 34886 256 34892
rect 584 34649 612 39520
rect 570 34640 626 34649
rect 570 34575 626 34584
rect 952 31521 980 39520
rect 1308 34944 1360 34950
rect 1308 34886 1360 34892
rect 1320 33266 1348 34886
rect 1412 34542 1440 39520
rect 1780 35057 1808 39520
rect 2148 35698 2176 39520
rect 2136 35692 2188 35698
rect 2136 35634 2188 35640
rect 1766 35048 1822 35057
rect 1766 34983 1822 34992
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 2608 33538 2636 39520
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 2424 33510 2636 33538
rect 1490 33416 1546 33425
rect 1490 33351 1546 33360
rect 1320 33238 1440 33266
rect 1412 32026 1440 33238
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 938 31512 994 31521
rect 938 31447 994 31456
rect 1504 27130 1532 33351
rect 1584 31884 1636 31890
rect 1584 31826 1636 31832
rect 1596 31142 1624 31826
rect 1584 31136 1636 31142
rect 1584 31078 1636 31084
rect 1492 27124 1544 27130
rect 1492 27066 1544 27072
rect 1596 10305 1624 31078
rect 2424 26314 2452 33510
rect 2700 31498 2728 35634
rect 2870 34640 2926 34649
rect 2870 34575 2926 34584
rect 2780 34536 2832 34542
rect 2780 34478 2832 34484
rect 2792 32570 2820 34478
rect 2780 32564 2832 32570
rect 2780 32506 2832 32512
rect 2884 32026 2912 34575
rect 2976 32065 3004 39520
rect 3344 35601 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3330 35592 3386 35601
rect 3330 35527 3386 35536
rect 3988 35193 4016 37182
rect 3974 35184 4030 35193
rect 3974 35119 4030 35128
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4172 34746 4200 39520
rect 4250 35048 4306 35057
rect 4250 34983 4306 34992
rect 4160 34740 4212 34746
rect 4160 34682 4212 34688
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3148 32360 3200 32366
rect 3148 32302 3200 32308
rect 2962 32056 3018 32065
rect 2872 32020 2924 32026
rect 2962 31991 3018 32000
rect 2872 31962 2924 31968
rect 2870 31512 2926 31521
rect 2700 31470 2820 31498
rect 2792 31414 2820 31470
rect 2870 31447 2872 31456
rect 2924 31447 2926 31456
rect 2872 31418 2924 31424
rect 2780 31408 2832 31414
rect 2780 31350 2832 31356
rect 2504 31136 2556 31142
rect 2504 31078 2556 31084
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 2318 9616 2374 9625
rect 2318 9551 2374 9560
rect 2134 3496 2190 3505
rect 2134 3431 2190 3440
rect 1398 3088 1454 3097
rect 1398 3023 1454 3032
rect 938 2952 994 2961
rect 938 2887 994 2896
rect 570 2816 626 2825
rect 570 2751 626 2760
rect 202 1456 258 1465
rect 202 1391 258 1400
rect 216 480 244 1391
rect 584 480 612 2751
rect 952 480 980 2887
rect 1412 480 1440 3023
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1780 480 1808 2314
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1872 1465 1900 2246
rect 1858 1456 1914 1465
rect 1858 1391 1914 1400
rect 2148 480 2176 3431
rect 2332 2650 2360 9551
rect 2516 9217 2544 31078
rect 2688 26784 2740 26790
rect 2740 26744 2820 26772
rect 2688 26726 2740 26732
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2502 9208 2558 9217
rect 2502 9143 2558 9152
rect 2608 8265 2636 26250
rect 2792 24682 2820 26744
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2780 24676 2832 24682
rect 2780 24618 2832 24624
rect 2884 24614 2912 24754
rect 2872 24608 2924 24614
rect 2872 24550 2924 24556
rect 2884 20097 2912 24550
rect 2870 20088 2926 20097
rect 2870 20023 2926 20032
rect 3160 19417 3188 32302
rect 4264 32026 4292 34983
rect 4540 32570 4568 39520
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 5000 32473 5028 39520
rect 5276 39494 5396 39520
rect 4986 32464 5042 32473
rect 4986 32399 5042 32408
rect 5080 32360 5132 32366
rect 5080 32302 5132 32308
rect 4252 32020 4304 32026
rect 4252 31962 4304 31968
rect 4160 31884 4212 31890
rect 4160 31826 4212 31832
rect 3240 31748 3292 31754
rect 3240 31690 3292 31696
rect 3252 31142 3280 31690
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 4172 31142 4200 31826
rect 3240 31136 3292 31142
rect 3240 31078 3292 31084
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 4160 31136 4212 31142
rect 4160 31078 4212 31084
rect 4988 31136 5040 31142
rect 4988 31078 5040 31084
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 3252 19281 3280 31078
rect 3344 20913 3372 31078
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3436 24750 3464 25434
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 24070 3556 24550
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3988 21690 4016 24006
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3330 20904 3386 20913
rect 3330 20839 3386 20848
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3974 20360 4030 20369
rect 3332 20324 3384 20330
rect 3974 20295 3976 20304
rect 3332 20266 3384 20272
rect 4028 20295 4030 20304
rect 3976 20266 4028 20272
rect 3344 20233 3372 20266
rect 3330 20224 3386 20233
rect 3330 20159 3386 20168
rect 3344 20058 3372 20159
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3988 19514 4016 20266
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3238 19272 3294 19281
rect 3238 19207 3294 19216
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 4080 15586 4108 30534
rect 4172 28966 4200 31078
rect 4342 30832 4398 30841
rect 4342 30767 4344 30776
rect 4396 30767 4398 30776
rect 4344 30738 4396 30744
rect 4356 30394 4384 30738
rect 4344 30388 4396 30394
rect 4344 30330 4396 30336
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 4620 28960 4672 28966
rect 4620 28902 4672 28908
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21486 4568 21830
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4540 21146 4568 21422
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 20097 4476 20198
rect 4434 20088 4490 20097
rect 4434 20023 4490 20032
rect 4632 19990 4660 28902
rect 4802 27976 4858 27985
rect 4802 27911 4858 27920
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4448 19394 4476 19926
rect 2976 15558 4108 15586
rect 4264 19366 4476 19394
rect 2594 8256 2650 8265
rect 2594 8191 2650 8200
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2608 480 2636 3062
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 2792 2854 2820 2887
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2976 480 3004 15558
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 3068 2650 3096 2751
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3344 480 3372 12271
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3528 3194 3556 8327
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3528 2990 3556 3130
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3516 2576 3568 2582
rect 3514 2544 3516 2553
rect 3568 2544 3570 2553
rect 3514 2479 3570 2488
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3988 1986 4016 15399
rect 4264 10169 4292 19366
rect 4816 18986 4844 27911
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25498 4936 25638
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 5000 23225 5028 31078
rect 5092 26874 5120 32302
rect 5170 32056 5226 32065
rect 5170 31991 5172 32000
rect 5224 31991 5226 32000
rect 5172 31962 5224 31968
rect 5172 31884 5224 31890
rect 5172 31826 5224 31832
rect 5184 31142 5212 31826
rect 5276 31249 5304 39494
rect 5448 34740 5500 34746
rect 5448 34682 5500 34688
rect 5460 31396 5488 34682
rect 5736 33017 5764 39520
rect 5906 34096 5962 34105
rect 5906 34031 5962 34040
rect 5722 33008 5778 33017
rect 5722 32943 5778 32952
rect 5540 31408 5592 31414
rect 5460 31368 5540 31396
rect 5540 31350 5592 31356
rect 5262 31240 5318 31249
rect 5262 31175 5318 31184
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 5092 26846 5212 26874
rect 5080 25900 5132 25906
rect 5080 25842 5132 25848
rect 5092 25498 5120 25842
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 5184 23361 5212 26846
rect 5814 26344 5870 26353
rect 5356 26308 5408 26314
rect 5814 26279 5870 26288
rect 5356 26250 5408 26256
rect 5368 25838 5396 26250
rect 5356 25832 5408 25838
rect 5356 25774 5408 25780
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 5170 23352 5226 23361
rect 5170 23287 5226 23296
rect 4986 23216 5042 23225
rect 4986 23151 5042 23160
rect 5276 21554 5304 25706
rect 5538 23352 5594 23361
rect 5538 23287 5594 23296
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 4908 20806 4936 21286
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 5276 20233 5304 21490
rect 5552 21078 5580 23287
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5552 20890 5580 21014
rect 5552 20862 5672 20890
rect 5448 20800 5500 20806
rect 5500 20748 5580 20754
rect 5448 20742 5580 20748
rect 5460 20726 5580 20742
rect 5262 20224 5318 20233
rect 5262 20159 5318 20168
rect 5276 19174 5304 20159
rect 5552 20058 5580 20726
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5552 19310 5580 19722
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 4816 18958 5488 18986
rect 5552 18970 5580 19246
rect 5354 14512 5410 14521
rect 5354 14447 5410 14456
rect 4250 10160 4306 10169
rect 4250 10095 4306 10104
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4068 6792 4120 6798
rect 4172 6769 4200 6802
rect 4068 6734 4120 6740
rect 4158 6760 4214 6769
rect 4080 6390 4108 6734
rect 4158 6695 4214 6704
rect 4172 6458 4200 6695
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4158 3496 4214 3505
rect 4158 3431 4160 3440
rect 4212 3431 4214 3440
rect 4160 3402 4212 3408
rect 4158 3224 4214 3233
rect 4264 3194 4292 8191
rect 5264 6656 5316 6662
rect 5262 6624 5264 6633
rect 5316 6624 5318 6633
rect 5262 6559 5318 6568
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4158 3159 4214 3168
rect 4252 3188 4304 3194
rect 3804 1958 4016 1986
rect 3804 480 3832 1958
rect 4172 480 4200 3159
rect 4252 3130 4304 3136
rect 4250 3088 4306 3097
rect 4250 3023 4306 3032
rect 4264 2650 4292 3023
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4540 480 4568 3334
rect 4618 2952 4674 2961
rect 4618 2887 4620 2896
rect 4672 2887 4674 2896
rect 4620 2858 4672 2864
rect 5000 480 5028 4082
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5092 3369 5120 3470
rect 5078 3360 5134 3369
rect 5078 3295 5134 3304
rect 5092 3194 5120 3295
rect 5184 3194 5212 3538
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5368 480 5396 14447
rect 5460 4146 5488 18958
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5644 18766 5672 20862
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5736 18698 5764 19110
rect 5828 18834 5856 26279
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5736 18426 5764 18634
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5552 6474 5580 9590
rect 5644 6769 5672 18022
rect 5630 6760 5686 6769
rect 5630 6695 5686 6704
rect 5552 6446 5672 6474
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5370 5580 6326
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 4729 5672 6446
rect 5630 4720 5686 4729
rect 5630 4655 5686 4664
rect 5736 4298 5764 18090
rect 5814 10568 5870 10577
rect 5814 10503 5870 10512
rect 5828 9178 5856 10503
rect 5920 10198 5948 34031
rect 6196 31793 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6776 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6748 31906 6776 37726
rect 6932 35850 6960 39520
rect 6840 35822 6960 35850
rect 6840 32026 6868 35822
rect 7194 35728 7250 35737
rect 7194 35663 7250 35672
rect 7102 35592 7158 35601
rect 7102 35527 7158 35536
rect 7012 32224 7064 32230
rect 7012 32166 7064 32172
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6932 31906 6960 31962
rect 6748 31878 6960 31906
rect 6182 31784 6238 31793
rect 6182 31719 6238 31728
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 6184 31136 6236 31142
rect 6184 31078 6236 31084
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 6104 20602 6132 21014
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6012 19446 6040 19790
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 6012 18970 6040 19382
rect 6104 18970 6132 19926
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 12238 6040 18702
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5998 10296 6054 10305
rect 5998 10231 6054 10240
rect 6012 10198 6040 10231
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5920 9722 5948 10134
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5920 9625 5948 9658
rect 6012 9654 6040 10134
rect 6000 9648 6052 9654
rect 5906 9616 5962 9625
rect 6000 9590 6052 9596
rect 5906 9551 5962 9560
rect 5998 9208 6054 9217
rect 5816 9172 5868 9178
rect 5998 9143 6000 9152
rect 5816 9114 5868 9120
rect 6052 9143 6054 9152
rect 6000 9114 6052 9120
rect 6012 8634 6040 9114
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6012 8537 6040 8570
rect 5998 8528 6054 8537
rect 5998 8463 6054 8472
rect 6104 4842 6132 18770
rect 6196 12753 6224 31078
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6642 29064 6698 29073
rect 6642 28999 6698 29008
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20505 6500 20810
rect 6458 20496 6514 20505
rect 6458 20431 6460 20440
rect 6512 20431 6514 20440
rect 6460 20402 6512 20408
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6550 19272 6606 19281
rect 6550 19207 6552 19216
rect 6604 19207 6606 19216
rect 6552 19178 6604 19184
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6182 9480 6238 9489
rect 6182 9415 6238 9424
rect 6196 9042 6224 9415
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8430 6224 8978
rect 6184 8424 6236 8430
rect 6182 8392 6184 8401
rect 6236 8392 6238 8401
rect 6182 8327 6238 8336
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6104 4814 6224 4842
rect 5552 4270 5764 4298
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5552 2666 5580 4270
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5460 2650 5580 2666
rect 5448 2644 5580 2650
rect 5500 2638 5580 2644
rect 5448 2586 5500 2592
rect 5736 480 5764 4082
rect 6090 3088 6146 3097
rect 6090 3023 6092 3032
rect 6144 3023 6146 3032
rect 6092 2994 6144 3000
rect 6196 480 6224 4814
rect 6656 4146 6684 28999
rect 6840 24857 6868 31214
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6932 26042 6960 26522
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 6826 24848 6882 24857
rect 6826 24783 6882 24792
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6748 20398 6776 20946
rect 6826 20496 6882 20505
rect 6826 20431 6882 20440
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6748 20058 6776 20334
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6840 19854 6868 20431
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6826 19408 6882 19417
rect 6826 19343 6882 19352
rect 6840 19258 6868 19343
rect 6840 19230 6960 19258
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6840 18850 6868 18906
rect 6932 18850 6960 19230
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6840 18822 6960 18850
rect 6748 18154 6776 18770
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6840 18086 6868 18822
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 7024 12345 7052 32166
rect 7116 31482 7144 35527
rect 7104 31476 7156 31482
rect 7104 31418 7156 31424
rect 7208 26874 7236 35663
rect 7286 35048 7342 35057
rect 7286 34983 7342 34992
rect 7116 26846 7236 26874
rect 7116 19922 7144 26846
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7208 26450 7236 26726
rect 7196 26444 7248 26450
rect 7196 26386 7248 26392
rect 7208 25498 7236 26386
rect 7300 25906 7328 34983
rect 7392 32337 7420 39520
rect 7470 32872 7526 32881
rect 7470 32807 7526 32816
rect 7484 32570 7512 32807
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7484 32366 7512 32506
rect 7472 32360 7524 32366
rect 7378 32328 7434 32337
rect 7472 32302 7524 32308
rect 7378 32263 7434 32272
rect 7656 32224 7708 32230
rect 7656 32166 7708 32172
rect 7380 31748 7432 31754
rect 7380 31690 7432 31696
rect 7392 31142 7420 31690
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7300 25430 7328 25842
rect 7392 25702 7420 31078
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7380 25696 7432 25702
rect 7380 25638 7432 25644
rect 7288 25424 7340 25430
rect 7288 25366 7340 25372
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7116 19310 7144 19858
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7010 12336 7066 12345
rect 7010 12271 7066 12280
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 7857 6776 12174
rect 7116 11626 7144 19246
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 6826 11520 6882 11529
rect 6826 11455 6882 11464
rect 6840 10810 6868 11455
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6932 10606 6960 10950
rect 6920 10600 6972 10606
rect 6918 10568 6920 10577
rect 6972 10568 6974 10577
rect 6918 10503 6974 10512
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6932 10198 6960 10406
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 7010 10160 7066 10169
rect 7010 10095 7066 10104
rect 7024 10062 7052 10095
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6840 9466 6868 9998
rect 6840 9438 6960 9466
rect 6932 9382 6960 9438
rect 7024 9382 7052 9998
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6932 8974 6960 9318
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8362 6960 8910
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6734 7848 6790 7857
rect 6734 7783 6790 7792
rect 6932 6633 6960 8298
rect 6918 6624 6974 6633
rect 6918 6559 6974 6568
rect 6932 5098 6960 6559
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6932 4826 6960 5034
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7024 4185 7052 9318
rect 7010 4176 7066 4185
rect 6644 4140 6696 4146
rect 7010 4111 7066 4120
rect 6644 4082 6696 4088
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6564 480 6592 2314
rect 6932 480 6960 2790
rect 7116 2650 7144 9658
rect 7208 3369 7236 11698
rect 7194 3360 7250 3369
rect 7194 3295 7250 3304
rect 7300 3194 7328 25366
rect 7392 22001 7420 25638
rect 7378 21992 7434 22001
rect 7378 21927 7434 21936
rect 7378 20904 7434 20913
rect 7378 20839 7434 20848
rect 7392 20058 7420 20839
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7392 19514 7420 19994
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7392 11762 7420 18906
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 3346 7420 11562
rect 7484 10198 7512 26862
rect 7564 26376 7616 26382
rect 7564 26318 7616 26324
rect 7576 25906 7604 26318
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7576 25702 7604 25842
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7576 25158 7604 25638
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7576 20505 7604 25094
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7576 10713 7604 19450
rect 7668 15473 7696 32166
rect 7760 31385 7788 39520
rect 7930 35592 7986 35601
rect 7930 35527 7986 35536
rect 7840 31884 7892 31890
rect 7840 31826 7892 31832
rect 7746 31376 7802 31385
rect 7746 31311 7802 31320
rect 7852 31142 7880 31826
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7746 20088 7802 20097
rect 7746 20023 7802 20032
rect 7760 19990 7788 20023
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7760 18970 7788 19926
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7654 15464 7710 15473
rect 7654 15399 7710 15408
rect 7852 13841 7880 31078
rect 7944 26586 7972 35527
rect 8022 34504 8078 34513
rect 8022 34439 8078 34448
rect 8036 26926 8064 34439
rect 8220 34105 8248 39520
rect 8588 35737 8616 39520
rect 8956 37210 8984 39520
rect 8772 37182 8984 37210
rect 8574 35728 8630 35737
rect 8574 35663 8630 35672
rect 8298 35184 8354 35193
rect 8298 35119 8354 35128
rect 8206 34096 8262 34105
rect 8206 34031 8262 34040
rect 8312 31482 8340 35119
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7838 13832 7894 13841
rect 7838 13767 7894 13776
rect 7562 10704 7618 10713
rect 7562 10639 7618 10648
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7484 9722 7512 10134
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7838 4584 7894 4593
rect 7838 4519 7894 4528
rect 7746 3496 7802 3505
rect 7746 3431 7802 3440
rect 7392 3318 7512 3346
rect 7378 3224 7434 3233
rect 7288 3188 7340 3194
rect 7378 3159 7434 3168
rect 7288 3130 7340 3136
rect 7286 2816 7342 2825
rect 7286 2751 7342 2760
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7300 2530 7328 2751
rect 7392 2650 7420 3159
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7484 2553 7512 3318
rect 7470 2544 7526 2553
rect 7300 2502 7420 2530
rect 7392 480 7420 2502
rect 7470 2479 7526 2488
rect 7760 480 7788 3431
rect 7852 2650 7880 4519
rect 7944 3194 7972 26522
rect 8206 20360 8262 20369
rect 8206 20295 8262 20304
rect 8220 20262 8248 20295
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8404 18834 8432 26862
rect 8576 20324 8628 20330
rect 8576 20266 8628 20272
rect 8588 19718 8616 20266
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19514 8616 19654
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8298 12744 8354 12753
rect 8298 12679 8354 12688
rect 8312 10810 8340 12679
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 10810 8524 11562
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8312 10606 8340 10746
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 5681 8524 10542
rect 8482 5672 8538 5681
rect 8482 5607 8538 5616
rect 8206 4720 8262 4729
rect 8206 4655 8262 4664
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8220 480 8248 4655
rect 8680 3482 8708 19178
rect 8772 9489 8800 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9310 34640 9366 34649
rect 9310 34575 9366 34584
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 9324 32570 9352 34575
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9324 32366 9352 32506
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9312 31136 9364 31142
rect 9312 31078 9364 31084
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 17921 9352 31078
rect 9416 26926 9444 39520
rect 9784 34513 9812 39520
rect 10046 35184 10102 35193
rect 10046 35119 10102 35128
rect 9770 34504 9826 34513
rect 9770 34439 9826 34448
rect 9770 33008 9826 33017
rect 9770 32943 9826 32952
rect 9678 31920 9734 31929
rect 9678 31855 9734 31864
rect 9692 31482 9720 31855
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9692 31278 9720 31418
rect 9680 31272 9732 31278
rect 9680 31214 9732 31220
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9692 29073 9720 29446
rect 9784 29238 9812 32943
rect 9862 32464 9918 32473
rect 9862 32399 9918 32408
rect 9876 32026 9904 32399
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9954 31240 10010 31249
rect 9954 31175 10010 31184
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9678 29064 9734 29073
rect 9678 28999 9734 29008
rect 9876 27985 9904 31078
rect 9968 30938 9996 31175
rect 9956 30932 10008 30938
rect 9956 30874 10008 30880
rect 10060 30326 10088 35119
rect 10048 30320 10100 30326
rect 10048 30262 10100 30268
rect 9956 30048 10008 30054
rect 9956 29990 10008 29996
rect 9862 27976 9918 27985
rect 9862 27911 9918 27920
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9770 23216 9826 23225
rect 9770 23151 9826 23160
rect 9680 20528 9732 20534
rect 9678 20496 9680 20505
rect 9732 20496 9734 20505
rect 9678 20431 9734 20440
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9692 19854 9720 20198
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9692 19174 9720 19790
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9310 17912 9366 17921
rect 9310 17847 9366 17856
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9600 12646 9628 13330
rect 9692 13326 9720 19110
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11558 8892 12038
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11665 9076 11698
rect 9600 11665 9628 12582
rect 9034 11656 9090 11665
rect 9034 11591 9090 11600
rect 9586 11656 9642 11665
rect 9586 11591 9642 11600
rect 8852 11552 8904 11558
rect 8850 11520 8852 11529
rect 8904 11520 8906 11529
rect 8850 11455 8906 11464
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8864 10470 8892 10950
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 10266 8892 10406
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8956 10010 8984 10610
rect 8864 9982 8984 10010
rect 9678 10024 9734 10033
rect 8864 9926 8892 9982
rect 9678 9959 9734 9968
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8758 9480 8814 9489
rect 8758 9415 8814 9424
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8588 3454 8708 3482
rect 8588 480 8616 3454
rect 8772 1986 8800 8327
rect 8864 5370 8892 9862
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9402 6760 9458 6769
rect 9402 6695 9458 6704
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8772 1958 8984 1986
rect 8956 480 8984 1958
rect 9416 480 9444 6695
rect 9692 5710 9720 9959
rect 9680 5704 9732 5710
rect 9600 5652 9680 5658
rect 9600 5646 9732 5652
rect 9600 5630 9720 5646
rect 9600 5166 9628 5630
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9678 4176 9734 4185
rect 9600 2650 9628 4150
rect 9678 4111 9734 4120
rect 9692 3346 9720 4111
rect 9784 3534 9812 23151
rect 9968 14521 9996 29990
rect 10152 26926 10180 39520
rect 10612 39494 10732 39520
rect 10230 34912 10286 34921
rect 10230 34847 10286 34856
rect 10244 29714 10272 34847
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10336 31142 10364 31826
rect 10704 31226 10732 39494
rect 10874 34776 10930 34785
rect 10874 34711 10930 34720
rect 10612 31198 10732 31226
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10428 30054 10456 30738
rect 10416 30048 10468 30054
rect 10416 29990 10468 29996
rect 10232 29708 10284 29714
rect 10232 29650 10284 29656
rect 10244 29306 10272 29650
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10232 29096 10284 29102
rect 10232 29038 10284 29044
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 10060 19174 10088 19926
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9954 14512 10010 14521
rect 9954 14447 10010 14456
rect 10060 13530 10088 19110
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9876 12646 9904 13262
rect 10060 12850 10088 13466
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9876 10033 9904 12582
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9968 6458 9996 12582
rect 10060 12442 10088 12786
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5234 9996 5714
rect 10060 5250 10088 10639
rect 10244 9625 10272 29038
rect 10428 28665 10456 29990
rect 10414 28656 10470 28665
rect 10414 28591 10470 28600
rect 10612 27062 10640 31198
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10336 19378 10364 26998
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10612 20097 10640 26862
rect 10704 23633 10732 31078
rect 10888 30326 10916 34711
rect 10980 30841 11008 39520
rect 11348 32881 11376 39520
rect 11808 37754 11836 39520
rect 11532 37726 11836 37754
rect 11532 34649 11560 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11518 34640 11574 34649
rect 11518 34575 11574 34584
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11334 32872 11390 32881
rect 11334 32807 11390 32816
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11058 31784 11114 31793
rect 11058 31719 11114 31728
rect 11072 30938 11100 31719
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 10966 30832 11022 30841
rect 10966 30767 11022 30776
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 10876 30320 10928 30326
rect 10876 30262 10928 30268
rect 11440 30054 11468 30738
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11428 30048 11480 30054
rect 11428 29990 11480 29996
rect 11072 26353 11100 29990
rect 11058 26344 11114 26353
rect 11058 26279 11114 26288
rect 11150 24848 11206 24857
rect 11150 24783 11206 24792
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 10690 23624 10746 23633
rect 10690 23559 10746 23568
rect 11072 20754 11100 24550
rect 10888 20726 11100 20754
rect 10888 20618 10916 20726
rect 10796 20590 10916 20618
rect 10598 20088 10654 20097
rect 10598 20023 10654 20032
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10428 12102 10456 12718
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11898 10456 12038
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 9956 5228 10008 5234
rect 10060 5222 10180 5250
rect 9956 5170 10008 5176
rect 9968 4282 9996 5170
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4826 10088 5102
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10060 4593 10088 4762
rect 10046 4584 10102 4593
rect 10046 4519 10102 4528
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9692 3318 9812 3346
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9784 480 9812 3318
rect 10152 480 10180 5222
rect 10244 4826 10272 6122
rect 10428 6118 10456 6598
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5370 10456 6054
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10336 4185 10364 4966
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10520 3097 10548 19314
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10704 6882 10732 13767
rect 10796 12986 10824 20590
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10966 11656 11022 11665
rect 10966 11591 11022 11600
rect 10612 6854 10732 6882
rect 10612 5030 10640 6854
rect 10980 6322 11008 11591
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5914 11008 6258
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10690 5128 10746 5137
rect 10690 5063 10746 5072
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10704 4826 10732 5063
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 4146 10640 4626
rect 10704 4282 10732 4762
rect 10796 4622 10824 5170
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11164 3482 11192 24783
rect 11336 22160 11388 22166
rect 11336 22102 11388 22108
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11256 3618 11284 17847
rect 11348 5166 11376 22102
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11440 4049 11468 29990
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12084 24614 12112 25298
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 12176 22166 12204 39520
rect 12544 35057 12572 39520
rect 12530 35048 12586 35057
rect 12530 34983 12586 34992
rect 12438 32328 12494 32337
rect 12438 32263 12494 32272
rect 12452 32026 12480 32263
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 12532 31408 12584 31414
rect 12530 31376 12532 31385
rect 12584 31376 12586 31385
rect 12530 31311 12586 31320
rect 12254 30016 12310 30025
rect 12254 29951 12310 29960
rect 12268 25498 12296 29951
rect 12438 28656 12494 28665
rect 12438 28591 12494 28600
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 12452 7954 12480 28591
rect 12530 23624 12586 23633
rect 12530 23559 12586 23568
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12438 7848 12494 7857
rect 12438 7783 12494 7792
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11426 4040 11482 4049
rect 11426 3975 11482 3984
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11256 3590 11560 3618
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 10598 2952 10654 2961
rect 10598 2887 10654 2896
rect 10612 480 10640 2887
rect 10980 480 11008 3470
rect 11164 3454 11376 3482
rect 11348 480 11376 3454
rect 11532 2530 11560 3590
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11532 2502 11836 2530
rect 11808 480 11836 2502
rect 12176 480 12204 5607
rect 12452 3210 12480 7783
rect 12544 3346 12572 23559
rect 12636 3505 12664 32166
rect 13004 31929 13032 39520
rect 13372 35193 13400 39520
rect 13358 35184 13414 35193
rect 13358 35119 13414 35128
rect 13082 35048 13138 35057
rect 13082 34983 13138 34992
rect 13096 32570 13124 34983
rect 13740 34921 13768 39520
rect 14200 37754 14228 39520
rect 14016 37726 14228 37754
rect 13726 34912 13782 34921
rect 13726 34847 13782 34856
rect 14016 34785 14044 37726
rect 14568 37618 14596 39520
rect 14108 37590 14596 37618
rect 14002 34776 14058 34785
rect 14002 34711 14058 34720
rect 13358 34640 13414 34649
rect 13358 34575 13414 34584
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 13096 32366 13124 32506
rect 13084 32360 13136 32366
rect 13084 32302 13136 32308
rect 12990 31920 13046 31929
rect 13372 31890 13400 34575
rect 12990 31855 13046 31864
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 13004 31142 13032 31690
rect 13372 31482 13400 31826
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 13004 3913 13032 31078
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 12990 3904 13046 3913
rect 12990 3839 13046 3848
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12544 3318 12664 3346
rect 12636 3210 12664 3318
rect 12452 3182 12572 3210
rect 12636 3182 13032 3210
rect 12544 480 12572 3182
rect 13004 480 13032 3182
rect 13372 480 13400 7890
rect 13556 2961 13584 31622
rect 14002 21992 14058 22001
rect 14002 21927 14058 21936
rect 13818 12472 13874 12481
rect 13818 12407 13874 12416
rect 13726 9616 13782 9625
rect 13726 9551 13782 9560
rect 13542 2952 13598 2961
rect 13542 2887 13598 2896
rect 13740 480 13768 9551
rect 13832 7546 13860 12407
rect 14016 7750 14044 21927
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14108 5137 14136 37590
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14936 35601 14964 39520
rect 14922 35592 14978 35601
rect 14922 35527 14978 35536
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 15396 34649 15424 39520
rect 15764 35057 15792 39520
rect 15750 35048 15806 35057
rect 15750 34983 15806 34992
rect 15382 34640 15438 34649
rect 15382 34575 15438 34584
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 14200 12481 14228 31214
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14186 12472 14242 12481
rect 14186 12407 14242 12416
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14094 5128 14150 5137
rect 14094 5063 14150 5072
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14186 4040 14242 4049
rect 14186 3975 14242 3984
rect 14200 480 14228 3975
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 1986 14688 4111
rect 14568 1958 14688 1986
rect 14568 480 14596 1958
rect 14936 480 14964 7686
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15396 480 15424 3839
rect 15764 480 15792 7482
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 570 34584 626 34640
rect 1766 34992 1822 35048
rect 1490 33360 1546 33416
rect 938 31456 994 31512
rect 2870 34584 2926 34640
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3330 35536 3386 35592
rect 3974 35128 4030 35184
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 4250 34992 4306 35048
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 2962 32000 3018 32056
rect 2870 31476 2926 31512
rect 2870 31456 2872 31476
rect 2872 31456 2924 31476
rect 2924 31456 2926 31476
rect 1582 10240 1638 10296
rect 2318 9560 2374 9616
rect 2134 3440 2190 3496
rect 1398 3032 1454 3088
rect 938 2896 994 2952
rect 570 2760 626 2816
rect 202 1400 258 1456
rect 1858 1400 1914 1456
rect 2502 9152 2558 9208
rect 2870 20032 2926 20088
rect 4986 32408 5042 32464
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3146 19352 3202 19408
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3330 20848 3386 20904
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3974 20324 4030 20360
rect 3974 20304 3976 20324
rect 3976 20304 4028 20324
rect 4028 20304 4030 20324
rect 3330 20168 3386 20224
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3238 19216 3294 19272
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 4342 30796 4398 30832
rect 4342 30776 4344 30796
rect 4344 30776 4396 30796
rect 4396 30776 4398 30796
rect 4434 20032 4490 20088
rect 4802 27920 4858 27976
rect 2594 8200 2650 8256
rect 2778 2896 2834 2952
rect 3974 15408 4030 15464
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3330 12280 3386 12336
rect 3054 2760 3110 2816
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3514 8336 3570 8392
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3514 2524 3516 2544
rect 3516 2524 3568 2544
rect 3568 2524 3570 2544
rect 3514 2488 3570 2524
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 5170 32020 5226 32056
rect 5170 32000 5172 32020
rect 5172 32000 5224 32020
rect 5224 32000 5226 32020
rect 5906 34040 5962 34096
rect 5722 32952 5778 33008
rect 5262 31184 5318 31240
rect 5814 26288 5870 26344
rect 5170 23296 5226 23352
rect 4986 23160 5042 23216
rect 5538 23296 5594 23352
rect 5262 20168 5318 20224
rect 5354 14456 5410 14512
rect 4250 10104 4306 10160
rect 4250 8200 4306 8256
rect 4158 6704 4214 6760
rect 4158 3460 4214 3496
rect 4158 3440 4160 3460
rect 4160 3440 4212 3460
rect 4212 3440 4214 3460
rect 4158 3168 4214 3224
rect 5262 6604 5264 6624
rect 5264 6604 5316 6624
rect 5316 6604 5318 6624
rect 5262 6568 5318 6604
rect 4250 3032 4306 3088
rect 4618 2916 4674 2952
rect 4618 2896 4620 2916
rect 4620 2896 4672 2916
rect 4672 2896 4674 2916
rect 5078 3304 5134 3360
rect 5630 6704 5686 6760
rect 5630 4664 5686 4720
rect 5814 10512 5870 10568
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 7194 35672 7250 35728
rect 7102 35536 7158 35592
rect 6182 31728 6238 31784
rect 5998 10240 6054 10296
rect 5906 9560 5962 9616
rect 5998 9172 6054 9208
rect 5998 9152 6000 9172
rect 6000 9152 6052 9172
rect 6052 9152 6054 9172
rect 5998 8472 6054 8528
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6642 29008 6698 29064
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6458 20460 6514 20496
rect 6458 20440 6460 20460
rect 6460 20440 6512 20460
rect 6512 20440 6514 20460
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6550 19236 6606 19272
rect 6550 19216 6552 19236
rect 6552 19216 6604 19236
rect 6604 19216 6606 19236
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6182 12688 6238 12744
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6182 9424 6238 9480
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6182 8372 6184 8392
rect 6184 8372 6236 8392
rect 6236 8372 6238 8392
rect 6182 8336 6238 8372
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6090 3052 6146 3088
rect 6090 3032 6092 3052
rect 6092 3032 6144 3052
rect 6144 3032 6146 3052
rect 6826 24792 6882 24848
rect 6826 20440 6882 20496
rect 6826 19352 6882 19408
rect 7286 34992 7342 35048
rect 7470 32816 7526 32872
rect 7378 32272 7434 32328
rect 7010 12280 7066 12336
rect 6826 11464 6882 11520
rect 6918 10548 6920 10568
rect 6920 10548 6972 10568
rect 6972 10548 6974 10568
rect 6918 10512 6974 10548
rect 7010 10104 7066 10160
rect 6734 7792 6790 7848
rect 6918 6568 6974 6624
rect 7010 4120 7066 4176
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7194 3304 7250 3360
rect 7378 21936 7434 21992
rect 7378 20848 7434 20904
rect 7562 20440 7618 20496
rect 7930 35536 7986 35592
rect 7746 31320 7802 31376
rect 7746 20032 7802 20088
rect 7654 15408 7710 15464
rect 8022 34448 8078 34504
rect 8574 35672 8630 35728
rect 8298 35128 8354 35184
rect 8206 34040 8262 34096
rect 7838 13776 7894 13832
rect 7562 10648 7618 10704
rect 7838 4528 7894 4584
rect 7746 3440 7802 3496
rect 7378 3168 7434 3224
rect 7286 2760 7342 2816
rect 7470 2488 7526 2544
rect 8206 20304 8262 20360
rect 8298 12688 8354 12744
rect 8482 5616 8538 5672
rect 8206 4664 8262 4720
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 9310 34584 9366 34640
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 10046 35128 10102 35184
rect 9770 34448 9826 34504
rect 9770 32952 9826 33008
rect 9678 31864 9734 31920
rect 9862 32408 9918 32464
rect 9954 31184 10010 31240
rect 9678 29008 9734 29064
rect 9862 27920 9918 27976
rect 9770 23160 9826 23216
rect 9678 20476 9680 20496
rect 9680 20476 9732 20496
rect 9732 20476 9734 20496
rect 9678 20440 9734 20476
rect 9310 17856 9366 17912
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 9034 11600 9090 11656
rect 9586 11600 9642 11656
rect 8850 11500 8852 11520
rect 8852 11500 8904 11520
rect 8904 11500 8906 11520
rect 8850 11464 8906 11500
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 9678 9968 9734 10024
rect 8758 9424 8814 9480
rect 8758 8336 8814 8392
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 9402 6704 9458 6760
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9678 4120 9734 4176
rect 10230 34856 10286 34912
rect 10874 34720 10930 34776
rect 9954 14456 10010 14512
rect 9862 9968 9918 10024
rect 10046 10648 10102 10704
rect 10414 28600 10470 28656
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11518 34584 11574 34640
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11334 32816 11390 32872
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11058 31728 11114 31784
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 10966 30776 11022 30832
rect 11058 26288 11114 26344
rect 11150 24792 11206 24848
rect 10690 23568 10746 23624
rect 10598 20032 10654 20088
rect 10230 9560 10286 9616
rect 10046 4528 10102 4584
rect 10322 4120 10378 4176
rect 10690 13776 10746 13832
rect 10966 11600 11022 11656
rect 10690 5072 10746 5128
rect 11242 17856 11298 17912
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 12530 34992 12586 35048
rect 12438 32272 12494 32328
rect 12530 31356 12532 31376
rect 12532 31356 12584 31376
rect 12584 31356 12586 31376
rect 12530 31320 12586 31356
rect 12254 29960 12310 30016
rect 12438 28600 12494 28656
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 12530 23568 12586 23624
rect 12438 7792 12494 7848
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 12162 5616 12218 5672
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11426 3984 11482 4040
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 10506 3032 10562 3088
rect 10598 2896 10654 2952
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 13358 35128 13414 35184
rect 13082 34992 13138 35048
rect 13726 34856 13782 34912
rect 14002 34720 14058 34776
rect 13358 34584 13414 34640
rect 12990 31864 13046 31920
rect 12990 3848 13046 3904
rect 12622 3440 12678 3496
rect 14002 21936 14058 21992
rect 13818 12416 13874 12472
rect 13726 9560 13782 9616
rect 13542 2896 13598 2952
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14922 35536 14978 35592
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 15750 34992 15806 35048
rect 15382 34584 15438 34640
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14186 12416 14242 12472
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14094 5072 14150 5128
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14646 4120 14702 4176
rect 14186 3984 14242 4040
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15382 3848 15438 3904
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 7189 35730 7255 35733
rect 8569 35730 8635 35733
rect 7189 35728 8635 35730
rect 7189 35672 7194 35728
rect 7250 35672 8574 35728
rect 8630 35672 8635 35728
rect 7189 35670 8635 35672
rect 7189 35667 7255 35670
rect 8569 35667 8635 35670
rect 3325 35594 3391 35597
rect 7097 35594 7163 35597
rect 3325 35592 7163 35594
rect 3325 35536 3330 35592
rect 3386 35536 7102 35592
rect 7158 35536 7163 35592
rect 3325 35534 7163 35536
rect 3325 35531 3391 35534
rect 7097 35531 7163 35534
rect 7925 35594 7991 35597
rect 14917 35594 14983 35597
rect 7925 35592 14983 35594
rect 7925 35536 7930 35592
rect 7986 35536 14922 35592
rect 14978 35536 14983 35592
rect 7925 35534 14983 35536
rect 7925 35531 7991 35534
rect 14917 35531 14983 35534
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3969 35186 4035 35189
rect 8293 35186 8359 35189
rect 3969 35184 8359 35186
rect 3969 35128 3974 35184
rect 4030 35128 8298 35184
rect 8354 35128 8359 35184
rect 3969 35126 8359 35128
rect 3969 35123 4035 35126
rect 8293 35123 8359 35126
rect 10041 35186 10107 35189
rect 13353 35186 13419 35189
rect 10041 35184 13419 35186
rect 10041 35128 10046 35184
rect 10102 35128 13358 35184
rect 13414 35128 13419 35184
rect 10041 35126 13419 35128
rect 10041 35123 10107 35126
rect 13353 35123 13419 35126
rect 1761 35050 1827 35053
rect 4245 35050 4311 35053
rect 1761 35048 4311 35050
rect 1761 34992 1766 35048
rect 1822 34992 4250 35048
rect 4306 34992 4311 35048
rect 1761 34990 4311 34992
rect 1761 34987 1827 34990
rect 4245 34987 4311 34990
rect 7281 35050 7347 35053
rect 12525 35050 12591 35053
rect 7281 35048 12591 35050
rect 7281 34992 7286 35048
rect 7342 34992 12530 35048
rect 12586 34992 12591 35048
rect 7281 34990 12591 34992
rect 7281 34987 7347 34990
rect 12525 34987 12591 34990
rect 13077 35050 13143 35053
rect 15745 35050 15811 35053
rect 13077 35048 15811 35050
rect 13077 34992 13082 35048
rect 13138 34992 15750 35048
rect 15806 34992 15811 35048
rect 13077 34990 15811 34992
rect 13077 34987 13143 34990
rect 15745 34987 15811 34990
rect 10225 34914 10291 34917
rect 13721 34914 13787 34917
rect 10225 34912 13787 34914
rect 10225 34856 10230 34912
rect 10286 34856 13726 34912
rect 13782 34856 13787 34912
rect 10225 34854 13787 34856
rect 10225 34851 10291 34854
rect 13721 34851 13787 34854
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 10869 34778 10935 34781
rect 13997 34778 14063 34781
rect 10869 34776 14063 34778
rect 10869 34720 10874 34776
rect 10930 34720 14002 34776
rect 14058 34720 14063 34776
rect 10869 34718 14063 34720
rect 10869 34715 10935 34718
rect 13997 34715 14063 34718
rect 565 34642 631 34645
rect 2865 34642 2931 34645
rect 565 34640 2931 34642
rect 565 34584 570 34640
rect 626 34584 2870 34640
rect 2926 34584 2931 34640
rect 565 34582 2931 34584
rect 565 34579 631 34582
rect 2865 34579 2931 34582
rect 9305 34642 9371 34645
rect 11513 34642 11579 34645
rect 9305 34640 11579 34642
rect 9305 34584 9310 34640
rect 9366 34584 11518 34640
rect 11574 34584 11579 34640
rect 9305 34582 11579 34584
rect 9305 34579 9371 34582
rect 11513 34579 11579 34582
rect 13353 34642 13419 34645
rect 15377 34642 15443 34645
rect 13353 34640 15443 34642
rect 13353 34584 13358 34640
rect 13414 34584 15382 34640
rect 15438 34584 15443 34640
rect 13353 34582 15443 34584
rect 13353 34579 13419 34582
rect 15377 34579 15443 34582
rect 8017 34506 8083 34509
rect 9765 34506 9831 34509
rect 8017 34504 9831 34506
rect 8017 34448 8022 34504
rect 8078 34448 9770 34504
rect 9826 34448 9831 34504
rect 8017 34446 9831 34448
rect 8017 34443 8083 34446
rect 9765 34443 9831 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 5901 34098 5967 34101
rect 8201 34098 8267 34101
rect 5901 34096 8267 34098
rect 5901 34040 5906 34096
rect 5962 34040 8206 34096
rect 8262 34040 8267 34096
rect 5901 34038 8267 34040
rect 5901 34035 5967 34038
rect 8201 34035 8267 34038
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 0 33418 480 33448
rect 1485 33418 1551 33421
rect 0 33416 1551 33418
rect 0 33360 1490 33416
rect 1546 33360 1551 33416
rect 0 33358 1551 33360
rect 0 33328 480 33358
rect 1485 33355 1551 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 5717 33010 5783 33013
rect 9765 33010 9831 33013
rect 5717 33008 9831 33010
rect 5717 32952 5722 33008
rect 5778 32952 9770 33008
rect 9826 32952 9831 33008
rect 5717 32950 9831 32952
rect 5717 32947 5783 32950
rect 9765 32947 9831 32950
rect 7465 32874 7531 32877
rect 11329 32874 11395 32877
rect 7465 32872 11395 32874
rect 7465 32816 7470 32872
rect 7526 32816 11334 32872
rect 11390 32816 11395 32872
rect 7465 32814 11395 32816
rect 7465 32811 7531 32814
rect 11329 32811 11395 32814
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 4981 32466 5047 32469
rect 9857 32466 9923 32469
rect 4981 32464 9923 32466
rect 4981 32408 4986 32464
rect 5042 32408 9862 32464
rect 9918 32408 9923 32464
rect 4981 32406 9923 32408
rect 4981 32403 5047 32406
rect 9857 32403 9923 32406
rect 7373 32330 7439 32333
rect 12433 32330 12499 32333
rect 7373 32328 12499 32330
rect 7373 32272 7378 32328
rect 7434 32272 12438 32328
rect 12494 32272 12499 32328
rect 7373 32270 12499 32272
rect 7373 32267 7439 32270
rect 12433 32267 12499 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 2957 32058 3023 32061
rect 5165 32058 5231 32061
rect 2957 32056 5231 32058
rect 2957 32000 2962 32056
rect 3018 32000 5170 32056
rect 5226 32000 5231 32056
rect 2957 31998 5231 32000
rect 2957 31995 3023 31998
rect 5165 31995 5231 31998
rect 9673 31922 9739 31925
rect 12985 31922 13051 31925
rect 9673 31920 13051 31922
rect 9673 31864 9678 31920
rect 9734 31864 12990 31920
rect 13046 31864 13051 31920
rect 9673 31862 13051 31864
rect 9673 31859 9739 31862
rect 12985 31859 13051 31862
rect 6177 31786 6243 31789
rect 11053 31786 11119 31789
rect 6177 31784 11119 31786
rect 6177 31728 6182 31784
rect 6238 31728 11058 31784
rect 11114 31728 11119 31784
rect 6177 31726 11119 31728
rect 6177 31723 6243 31726
rect 11053 31723 11119 31726
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 933 31514 999 31517
rect 2865 31514 2931 31517
rect 933 31512 2931 31514
rect 933 31456 938 31512
rect 994 31456 2870 31512
rect 2926 31456 2931 31512
rect 933 31454 2931 31456
rect 933 31451 999 31454
rect 2865 31451 2931 31454
rect 7741 31378 7807 31381
rect 12525 31378 12591 31381
rect 7741 31376 12591 31378
rect 7741 31320 7746 31376
rect 7802 31320 12530 31376
rect 12586 31320 12591 31376
rect 7741 31318 12591 31320
rect 7741 31315 7807 31318
rect 12525 31315 12591 31318
rect 5257 31242 5323 31245
rect 9949 31242 10015 31245
rect 5257 31240 10015 31242
rect 5257 31184 5262 31240
rect 5318 31184 9954 31240
rect 10010 31184 10015 31240
rect 5257 31182 10015 31184
rect 5257 31179 5323 31182
rect 9949 31179 10015 31182
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 4337 30834 4403 30837
rect 10961 30834 11027 30837
rect 4337 30832 11027 30834
rect 4337 30776 4342 30832
rect 4398 30776 10966 30832
rect 11022 30776 11027 30832
rect 4337 30774 11027 30776
rect 4337 30771 4403 30774
rect 10961 30771 11027 30774
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 12249 30018 12315 30021
rect 15520 30018 16000 30048
rect 12249 30016 16000 30018
rect 12249 29960 12254 30016
rect 12310 29960 16000 30016
rect 12249 29958 16000 29960
rect 12249 29955 12315 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6637 29066 6703 29069
rect 9673 29066 9739 29069
rect 6637 29064 9739 29066
rect 6637 29008 6642 29064
rect 6698 29008 9678 29064
rect 9734 29008 9739 29064
rect 6637 29006 9739 29008
rect 6637 29003 6703 29006
rect 9673 29003 9739 29006
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 10409 28658 10475 28661
rect 12433 28658 12499 28661
rect 10409 28656 12499 28658
rect 10409 28600 10414 28656
rect 10470 28600 12438 28656
rect 12494 28600 12499 28656
rect 10409 28598 12499 28600
rect 10409 28595 10475 28598
rect 12433 28595 12499 28598
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 4797 27978 4863 27981
rect 9857 27978 9923 27981
rect 4797 27976 9923 27978
rect 4797 27920 4802 27976
rect 4858 27920 9862 27976
rect 9918 27920 9923 27976
rect 4797 27918 9923 27920
rect 4797 27915 4863 27918
rect 9857 27915 9923 27918
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 5809 26346 5875 26349
rect 11053 26346 11119 26349
rect 5809 26344 11119 26346
rect 5809 26288 5814 26344
rect 5870 26288 11058 26344
rect 11114 26288 11119 26344
rect 5809 26286 11119 26288
rect 5809 26283 5875 26286
rect 11053 26283 11119 26286
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6821 24850 6887 24853
rect 11145 24850 11211 24853
rect 6821 24848 11211 24850
rect 6821 24792 6826 24848
rect 6882 24792 11150 24848
rect 11206 24792 11211 24848
rect 6821 24790 11211 24792
rect 6821 24787 6887 24790
rect 11145 24787 11211 24790
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 10685 23626 10751 23629
rect 12525 23626 12591 23629
rect 10685 23624 12591 23626
rect 10685 23568 10690 23624
rect 10746 23568 12530 23624
rect 12586 23568 12591 23624
rect 10685 23566 12591 23568
rect 10685 23563 10751 23566
rect 12525 23563 12591 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 5165 23354 5231 23357
rect 5533 23354 5599 23357
rect 5165 23352 5599 23354
rect 5165 23296 5170 23352
rect 5226 23296 5538 23352
rect 5594 23296 5599 23352
rect 5165 23294 5599 23296
rect 5165 23291 5231 23294
rect 5533 23291 5599 23294
rect 4981 23218 5047 23221
rect 9765 23218 9831 23221
rect 4981 23216 9831 23218
rect 4981 23160 4986 23216
rect 5042 23160 9770 23216
rect 9826 23160 9831 23216
rect 4981 23158 9831 23160
rect 4981 23155 5047 23158
rect 9765 23155 9831 23158
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 7373 21994 7439 21997
rect 13997 21994 14063 21997
rect 7373 21992 14063 21994
rect 7373 21936 7378 21992
rect 7434 21936 14002 21992
rect 14058 21936 14063 21992
rect 7373 21934 14063 21936
rect 7373 21931 7439 21934
rect 13997 21931 14063 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3325 20906 3391 20909
rect 7373 20906 7439 20909
rect 3325 20904 7439 20906
rect 3325 20848 3330 20904
rect 3386 20848 7378 20904
rect 7434 20848 7439 20904
rect 3325 20846 7439 20848
rect 3325 20843 3391 20846
rect 7373 20843 7439 20846
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 6453 20498 6519 20501
rect 6821 20498 6887 20501
rect 7557 20498 7623 20501
rect 9673 20498 9739 20501
rect 6453 20496 9739 20498
rect 6453 20440 6458 20496
rect 6514 20440 6826 20496
rect 6882 20440 7562 20496
rect 7618 20440 9678 20496
rect 9734 20440 9739 20496
rect 6453 20438 9739 20440
rect 6453 20435 6519 20438
rect 6821 20435 6887 20438
rect 7557 20435 7623 20438
rect 9673 20435 9739 20438
rect 3969 20362 4035 20365
rect 8201 20362 8267 20365
rect 3969 20360 8267 20362
rect 3969 20304 3974 20360
rect 4030 20304 8206 20360
rect 8262 20304 8267 20360
rect 3969 20302 8267 20304
rect 3969 20299 4035 20302
rect 8201 20299 8267 20302
rect 3325 20226 3391 20229
rect 5257 20226 5323 20229
rect 3325 20224 5323 20226
rect 3325 20168 3330 20224
rect 3386 20168 5262 20224
rect 5318 20168 5323 20224
rect 3325 20166 5323 20168
rect 3325 20163 3391 20166
rect 5257 20163 5323 20166
rect 6277 20160 6597 20161
rect 0 20090 480 20120
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 2865 20090 2931 20093
rect 4429 20090 4495 20093
rect 0 20088 4495 20090
rect 0 20032 2870 20088
rect 2926 20032 4434 20088
rect 4490 20032 4495 20088
rect 0 20030 4495 20032
rect 0 20000 480 20030
rect 2865 20027 2931 20030
rect 4429 20027 4495 20030
rect 7741 20090 7807 20093
rect 10593 20090 10659 20093
rect 7741 20088 10659 20090
rect 7741 20032 7746 20088
rect 7802 20032 10598 20088
rect 10654 20032 10659 20088
rect 7741 20030 10659 20032
rect 7741 20027 7807 20030
rect 10593 20027 10659 20030
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 3141 19410 3207 19413
rect 6821 19410 6887 19413
rect 3141 19408 6887 19410
rect 3141 19352 3146 19408
rect 3202 19352 6826 19408
rect 6882 19352 6887 19408
rect 3141 19350 6887 19352
rect 3141 19347 3207 19350
rect 6821 19347 6887 19350
rect 3233 19274 3299 19277
rect 6545 19274 6611 19277
rect 3233 19272 6611 19274
rect 3233 19216 3238 19272
rect 3294 19216 6550 19272
rect 6606 19216 6611 19272
rect 3233 19214 6611 19216
rect 3233 19211 3299 19214
rect 6545 19211 6611 19214
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 9305 17914 9371 17917
rect 11237 17914 11303 17917
rect 9305 17912 11303 17914
rect 9305 17856 9310 17912
rect 9366 17856 11242 17912
rect 11298 17856 11303 17912
rect 9305 17854 11303 17856
rect 9305 17851 9371 17854
rect 11237 17851 11303 17854
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3969 15466 4035 15469
rect 7649 15466 7715 15469
rect 3969 15464 7715 15466
rect 3969 15408 3974 15464
rect 4030 15408 7654 15464
rect 7710 15408 7715 15464
rect 3969 15406 7715 15408
rect 3969 15403 4035 15406
rect 7649 15403 7715 15406
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 5349 14514 5415 14517
rect 9949 14514 10015 14517
rect 5349 14512 10015 14514
rect 5349 14456 5354 14512
rect 5410 14456 9954 14512
rect 10010 14456 10015 14512
rect 5349 14454 10015 14456
rect 5349 14451 5415 14454
rect 9949 14451 10015 14454
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 7833 13834 7899 13837
rect 10685 13834 10751 13837
rect 7833 13832 10751 13834
rect 7833 13776 7838 13832
rect 7894 13776 10690 13832
rect 10746 13776 10751 13832
rect 7833 13774 10751 13776
rect 7833 13771 7899 13774
rect 10685 13771 10751 13774
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 6177 12746 6243 12749
rect 8293 12746 8359 12749
rect 6177 12744 8359 12746
rect 6177 12688 6182 12744
rect 6238 12688 8298 12744
rect 8354 12688 8359 12744
rect 6177 12686 8359 12688
rect 6177 12683 6243 12686
rect 8293 12683 8359 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 13813 12474 13879 12477
rect 14181 12474 14247 12477
rect 13813 12472 14247 12474
rect 13813 12416 13818 12472
rect 13874 12416 14186 12472
rect 14242 12416 14247 12472
rect 13813 12414 14247 12416
rect 13813 12411 13879 12414
rect 14181 12411 14247 12414
rect 3325 12338 3391 12341
rect 7005 12338 7071 12341
rect 3325 12336 7071 12338
rect 3325 12280 3330 12336
rect 3386 12280 7010 12336
rect 7066 12280 7071 12336
rect 3325 12278 7071 12280
rect 3325 12275 3391 12278
rect 7005 12275 7071 12278
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 9029 11658 9095 11661
rect 9581 11658 9647 11661
rect 10961 11658 11027 11661
rect 9029 11656 11027 11658
rect 9029 11600 9034 11656
rect 9090 11600 9586 11656
rect 9642 11600 10966 11656
rect 11022 11600 11027 11656
rect 9029 11598 11027 11600
rect 9029 11595 9095 11598
rect 9581 11595 9647 11598
rect 10961 11595 11027 11598
rect 6821 11522 6887 11525
rect 8845 11522 8911 11525
rect 6821 11520 8911 11522
rect 6821 11464 6826 11520
rect 6882 11464 8850 11520
rect 8906 11464 8911 11520
rect 6821 11462 8911 11464
rect 6821 11459 6887 11462
rect 8845 11459 8911 11462
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 7557 10706 7623 10709
rect 10041 10706 10107 10709
rect 7557 10704 10107 10706
rect 7557 10648 7562 10704
rect 7618 10648 10046 10704
rect 10102 10648 10107 10704
rect 7557 10646 10107 10648
rect 7557 10643 7623 10646
rect 10041 10643 10107 10646
rect 5809 10570 5875 10573
rect 6913 10570 6979 10573
rect 5809 10568 6979 10570
rect 5809 10512 5814 10568
rect 5870 10512 6918 10568
rect 6974 10512 6979 10568
rect 5809 10510 6979 10512
rect 5809 10507 5875 10510
rect 6913 10507 6979 10510
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 1577 10298 1643 10301
rect 5993 10298 6059 10301
rect 1577 10296 6059 10298
rect 1577 10240 1582 10296
rect 1638 10240 5998 10296
rect 6054 10240 6059 10296
rect 1577 10238 6059 10240
rect 1577 10235 1643 10238
rect 5993 10235 6059 10238
rect 4245 10162 4311 10165
rect 7005 10162 7071 10165
rect 4245 10160 7071 10162
rect 4245 10104 4250 10160
rect 4306 10104 7010 10160
rect 7066 10104 7071 10160
rect 4245 10102 7071 10104
rect 4245 10099 4311 10102
rect 7005 10099 7071 10102
rect 9673 10026 9739 10029
rect 9857 10026 9923 10029
rect 15520 10026 16000 10056
rect 9673 10024 16000 10026
rect 9673 9968 9678 10024
rect 9734 9968 9862 10024
rect 9918 9968 16000 10024
rect 9673 9966 16000 9968
rect 9673 9963 9739 9966
rect 9857 9963 9923 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 2313 9618 2379 9621
rect 5901 9618 5967 9621
rect 2313 9616 5967 9618
rect 2313 9560 2318 9616
rect 2374 9560 5906 9616
rect 5962 9560 5967 9616
rect 2313 9558 5967 9560
rect 2313 9555 2379 9558
rect 5901 9555 5967 9558
rect 10225 9618 10291 9621
rect 13721 9618 13787 9621
rect 10225 9616 13787 9618
rect 10225 9560 10230 9616
rect 10286 9560 13726 9616
rect 13782 9560 13787 9616
rect 10225 9558 13787 9560
rect 10225 9555 10291 9558
rect 13721 9555 13787 9558
rect 6177 9482 6243 9485
rect 8753 9482 8819 9485
rect 6177 9480 8819 9482
rect 6177 9424 6182 9480
rect 6238 9424 8758 9480
rect 8814 9424 8819 9480
rect 6177 9422 8819 9424
rect 6177 9419 6243 9422
rect 8753 9419 8819 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 2497 9210 2563 9213
rect 5993 9210 6059 9213
rect 2497 9208 6059 9210
rect 2497 9152 2502 9208
rect 2558 9152 5998 9208
rect 6054 9152 6059 9208
rect 2497 9150 6059 9152
rect 2497 9147 2563 9150
rect 5993 9147 6059 9150
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 5993 8530 6059 8533
rect 5993 8528 6378 8530
rect 5993 8472 5998 8528
rect 6054 8472 6378 8528
rect 5993 8470 6378 8472
rect 5993 8467 6059 8470
rect 3509 8394 3575 8397
rect 6177 8394 6243 8397
rect 3509 8392 6243 8394
rect 3509 8336 3514 8392
rect 3570 8336 6182 8392
rect 6238 8336 6243 8392
rect 3509 8334 6243 8336
rect 6318 8394 6378 8470
rect 8753 8394 8819 8397
rect 6318 8392 8819 8394
rect 6318 8336 8758 8392
rect 8814 8336 8819 8392
rect 6318 8334 8819 8336
rect 3509 8331 3575 8334
rect 6177 8331 6243 8334
rect 8753 8331 8819 8334
rect 2589 8258 2655 8261
rect 4245 8258 4311 8261
rect 2589 8256 4311 8258
rect 2589 8200 2594 8256
rect 2650 8200 4250 8256
rect 4306 8200 4311 8256
rect 2589 8198 4311 8200
rect 2589 8195 2655 8198
rect 4245 8195 4311 8198
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 6729 7850 6795 7853
rect 12433 7850 12499 7853
rect 6729 7848 12499 7850
rect 6729 7792 6734 7848
rect 6790 7792 12438 7848
rect 12494 7792 12499 7848
rect 6729 7790 12499 7792
rect 6729 7787 6795 7790
rect 12433 7787 12499 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 0 6762 480 6792
rect 4153 6762 4219 6765
rect 0 6760 4219 6762
rect 0 6704 4158 6760
rect 4214 6704 4219 6760
rect 0 6702 4219 6704
rect 0 6672 480 6702
rect 4153 6699 4219 6702
rect 5625 6762 5691 6765
rect 9397 6762 9463 6765
rect 5625 6760 9463 6762
rect 5625 6704 5630 6760
rect 5686 6704 9402 6760
rect 9458 6704 9463 6760
rect 5625 6702 9463 6704
rect 5625 6699 5691 6702
rect 9397 6699 9463 6702
rect 5257 6626 5323 6629
rect 6913 6626 6979 6629
rect 5257 6624 6979 6626
rect 5257 6568 5262 6624
rect 5318 6568 6918 6624
rect 6974 6568 6979 6624
rect 5257 6566 6979 6568
rect 5257 6563 5323 6566
rect 6913 6563 6979 6566
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 8477 5674 8543 5677
rect 12157 5674 12223 5677
rect 8477 5672 12223 5674
rect 8477 5616 8482 5672
rect 8538 5616 12162 5672
rect 12218 5616 12223 5672
rect 8477 5614 12223 5616
rect 8477 5611 8543 5614
rect 12157 5611 12223 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 10685 5130 10751 5133
rect 14089 5130 14155 5133
rect 10685 5128 14155 5130
rect 10685 5072 10690 5128
rect 10746 5072 14094 5128
rect 14150 5072 14155 5128
rect 10685 5070 14155 5072
rect 10685 5067 10751 5070
rect 14089 5067 14155 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 5625 4722 5691 4725
rect 8201 4722 8267 4725
rect 5625 4720 8267 4722
rect 5625 4664 5630 4720
rect 5686 4664 8206 4720
rect 8262 4664 8267 4720
rect 5625 4662 8267 4664
rect 5625 4659 5691 4662
rect 8201 4659 8267 4662
rect 7833 4586 7899 4589
rect 10041 4586 10107 4589
rect 7833 4584 10107 4586
rect 7833 4528 7838 4584
rect 7894 4528 10046 4584
rect 10102 4528 10107 4584
rect 7833 4526 10107 4528
rect 7833 4523 7899 4526
rect 10041 4523 10107 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 7005 4178 7071 4181
rect 9673 4178 9739 4181
rect 7005 4176 9739 4178
rect 7005 4120 7010 4176
rect 7066 4120 9678 4176
rect 9734 4120 9739 4176
rect 7005 4118 9739 4120
rect 7005 4115 7071 4118
rect 9673 4115 9739 4118
rect 10317 4178 10383 4181
rect 14641 4178 14707 4181
rect 10317 4176 14707 4178
rect 10317 4120 10322 4176
rect 10378 4120 14646 4176
rect 14702 4120 14707 4176
rect 10317 4118 14707 4120
rect 10317 4115 10383 4118
rect 14641 4115 14707 4118
rect 11421 4042 11487 4045
rect 14181 4042 14247 4045
rect 11421 4040 14247 4042
rect 11421 3984 11426 4040
rect 11482 3984 14186 4040
rect 14242 3984 14247 4040
rect 11421 3982 14247 3984
rect 11421 3979 11487 3982
rect 14181 3979 14247 3982
rect 12985 3906 13051 3909
rect 15377 3906 15443 3909
rect 12985 3904 15443 3906
rect 12985 3848 12990 3904
rect 13046 3848 15382 3904
rect 15438 3848 15443 3904
rect 12985 3846 15443 3848
rect 12985 3843 13051 3846
rect 15377 3843 15443 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 2129 3498 2195 3501
rect 4153 3498 4219 3501
rect 2129 3496 4219 3498
rect 2129 3440 2134 3496
rect 2190 3440 4158 3496
rect 4214 3440 4219 3496
rect 2129 3438 4219 3440
rect 2129 3435 2195 3438
rect 4153 3435 4219 3438
rect 7741 3498 7807 3501
rect 12617 3498 12683 3501
rect 7741 3496 12683 3498
rect 7741 3440 7746 3496
rect 7802 3440 12622 3496
rect 12678 3440 12683 3496
rect 7741 3438 12683 3440
rect 7741 3435 7807 3438
rect 12617 3435 12683 3438
rect 5073 3362 5139 3365
rect 7189 3362 7255 3365
rect 5073 3360 7255 3362
rect 5073 3304 5078 3360
rect 5134 3304 7194 3360
rect 7250 3304 7255 3360
rect 5073 3302 7255 3304
rect 5073 3299 5139 3302
rect 7189 3299 7255 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 4153 3226 4219 3229
rect 7373 3226 7439 3229
rect 4153 3224 7439 3226
rect 4153 3168 4158 3224
rect 4214 3168 7378 3224
rect 7434 3168 7439 3224
rect 4153 3166 7439 3168
rect 4153 3163 4219 3166
rect 7373 3163 7439 3166
rect 1393 3090 1459 3093
rect 4245 3090 4311 3093
rect 1393 3088 4311 3090
rect 1393 3032 1398 3088
rect 1454 3032 4250 3088
rect 4306 3032 4311 3088
rect 1393 3030 4311 3032
rect 1393 3027 1459 3030
rect 4245 3027 4311 3030
rect 6085 3090 6151 3093
rect 10501 3090 10567 3093
rect 6085 3088 10567 3090
rect 6085 3032 6090 3088
rect 6146 3032 10506 3088
rect 10562 3032 10567 3088
rect 6085 3030 10567 3032
rect 6085 3027 6151 3030
rect 10501 3027 10567 3030
rect 933 2954 999 2957
rect 2773 2954 2839 2957
rect 933 2952 2839 2954
rect 933 2896 938 2952
rect 994 2896 2778 2952
rect 2834 2896 2839 2952
rect 933 2894 2839 2896
rect 933 2891 999 2894
rect 2773 2891 2839 2894
rect 4613 2954 4679 2957
rect 10593 2954 10659 2957
rect 13537 2954 13603 2957
rect 4613 2952 10659 2954
rect 4613 2896 4618 2952
rect 4674 2896 10598 2952
rect 10654 2896 10659 2952
rect 4613 2894 10659 2896
rect 4613 2891 4679 2894
rect 10593 2891 10659 2894
rect 10734 2952 13603 2954
rect 10734 2896 13542 2952
rect 13598 2896 13603 2952
rect 10734 2894 13603 2896
rect 565 2818 631 2821
rect 3049 2818 3115 2821
rect 565 2816 3115 2818
rect 565 2760 570 2816
rect 626 2760 3054 2816
rect 3110 2760 3115 2816
rect 565 2758 3115 2760
rect 565 2755 631 2758
rect 3049 2755 3115 2758
rect 7281 2818 7347 2821
rect 10734 2818 10794 2894
rect 13537 2891 13603 2894
rect 7281 2816 10794 2818
rect 7281 2760 7286 2816
rect 7342 2760 10794 2816
rect 7281 2758 10794 2760
rect 7281 2755 7347 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 3509 2546 3575 2549
rect 7465 2546 7531 2549
rect 3509 2544 7531 2546
rect 3509 2488 3514 2544
rect 3570 2488 7470 2544
rect 7526 2488 7531 2544
rect 3509 2486 7531 2488
rect 3509 2483 3575 2486
rect 7465 2483 7531 2486
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 197 1458 263 1461
rect 1853 1458 1919 1461
rect 197 1456 1919 1458
rect 197 1400 202 1456
rect 258 1400 1858 1456
rect 1914 1400 1919 1456
rect 197 1398 1919 1400
rect 197 1395 263 1398
rect 1853 1395 1919 1398
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__decap_3  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2760 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14
timestamp 1604666999
transform 1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604666999
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604666999
transform 1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1604666999
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604666999
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1604666999
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604666999
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604666999
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604666999
transform 1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1604666999
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1604666999
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604666999
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604666999
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 1604666999
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1604666999
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1604666999
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604666999
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604666999
transform 1 0 5060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_55 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_51
timestamp 1604666999
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5888 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604666999
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604666999
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604666999
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_66
timestamp 1604666999
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604666999
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604666999
transform 1 0 7176 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1604666999
transform 1 0 7912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1604666999
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604666999
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604666999
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1604666999
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604666999
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1604666999
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86
timestamp 1604666999
transform 1 0 9016 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1604666999
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1604666999
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1604666999
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_106
timestamp 1604666999
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1604666999
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp 1604666999
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_36
timestamp 1604666999
transform 1 0 4416 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_48
timestamp 1604666999
transform 1 0 5520 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_60
timestamp 1604666999
transform 1 0 6624 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1604666999
transform 1 0 7728 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1604666999
transform 1 0 9752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_97
timestamp 1604666999
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _02_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_101
timestamp 1604666999
transform 1 0 10396 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1604666999
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_109
timestamp 1604666999
transform 1 0 11132 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1604666999
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp 1604666999
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_64
timestamp 1604666999
transform 1 0 6992 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_76
timestamp 1604666999
transform 1 0 8096 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1604666999
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1604666999
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_108
timestamp 1604666999
transform 1 0 11040 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_120
timestamp 1604666999
transform 1 0 12144 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_132
timestamp 1604666999
transform 1 0 13248 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1604666999
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604666999
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_81
timestamp 1604666999
transform 1 0 8556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1604666999
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1604666999
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_104
timestamp 1604666999
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1604666999
transform 1 0 11040 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp 1604666999
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1604666999
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1604666999
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1604666999
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_50
timestamp 1604666999
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 9936 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1604666999
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_112
timestamp 1604666999
transform 1 0 11408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1604666999
transform 1 0 10764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1604666999
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_124
timestamp 1604666999
transform 1 0 12512 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_136
timestamp 1604666999
transform 1 0 13616 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604666999
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1604666999
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp 1604666999
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_51
timestamp 1604666999
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_63
timestamp 1604666999
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_75
timestamp 1604666999
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1604666999
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604666999
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_98
timestamp 1604666999
transform 1 0 10120 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_110
timestamp 1604666999
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_122
timestamp 1604666999
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_134
timestamp 1604666999
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604666999
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604666999
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604666999
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604666999
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604666999
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604666999
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604666999
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604666999
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604666999
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604666999
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604666999
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604666999
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604666999
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1604666999
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_60
timestamp 1604666999
transform 1 0 6624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_72
timestamp 1604666999
transform 1 0 7728 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604666999
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604666999
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604666999
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1604666999
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1604666999
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604666999
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1604666999
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_47
timestamp 1604666999
transform 1 0 5428 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_57
timestamp 1604666999
transform 1 0 6348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1604666999
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1604666999
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1604666999
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1604666999
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp 1604666999
transform 1 0 6716 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_67
timestamp 1604666999
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7084 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1604666999
transform 1 0 8280 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1604666999
transform 1 0 7912 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604666999
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_75
timestamp 1604666999
transform 1 0 8004 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1604666999
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1604666999
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_81
timestamp 1604666999
transform 1 0 8556 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604666999
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1604666999
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1604666999
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604666999
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604666999
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604666999
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604666999
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604666999
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1604666999
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604666999
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604666999
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_71
timestamp 1604666999
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_88
timestamp 1604666999
transform 1 0 9200 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_100
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_112
timestamp 1604666999
transform 1 0 11408 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1604666999
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1604666999
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604666999
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1604666999
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_64
timestamp 1604666999
transform 1 0 6992 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_76
timestamp 1604666999
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_81
timestamp 1604666999
transform 1 0 8556 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1604666999
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604666999
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604666999
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1604666999
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604666999
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604666999
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_70
timestamp 1604666999
transform 1 0 7544 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1604666999
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_88
timestamp 1604666999
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1604666999
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1604666999
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1604666999
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1604666999
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604666999
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_68
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_76
timestamp 1604666999
transform 1 0 8096 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_81
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1604666999
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_99
timestamp 1604666999
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_103
timestamp 1604666999
transform 1 0 10580 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_115
timestamp 1604666999
transform 1 0 11684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1604666999
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_139
timestamp 1604666999
transform 1 0 13892 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604666999
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604666999
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604666999
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604666999
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1604666999
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1604666999
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1604666999
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1604666999
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604666999
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 10120 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_19_106
timestamp 1604666999
transform 1 0 10856 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604666999
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604666999
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1604666999
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1604666999
transform 1 0 14076 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604666999
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604666999
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604666999
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604666999
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604666999
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604666999
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1604666999
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1604666999
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604666999
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604666999
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604666999
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604666999
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604666999
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604666999
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604666999
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604666999
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604666999
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604666999
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_143
timestamp 1604666999
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604666999
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604666999
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604666999
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604666999
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604666999
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604666999
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604666999
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1604666999
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604666999
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604666999
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604666999
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604666999
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604666999
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604666999
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604666999
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604666999
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604666999
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604666999
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604666999
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604666999
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604666999
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1604666999
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1604666999
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604666999
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604666999
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604666999
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1604666999
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6440 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_51
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_56
timestamp 1604666999
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604666999
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_66
timestamp 1604666999
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_78
timestamp 1604666999
transform 1 0 8280 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_90
timestamp 1604666999
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_102
timestamp 1604666999
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1604666999
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6440 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_50
timestamp 1604666999
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1604666999
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604666999
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_71
timestamp 1604666999
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1604666999
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604666999
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604666999
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604666999
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604666999
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1604666999
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1604666999
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 3956 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1604666999
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_50
timestamp 1604666999
transform 1 0 5704 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_54
timestamp 1604666999
transform 1 0 6072 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604666999
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_75
timestamp 1604666999
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_79
timestamp 1604666999
transform 1 0 8372 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1604666999
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1604666999
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_99
timestamp 1604666999
transform 1 0 10212 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1604666999
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604666999
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1604666999
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1604666999
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5520 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1604666999
transform 1 0 6348 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7084 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1604666999
transform 1 0 6716 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1604666999
transform 1 0 6992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1604666999
transform 1 0 7912 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604666999
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_112
timestamp 1604666999
transform 1 0 11408 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_124
timestamp 1604666999
transform 1 0 12512 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_136
timestamp 1604666999
transform 1 0 13616 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1604666999
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 3036 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_38
timestamp 1604666999
transform 1 0 4600 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_48
timestamp 1604666999
transform 1 0 5520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_40
timestamp 1604666999
transform 1 0 4784 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_50
timestamp 1604666999
transform 1 0 5704 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_55
timestamp 1604666999
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1604666999
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5980 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8280 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1604666999
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_62
timestamp 1604666999
transform 1 0 6808 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_74
timestamp 1604666999
transform 1 0 7912 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_97
timestamp 1604666999
transform 1 0 10028 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1604666999
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_109
timestamp 1604666999
transform 1 0 11132 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604666999
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1604666999
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_143
timestamp 1604666999
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4416 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_33
timestamp 1604666999
transform 1 0 4140 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_45
timestamp 1604666999
transform 1 0 5244 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1604666999
transform 1 0 6348 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604666999
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604666999
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1604666999
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_143
timestamp 1604666999
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604666999
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_38
timestamp 1604666999
transform 1 0 4600 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_50
timestamp 1604666999
transform 1 0 5704 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_62
timestamp 1604666999
transform 1 0 6808 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_74
timestamp 1604666999
transform 1 0 7912 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_86
timestamp 1604666999
transform 1 0 9016 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604666999
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604666999
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604666999
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1604666999
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1604666999
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604666999
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604666999
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604666999
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604666999
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604666999
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604666999
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1604666999
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604666999
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604666999
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604666999
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604666999
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604666999
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604666999
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1604666999
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604666999
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_15
timestamp 1604666999
transform 1 0 2484 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604666999
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1604666999
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604666999
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604666999
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604666999
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604666999
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604666999
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604666999
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604666999
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_143
timestamp 1604666999
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1604666999
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1604666999
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3036 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1604666999
transform 1 0 3864 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1604666999
transform 1 0 4968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_54
timestamp 1604666999
transform 1 0 6072 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1604666999
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604666999
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604666999
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604666999
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12052 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_110
timestamp 1604666999
transform 1 0 11224 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_118
timestamp 1604666999
transform 1 0 11960 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1604666999
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_143
timestamp 1604666999
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_15
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_23
timestamp 1604666999
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_40
timestamp 1604666999
transform 1 0 4784 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604666999
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604666999
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7176 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7544 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_64
timestamp 1604666999
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_68
timestamp 1604666999
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_72
timestamp 1604666999
transform 1 0 7728 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_84
timestamp 1604666999
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 12052 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1604666999
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1604666999
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_122
timestamp 1604666999
transform 1 0 12328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_134
timestamp 1604666999
transform 1 0 13432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604666999
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604666999
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604666999
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604666999
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_39
timestamp 1604666999
transform 1 0 4692 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4968 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1604666999
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1604666999
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7820 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp 1604666999
transform 1 0 7636 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_75
timestamp 1604666999
transform 1 0 8004 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_87
timestamp 1604666999
transform 1 0 9108 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1604666999
transform 1 0 10212 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_111
timestamp 1604666999
transform 1 0 11316 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_119
timestamp 1604666999
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1604666999
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1604666999
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604666999
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_143
timestamp 1604666999
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604666999
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604666999
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604666999
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604666999
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_32
timestamp 1604666999
transform 1 0 4048 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4968 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_40
timestamp 1604666999
transform 1 0 4784 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1604666999
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_56
timestamp 1604666999
transform 1 0 6256 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6808 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1604666999
transform 1 0 7636 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_83
timestamp 1604666999
transform 1 0 8740 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1604666999
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1604666999
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1604666999
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1604666999
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1604666999
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604666999
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1604666999
transform 1 0 14076 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1604666999
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604666999
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_6
timestamp 1604666999
transform 1 0 1656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_10
timestamp 1604666999
transform 1 0 2024 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_22
timestamp 1604666999
transform 1 0 3128 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_34
timestamp 1604666999
transform 1 0 4232 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_46
timestamp 1604666999
transform 1 0 5336 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_58
timestamp 1604666999
transform 1 0 6440 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _03_
timestamp 1604666999
transform 1 0 7084 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_62
timestamp 1604666999
transform 1 0 6808 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_68
timestamp 1604666999
transform 1 0 7360 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_80
timestamp 1604666999
transform 1 0 8464 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_92
timestamp 1604666999
transform 1 0 9568 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_104
timestamp 1604666999
transform 1 0 10672 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_116
timestamp 1604666999
transform 1 0 11776 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604666999
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604666999
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604666999
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604666999
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604666999
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604666999
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604666999
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604666999
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1604666999
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604666999
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1604666999
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1604666999
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1604666999
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1604666999
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1604666999
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1604666999
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1604666999
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1604666999
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1604666999
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1604666999
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_74
timestamp 1604666999
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1604666999
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1604666999
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_86
timestamp 1604666999
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_98
timestamp 1604666999
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1604666999
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1604666999
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_110
timestamp 1604666999
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1604666999
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604666999
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604666999
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604666999
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604666999
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1604666999
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1604666999
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604666999
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604666999
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1604666999
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1604666999
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1604666999
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1604666999
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1604666999
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1604666999
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1604666999
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1604666999
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1604666999
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1604666999
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1604666999
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1604666999
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604666999
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1604666999
transform 1 0 14076 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1604666999
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604666999
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1604666999
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1604666999
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1604666999
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1604666999
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_51
timestamp 1604666999
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_59
timestamp 1604666999
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1604666999
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_74
timestamp 1604666999
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1604666999
transform 1 0 10212 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604666999
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_86
timestamp 1604666999
transform 1 0 9016 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_94
timestamp 1604666999
transform 1 0 9752 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1604666999
transform 1 0 10764 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_103
timestamp 1604666999
transform 1 0 10580 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_107
timestamp 1604666999
transform 1 0 10948 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_119
timestamp 1604666999
transform 1 0 12052 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604666999
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1604666999
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604666999
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1604666999
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604666999
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1604666999
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1604666999
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1604666999
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1604666999
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1604666999
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1604666999
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1604666999
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604666999
transform 1 0 10212 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_80
timestamp 1604666999
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_93
timestamp 1604666999
transform 1 0 9660 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_103
timestamp 1604666999
transform 1 0 10580 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_115
timestamp 1604666999
transform 1 0 11684 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_127
timestamp 1604666999
transform 1 0 12788 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604666999
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_139
timestamp 1604666999
transform 1 0 13892 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1604666999
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604666999
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1604666999
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1604666999
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604666999
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_27
timestamp 1604666999
transform 1 0 3588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_37
timestamp 1604666999
transform 1 0 4508 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_49
timestamp 1604666999
transform 1 0 5612 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1604666999
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_74
timestamp 1604666999
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604666999
transform 1 0 9752 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604666999
transform 1 0 9568 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_86
timestamp 1604666999
transform 1 0 9016 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_98
timestamp 1604666999
transform 1 0 10120 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604666999
transform 1 0 10856 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1604666999
transform 1 0 10304 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1604666999
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604666999
transform 1 0 10672 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_102
timestamp 1604666999
transform 1 0 10488 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1604666999
transform 1 0 11224 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_114
timestamp 1604666999
transform 1 0 11592 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604666999
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1604666999
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604666999
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1604666999
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604666999
transform 1 0 2668 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604666999
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604666999
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604666999
transform 1 0 1564 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604666999
transform 1 0 2484 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604666999
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1604666999
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1604666999
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_7
timestamp 1604666999
transform 1 0 1748 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_25
timestamp 1604666999
transform 1 0 3404 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_21
timestamp 1604666999
transform 1 0 3036 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1604666999
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1604666999
transform 1 0 3588 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604666999
transform 1 0 3220 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1604666999
transform 1 0 3772 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_37
timestamp 1604666999
transform 1 0 4508 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_33
timestamp 1604666999
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_32
timestamp 1604666999
transform 1 0 4048 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604666999
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604666999
transform 1 0 4324 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_39
timestamp 1604666999
transform 1 0 4692 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1604666999
transform 1 0 5612 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1604666999
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604666999
transform 1 0 5152 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604666999
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_51
timestamp 1604666999
transform 1 0 5796 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_43
timestamp 1604666999
transform 1 0 5060 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_46
timestamp 1604666999
transform 1 0 5336 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1604666999
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1604666999
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604666999
transform 1 0 6808 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1604666999
transform 1 0 7820 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604666999
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_63
timestamp 1604666999
transform 1 0 6900 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_75
timestamp 1604666999
transform 1 0 8004 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_66
timestamp 1604666999
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_70
timestamp 1604666999
transform 1 0 7544 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_75
timestamp 1604666999
transform 1 0 8004 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_86
timestamp 1604666999
transform 1 0 9016 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_81
timestamp 1604666999
transform 1 0 8556 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_87
timestamp 1604666999
transform 1 0 9108 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1604666999
transform 1 0 9200 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1604666999
transform 1 0 8648 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_90
timestamp 1604666999
transform 1 0 9384 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_93
timestamp 1604666999
transform 1 0 9660 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1604666999
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604666999
transform 1 0 9568 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604666999
transform 1 0 9752 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1604666999
transform 1 0 9752 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_98
timestamp 1604666999
transform 1 0 10120 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_98
timestamp 1604666999
transform 1 0 10120 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1604666999
transform 1 0 10856 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1604666999
transform 1 0 10304 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_110
timestamp 1604666999
transform 1 0 11224 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_102
timestamp 1604666999
transform 1 0 10488 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_114
timestamp 1604666999
transform 1 0 11592 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_127
timestamp 1604666999
transform 1 0 12788 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604666999
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604666999
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1604666999
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_131
timestamp 1604666999
transform 1 0 13156 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604666999
transform 1 0 13340 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604666999
transform 1 0 12972 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_134
timestamp 1604666999
transform 1 0 13432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_122
timestamp 1604666999
transform 1 0 12328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604666999
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604666999
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_143
timestamp 1604666999
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604666999
transform 1 0 2668 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604666999
transform 1 0 1564 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604666999
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1604666999
transform 1 0 1380 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_9
timestamp 1604666999
transform 1 0 1932 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604666999
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_21
timestamp 1604666999
transform 1 0 3036 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1604666999
transform 1 0 3772 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_36
timestamp 1604666999
transform 1 0 4416 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604666999
transform 1 0 5152 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_48
timestamp 1604666999
transform 1 0 5520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1604666999
transform 1 0 7820 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604666999
transform 1 0 6624 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_64
timestamp 1604666999
transform 1 0 6992 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_72
timestamp 1604666999
transform 1 0 7728 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_77
timestamp 1604666999
transform 1 0 8188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1604666999
transform 1 0 9660 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_89
timestamp 1604666999
transform 1 0 9292 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1604666999
transform 1 0 10028 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1604666999
transform 1 0 11132 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604666999
transform 1 0 13340 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604666999
transform 1 0 12236 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_125
timestamp 1604666999
transform 1 0 12604 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_137
timestamp 1604666999
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604666999
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1604666999
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604666999
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1604666999
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_15
timestamp 1604666999
transform 1 0 2484 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604666999
transform 1 0 3128 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604666999
transform 1 0 3680 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_21
timestamp 1604666999
transform 1 0 3036 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_26
timestamp 1604666999
transform 1 0 3496 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_30
timestamp 1604666999
transform 1 0 3864 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_38
timestamp 1604666999
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1604666999
transform 1 0 4784 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1604666999
transform 1 0 5336 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_44
timestamp 1604666999
transform 1 0 5152 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_48
timestamp 1604666999
transform 1 0 5520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604666999
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604666999
transform 1 0 7360 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_60
timestamp 1604666999
transform 1 0 6624 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_66
timestamp 1604666999
transform 1 0 7176 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1604666999
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604666999
transform 1 0 8648 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604666999
transform 1 0 9200 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_86
timestamp 1604666999
transform 1 0 9016 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_90
timestamp 1604666999
transform 1 0 9384 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_102
timestamp 1604666999
transform 1 0 10488 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_114
timestamp 1604666999
transform 1 0 11592 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604666999
transform 1 0 12420 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604666999
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_127
timestamp 1604666999
transform 1 0 12788 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_131
timestamp 1604666999
transform 1 0 13156 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604666999
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_143
timestamp 1604666999
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604666999
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604666999
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1604666999
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1604666999
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1604666999
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1604666999
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1604666999
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1604666999
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1604666999
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1604666999
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1604666999
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_117
timestamp 1604666999
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_129
timestamp 1604666999
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604666999
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1604666999
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1604666999
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604666999
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1604666999
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1604666999
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1604666999
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1604666999
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1604666999
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1604666999
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1604666999
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1604666999
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1604666999
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_98
timestamp 1604666999
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_110
timestamp 1604666999
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1604666999
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1604666999
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604666999
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_143
timestamp 1604666999
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604666999
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1604666999
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1604666999
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1604666999
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1604666999
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1604666999
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1604666999
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1604666999
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_80
timestamp 1604666999
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1604666999
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1604666999
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_117
timestamp 1604666999
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_129
timestamp 1604666999
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604666999
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1604666999
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1604666999
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604666999
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604666999
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1604666999
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1604666999
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1604666999
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1604666999
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1604666999
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1604666999
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604666999
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1604666999
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1604666999
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1604666999
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1604666999
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1604666999
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1604666999
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1604666999
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1604666999
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1604666999
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1604666999
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1604666999
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1604666999
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1604666999
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1604666999
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1604666999
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1604666999
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1604666999
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1604666999
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604666999
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604666999
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_143
timestamp 1604666999
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1604666999
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1604666999
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604666999
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604666999
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604666999
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604666999
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1604666999
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1604666999
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1604666999
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1604666999
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1604666999
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1604666999
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1604666999
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1604666999
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604666999
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604666999
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604666999
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604666999
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604666999
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604666999
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604666999
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604666999
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604666999
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604666999
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1604666999
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1604666999
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1604666999
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604666999
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604666999
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604666999
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604666999
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604666999
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604666999
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604666999
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604666999
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604666999
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604666999
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604666999
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604666999
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604666999
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604666999
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604666999
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604666999
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604666999
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604666999
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604666999
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604666999
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604666999
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604666999
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604666999
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604666999
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604666999
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604666999
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604666999
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604666999
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604666999
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604666999
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604666999
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604666999
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604666999
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604666999
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604666999
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604666999
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604666999
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604666999
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604666999
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604666999
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 6672 480 6792 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 20000 480 20120 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 33328 480 33448 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 prog_clk
port 83 nsew default input
rlabel metal3 s 15520 29928 16000 30048 6 right_grid_pin_52_
port 84 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 85 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 86 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
