VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__1_
  CLASS BLOCK ;
  FOREIGN sb_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 112.730 BY 123.450 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.400 4.040 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 121.050 3.130 123.450 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 121.050 8.650 123.450 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 3.440 112.730 4.040 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END bottom_right_grid_pin_11_
  PIN bottom_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 18.400 112.730 19.000 ;
    END
  END bottom_right_grid_pin_13_
  PIN bottom_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 2.400 ;
    END
  END bottom_right_grid_pin_15_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 121.050 14.630 123.450 ;
    END
  END bottom_right_grid_pin_1_
  PIN bottom_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END bottom_right_grid_pin_3_
  PIN bottom_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 10.920 112.730 11.520 ;
    END
  END bottom_right_grid_pin_5_
  PIN bottom_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END bottom_right_grid_pin_7_
  PIN bottom_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.330 121.050 20.610 123.450 ;
    END
  END bottom_right_grid_pin_9_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 26.560 112.730 27.160 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 34.040 112.730 34.640 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 41.520 112.730 42.120 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 121.050 26.590 123.450 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 2.400 51.640 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 121.050 32.570 123.450 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 121.050 38.550 123.450 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 49.680 112.730 50.280 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 57.160 112.730 57.760 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 121.050 44.530 123.450 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 65.320 112.730 65.920 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 121.050 50.510 123.450 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 121.050 56.490 123.450 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 72.800 112.730 73.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 121.050 62.010 123.450 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 80.280 112.730 80.880 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 121.050 67.990 123.450 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 88.440 112.730 89.040 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.400 86.320 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 121.050 73.970 123.450 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 121.050 79.950 123.450 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 121.050 85.930 123.450 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 121.050 91.910 123.450 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.330 95.920 112.730 96.520 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 121.050 97.890 123.450 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 2.400 99.920 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 121.050 103.870 123.450 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 2.400 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 2.400 ;
    END
  END left_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 121.050 109.850 123.450 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 103.400 112.730 104.000 ;
    END
  END top_right_grid_pin_11_
  PIN top_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 111.560 112.730 112.160 ;
    END
  END top_right_grid_pin_13_
  PIN top_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.330 119.040 112.730 119.640 ;
    END
  END top_right_grid_pin_15_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END top_right_grid_pin_1_
  PIN top_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END top_right_grid_pin_3_
  PIN top_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 2.400 120.320 ;
    END
  END top_right_grid_pin_5_
  PIN top_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END top_right_grid_pin_7_
  PIN top_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END top_right_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 23.510 10.640 25.110 111.760 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 42.295 10.640 43.895 111.760 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 107.180 111.605 ;
      LAYER met1 ;
        RECT 0.070 0.380 110.790 121.340 ;
      LAYER met2 ;
        RECT 0.090 120.770 2.570 121.450 ;
        RECT 3.410 120.770 8.090 121.450 ;
        RECT 8.930 120.770 14.070 121.450 ;
        RECT 14.910 120.770 20.050 121.450 ;
        RECT 20.890 120.770 26.030 121.450 ;
        RECT 26.870 120.770 32.010 121.450 ;
        RECT 32.850 120.770 37.990 121.450 ;
        RECT 38.830 120.770 43.970 121.450 ;
        RECT 44.810 120.770 49.950 121.450 ;
        RECT 50.790 120.770 55.930 121.450 ;
        RECT 56.770 120.770 61.450 121.450 ;
        RECT 62.290 120.770 67.430 121.450 ;
        RECT 68.270 120.770 73.410 121.450 ;
        RECT 74.250 120.770 79.390 121.450 ;
        RECT 80.230 120.770 85.370 121.450 ;
        RECT 86.210 120.770 91.350 121.450 ;
        RECT 92.190 120.770 97.330 121.450 ;
        RECT 98.170 120.770 103.310 121.450 ;
        RECT 104.150 120.770 109.290 121.450 ;
        RECT 110.130 120.770 110.770 121.450 ;
        RECT 0.090 2.680 110.770 120.770 ;
        RECT 0.090 0.155 1.650 2.680 ;
        RECT 2.490 0.155 5.330 2.680 ;
        RECT 6.170 0.155 9.010 2.680 ;
        RECT 9.850 0.155 12.690 2.680 ;
        RECT 13.530 0.155 16.370 2.680 ;
        RECT 17.210 0.155 20.050 2.680 ;
        RECT 20.890 0.155 24.190 2.680 ;
        RECT 25.030 0.155 27.870 2.680 ;
        RECT 28.710 0.155 31.550 2.680 ;
        RECT 32.390 0.155 35.230 2.680 ;
        RECT 36.070 0.155 38.910 2.680 ;
        RECT 39.750 0.155 42.590 2.680 ;
        RECT 43.430 0.155 46.730 2.680 ;
        RECT 47.570 0.155 50.410 2.680 ;
        RECT 51.250 0.155 54.090 2.680 ;
        RECT 54.930 0.155 57.770 2.680 ;
        RECT 58.610 0.155 61.450 2.680 ;
        RECT 62.290 0.155 65.130 2.680 ;
        RECT 65.970 0.155 69.270 2.680 ;
        RECT 70.110 0.155 72.950 2.680 ;
        RECT 73.790 0.155 76.630 2.680 ;
        RECT 77.470 0.155 80.310 2.680 ;
        RECT 81.150 0.155 83.990 2.680 ;
        RECT 84.830 0.155 87.670 2.680 ;
        RECT 88.510 0.155 91.810 2.680 ;
        RECT 92.650 0.155 95.490 2.680 ;
        RECT 96.330 0.155 99.170 2.680 ;
        RECT 100.010 0.155 102.850 2.680 ;
        RECT 103.690 0.155 106.530 2.680 ;
        RECT 107.370 0.155 110.210 2.680 ;
      LAYER met3 ;
        RECT 0.270 118.640 109.930 119.040 ;
        RECT 0.270 113.920 111.050 118.640 ;
        RECT 2.800 112.560 111.050 113.920 ;
        RECT 2.800 112.520 109.930 112.560 ;
        RECT 0.270 111.160 109.930 112.520 ;
        RECT 0.270 107.120 111.050 111.160 ;
        RECT 2.800 105.720 111.050 107.120 ;
        RECT 0.270 104.400 111.050 105.720 ;
        RECT 0.270 103.000 109.930 104.400 ;
        RECT 0.270 100.320 111.050 103.000 ;
        RECT 2.800 98.920 111.050 100.320 ;
        RECT 0.270 96.920 111.050 98.920 ;
        RECT 0.270 95.520 109.930 96.920 ;
        RECT 0.270 93.520 111.050 95.520 ;
        RECT 2.800 92.120 111.050 93.520 ;
        RECT 0.270 89.440 111.050 92.120 ;
        RECT 0.270 88.040 109.930 89.440 ;
        RECT 0.270 86.720 111.050 88.040 ;
        RECT 2.800 85.320 111.050 86.720 ;
        RECT 0.270 81.280 111.050 85.320 ;
        RECT 0.270 79.920 109.930 81.280 ;
        RECT 2.800 79.880 109.930 79.920 ;
        RECT 2.800 78.520 111.050 79.880 ;
        RECT 0.270 73.800 111.050 78.520 ;
        RECT 0.270 73.120 109.930 73.800 ;
        RECT 2.800 72.400 109.930 73.120 ;
        RECT 2.800 71.720 111.050 72.400 ;
        RECT 0.270 66.320 111.050 71.720 ;
        RECT 2.800 64.920 109.930 66.320 ;
        RECT 0.270 58.840 111.050 64.920 ;
        RECT 2.800 58.160 111.050 58.840 ;
        RECT 2.800 57.440 109.930 58.160 ;
        RECT 0.270 56.760 109.930 57.440 ;
        RECT 0.270 52.040 111.050 56.760 ;
        RECT 2.800 50.680 111.050 52.040 ;
        RECT 2.800 50.640 109.930 50.680 ;
        RECT 0.270 49.280 109.930 50.640 ;
        RECT 0.270 45.240 111.050 49.280 ;
        RECT 2.800 43.840 111.050 45.240 ;
        RECT 0.270 42.520 111.050 43.840 ;
        RECT 0.270 41.120 109.930 42.520 ;
        RECT 0.270 38.440 111.050 41.120 ;
        RECT 2.800 37.040 111.050 38.440 ;
        RECT 0.270 35.040 111.050 37.040 ;
        RECT 0.270 33.640 109.930 35.040 ;
        RECT 0.270 31.640 111.050 33.640 ;
        RECT 2.800 30.240 111.050 31.640 ;
        RECT 0.270 27.560 111.050 30.240 ;
        RECT 0.270 26.160 109.930 27.560 ;
        RECT 0.270 24.840 111.050 26.160 ;
        RECT 2.800 23.440 111.050 24.840 ;
        RECT 0.270 19.400 111.050 23.440 ;
        RECT 0.270 18.040 109.930 19.400 ;
        RECT 2.800 18.000 109.930 18.040 ;
        RECT 2.800 16.640 111.050 18.000 ;
        RECT 0.270 11.920 111.050 16.640 ;
        RECT 0.270 11.240 109.930 11.920 ;
        RECT 2.800 10.520 109.930 11.240 ;
        RECT 2.800 9.840 111.050 10.520 ;
        RECT 0.270 4.440 111.050 9.840 ;
        RECT 2.800 3.040 109.930 4.440 ;
        RECT 0.270 0.175 111.050 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.640 23.110 111.760 ;
        RECT 25.510 10.640 41.895 111.760 ;
        RECT 44.295 10.640 111.025 111.760 ;
  END
END sb_3__1_
END LIBRARY

