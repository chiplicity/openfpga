VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__2_
  CLASS BLOCK ;
  FOREIGN sb_0__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 137.600 70.290 140.000 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 68.040 140.000 68.640 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.760 140.000 105.360 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 107.480 140.000 108.080 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 110.880 140.000 111.480 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.280 140.000 114.880 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 117.680 140.000 118.280 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 124.480 140.000 125.080 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 127.880 140.000 128.480 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 131.280 140.000 131.880 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 71.440 140.000 72.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.160 140.000 74.760 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 77.560 140.000 78.160 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 84.360 140.000 84.960 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.760 140.000 88.360 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.160 140.000 91.760 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 94.560 140.000 95.160 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.960 140.000 98.560 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.720 140.000 35.320 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 37.440 140.000 38.040 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 40.840 140.000 41.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.640 140.000 48.240 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 51.040 140.000 51.640 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 54.440 140.000 55.040 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 57.840 140.000 58.440 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 61.240 140.000 61.840 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 64.640 140.000 65.240 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 7.520 140.000 8.120 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.920 140.000 11.520 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.320 140.000 14.920 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.720 140.000 18.320 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.120 140.000 21.720 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 24.520 140.000 25.120 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 27.920 140.000 28.520 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END prog_clk
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 134.680 140.000 135.280 ;
    END
  END right_top_grid_pin_1_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 4.670 2.760 134.320 133.580 ;
      LAYER met2 ;
        RECT 1.470 137.320 69.730 138.565 ;
        RECT 70.570 137.320 137.910 138.565 ;
        RECT 1.470 2.680 137.910 137.320 ;
        RECT 2.030 1.515 4.410 2.680 ;
        RECT 5.250 1.515 7.630 2.680 ;
        RECT 8.470 1.515 11.310 2.680 ;
        RECT 12.150 1.515 14.530 2.680 ;
        RECT 15.370 1.515 18.210 2.680 ;
        RECT 19.050 1.515 21.430 2.680 ;
        RECT 22.270 1.515 24.650 2.680 ;
        RECT 25.490 1.515 28.330 2.680 ;
        RECT 29.170 1.515 31.550 2.680 ;
        RECT 32.390 1.515 35.230 2.680 ;
        RECT 36.070 1.515 38.450 2.680 ;
        RECT 39.290 1.515 41.670 2.680 ;
        RECT 42.510 1.515 45.350 2.680 ;
        RECT 46.190 1.515 48.570 2.680 ;
        RECT 49.410 1.515 52.250 2.680 ;
        RECT 53.090 1.515 55.470 2.680 ;
        RECT 56.310 1.515 59.150 2.680 ;
        RECT 59.990 1.515 62.370 2.680 ;
        RECT 63.210 1.515 65.590 2.680 ;
        RECT 66.430 1.515 69.270 2.680 ;
        RECT 70.110 1.515 72.490 2.680 ;
        RECT 73.330 1.515 76.170 2.680 ;
        RECT 77.010 1.515 79.390 2.680 ;
        RECT 80.230 1.515 82.610 2.680 ;
        RECT 83.450 1.515 86.290 2.680 ;
        RECT 87.130 1.515 89.510 2.680 ;
        RECT 90.350 1.515 93.190 2.680 ;
        RECT 94.030 1.515 96.410 2.680 ;
        RECT 97.250 1.515 100.090 2.680 ;
        RECT 100.930 1.515 103.310 2.680 ;
        RECT 104.150 1.515 106.530 2.680 ;
        RECT 107.370 1.515 110.210 2.680 ;
        RECT 111.050 1.515 113.430 2.680 ;
        RECT 114.270 1.515 117.110 2.680 ;
        RECT 117.950 1.515 120.330 2.680 ;
        RECT 121.170 1.515 123.550 2.680 ;
        RECT 124.390 1.515 127.230 2.680 ;
        RECT 128.070 1.515 130.450 2.680 ;
        RECT 131.290 1.515 134.130 2.680 ;
        RECT 134.970 1.515 137.350 2.680 ;
      LAYER met3 ;
        RECT 1.445 137.680 137.200 138.545 ;
        RECT 1.445 135.680 137.935 137.680 ;
        RECT 1.445 134.280 137.200 135.680 ;
        RECT 1.445 132.280 137.935 134.280 ;
        RECT 1.445 130.880 137.200 132.280 ;
        RECT 1.445 128.880 137.935 130.880 ;
        RECT 1.445 127.480 137.200 128.880 ;
        RECT 1.445 125.480 137.935 127.480 ;
        RECT 1.445 124.080 137.200 125.480 ;
        RECT 1.445 122.080 137.935 124.080 ;
        RECT 1.445 120.680 137.200 122.080 ;
        RECT 1.445 118.680 137.935 120.680 ;
        RECT 1.445 117.280 137.200 118.680 ;
        RECT 1.445 115.280 137.935 117.280 ;
        RECT 1.445 113.880 137.200 115.280 ;
        RECT 1.445 111.880 137.935 113.880 ;
        RECT 1.445 110.480 137.200 111.880 ;
        RECT 1.445 108.480 137.935 110.480 ;
        RECT 1.445 107.080 137.200 108.480 ;
        RECT 1.445 105.760 137.935 107.080 ;
        RECT 1.445 104.360 137.200 105.760 ;
        RECT 1.445 102.360 137.935 104.360 ;
        RECT 1.445 100.960 137.200 102.360 ;
        RECT 1.445 98.960 137.935 100.960 ;
        RECT 1.445 97.560 137.200 98.960 ;
        RECT 1.445 95.560 137.935 97.560 ;
        RECT 1.445 94.160 137.200 95.560 ;
        RECT 1.445 92.160 137.935 94.160 ;
        RECT 1.445 90.760 137.200 92.160 ;
        RECT 1.445 88.760 137.935 90.760 ;
        RECT 1.445 87.360 137.200 88.760 ;
        RECT 1.445 85.360 137.935 87.360 ;
        RECT 1.445 83.960 137.200 85.360 ;
        RECT 1.445 81.960 137.935 83.960 ;
        RECT 1.445 80.560 137.200 81.960 ;
        RECT 1.445 78.560 137.935 80.560 ;
        RECT 1.445 77.160 137.200 78.560 ;
        RECT 1.445 75.160 137.935 77.160 ;
        RECT 1.445 73.760 137.200 75.160 ;
        RECT 1.445 72.440 137.935 73.760 ;
        RECT 1.445 71.080 137.200 72.440 ;
        RECT 2.800 71.040 137.200 71.080 ;
        RECT 2.800 69.680 137.935 71.040 ;
        RECT 1.445 69.040 137.935 69.680 ;
        RECT 1.445 67.640 137.200 69.040 ;
        RECT 1.445 65.640 137.935 67.640 ;
        RECT 1.445 64.240 137.200 65.640 ;
        RECT 1.445 62.240 137.935 64.240 ;
        RECT 1.445 60.840 137.200 62.240 ;
        RECT 1.445 58.840 137.935 60.840 ;
        RECT 1.445 57.440 137.200 58.840 ;
        RECT 1.445 55.440 137.935 57.440 ;
        RECT 1.445 54.040 137.200 55.440 ;
        RECT 1.445 52.040 137.935 54.040 ;
        RECT 1.445 50.640 137.200 52.040 ;
        RECT 1.445 48.640 137.935 50.640 ;
        RECT 1.445 47.240 137.200 48.640 ;
        RECT 1.445 45.240 137.935 47.240 ;
        RECT 1.445 43.840 137.200 45.240 ;
        RECT 1.445 41.840 137.935 43.840 ;
        RECT 1.445 40.440 137.200 41.840 ;
        RECT 1.445 38.440 137.935 40.440 ;
        RECT 1.445 37.040 137.200 38.440 ;
        RECT 1.445 35.720 137.935 37.040 ;
        RECT 1.445 34.320 137.200 35.720 ;
        RECT 1.445 32.320 137.935 34.320 ;
        RECT 1.445 30.920 137.200 32.320 ;
        RECT 1.445 28.920 137.935 30.920 ;
        RECT 1.445 27.520 137.200 28.920 ;
        RECT 1.445 25.520 137.935 27.520 ;
        RECT 1.445 24.120 137.200 25.520 ;
        RECT 1.445 22.120 137.935 24.120 ;
        RECT 1.445 20.720 137.200 22.120 ;
        RECT 1.445 18.720 137.935 20.720 ;
        RECT 1.445 17.320 137.200 18.720 ;
        RECT 1.445 15.320 137.935 17.320 ;
        RECT 1.445 13.920 137.200 15.320 ;
        RECT 1.445 11.920 137.935 13.920 ;
        RECT 1.445 10.520 137.200 11.920 ;
        RECT 1.445 8.520 137.935 10.520 ;
        RECT 1.445 7.120 137.200 8.520 ;
        RECT 1.445 5.120 137.935 7.120 ;
        RECT 1.445 3.720 137.200 5.120 ;
        RECT 1.445 2.400 137.935 3.720 ;
        RECT 1.445 1.535 137.200 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 123.905 128.080 ;
  END
END sb_0__2_
END LIBRARY

