VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_0__1_
  CLASS BLOCK ;
  FOREIGN cby_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 85.000 BY 100.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 96.000 1.290 100.000 ;
    END
  END IO_ISOL_N
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 61.920 85.000 62.520 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 96.000 44.530 100.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 96.000 65.230 100.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 96.000 67.530 100.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.090 96.000 69.370 100.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 96.000 71.670 100.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 96.000 73.510 100.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 96.000 75.810 100.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 96.000 77.650 100.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 96.000 79.950 100.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 96.000 81.790 100.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.810 96.000 84.090 100.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 96.000 46.830 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 96.000 50.970 100.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 96.000 52.810 100.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 96.000 56.950 100.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 96.000 59.250 100.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 96.000 61.090 100.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.110 96.000 63.390 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 96.000 3.130 100.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.550 96.000 23.830 100.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 96.000 26.130 100.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 96.000 27.970 100.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 96.000 30.270 100.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.830 96.000 32.110 100.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 96.000 34.410 100.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 96.000 36.250 100.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 96.000 38.550 100.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.110 96.000 40.390 100.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 96.000 42.690 100.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 96.000 5.430 100.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.990 96.000 7.270 100.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 96.000 9.570 100.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.130 96.000 11.410 100.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.430 96.000 13.710 100.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 96.000 15.550 100.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 96.000 17.850 100.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 21.710 96.000 21.990 100.000 ;
    END
  END chany_top_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN left_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END left_grid_pin_0_
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 81.000 36.760 85.000 37.360 ;
    END
  END prog_clk_0_E_in
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 12.280 85.000 12.880 ;
    END
  END right_width_0_height_0__pin_1_lower
  PIN right_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 81.000 87.080 85.000 87.680 ;
    END
  END right_width_0_height_0__pin_1_upper
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.045 10.640 18.645 87.280 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.375 10.640 30.975 87.280 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 79.120 87.125 ;
      LAYER met1 ;
        RECT 0.990 9.560 84.110 87.280 ;
      LAYER met2 ;
        RECT 1.570 95.720 2.570 96.000 ;
        RECT 3.410 95.720 4.870 96.000 ;
        RECT 5.710 95.720 6.710 96.000 ;
        RECT 7.550 95.720 9.010 96.000 ;
        RECT 9.850 95.720 10.850 96.000 ;
        RECT 11.690 95.720 13.150 96.000 ;
        RECT 13.990 95.720 14.990 96.000 ;
        RECT 15.830 95.720 17.290 96.000 ;
        RECT 18.130 95.720 19.130 96.000 ;
        RECT 19.970 95.720 21.430 96.000 ;
        RECT 22.270 95.720 23.270 96.000 ;
        RECT 24.110 95.720 25.570 96.000 ;
        RECT 26.410 95.720 27.410 96.000 ;
        RECT 28.250 95.720 29.710 96.000 ;
        RECT 30.550 95.720 31.550 96.000 ;
        RECT 32.390 95.720 33.850 96.000 ;
        RECT 34.690 95.720 35.690 96.000 ;
        RECT 36.530 95.720 37.990 96.000 ;
        RECT 38.830 95.720 39.830 96.000 ;
        RECT 40.670 95.720 42.130 96.000 ;
        RECT 42.970 95.720 43.970 96.000 ;
        RECT 44.810 95.720 46.270 96.000 ;
        RECT 47.110 95.720 48.110 96.000 ;
        RECT 48.950 95.720 50.410 96.000 ;
        RECT 51.250 95.720 52.250 96.000 ;
        RECT 53.090 95.720 54.550 96.000 ;
        RECT 55.390 95.720 56.390 96.000 ;
        RECT 57.230 95.720 58.690 96.000 ;
        RECT 59.530 95.720 60.530 96.000 ;
        RECT 61.370 95.720 62.830 96.000 ;
        RECT 63.670 95.720 64.670 96.000 ;
        RECT 65.510 95.720 66.970 96.000 ;
        RECT 67.810 95.720 68.810 96.000 ;
        RECT 69.650 95.720 71.110 96.000 ;
        RECT 71.950 95.720 72.950 96.000 ;
        RECT 73.790 95.720 75.250 96.000 ;
        RECT 76.090 95.720 77.090 96.000 ;
        RECT 77.930 95.720 79.390 96.000 ;
        RECT 80.230 95.720 81.230 96.000 ;
        RECT 82.070 95.720 83.530 96.000 ;
        RECT 1.020 4.280 84.080 95.720 ;
        RECT 1.570 4.000 2.570 4.280 ;
        RECT 3.410 4.000 4.870 4.280 ;
        RECT 5.710 4.000 6.710 4.280 ;
        RECT 7.550 4.000 9.010 4.280 ;
        RECT 9.850 4.000 11.310 4.280 ;
        RECT 12.150 4.000 13.150 4.280 ;
        RECT 13.990 4.000 15.450 4.280 ;
        RECT 16.290 4.000 17.750 4.280 ;
        RECT 18.590 4.000 19.590 4.280 ;
        RECT 20.430 4.000 21.890 4.280 ;
        RECT 22.730 4.000 23.730 4.280 ;
        RECT 24.570 4.000 26.030 4.280 ;
        RECT 26.870 4.000 28.330 4.280 ;
        RECT 29.170 4.000 30.170 4.280 ;
        RECT 31.010 4.000 32.470 4.280 ;
        RECT 33.310 4.000 34.770 4.280 ;
        RECT 35.610 4.000 36.610 4.280 ;
        RECT 37.450 4.000 38.910 4.280 ;
        RECT 39.750 4.000 40.750 4.280 ;
        RECT 41.590 4.000 43.050 4.280 ;
        RECT 43.890 4.000 45.350 4.280 ;
        RECT 46.190 4.000 47.190 4.280 ;
        RECT 48.030 4.000 49.490 4.280 ;
        RECT 50.330 4.000 51.790 4.280 ;
        RECT 52.630 4.000 53.630 4.280 ;
        RECT 54.470 4.000 55.930 4.280 ;
        RECT 56.770 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.070 4.280 ;
        RECT 60.910 4.000 62.370 4.280 ;
        RECT 63.210 4.000 64.210 4.280 ;
        RECT 65.050 4.000 66.510 4.280 ;
        RECT 67.350 4.000 68.810 4.280 ;
        RECT 69.650 4.000 70.650 4.280 ;
        RECT 71.490 4.000 72.950 4.280 ;
        RECT 73.790 4.000 74.790 4.280 ;
        RECT 75.630 4.000 77.090 4.280 ;
        RECT 77.930 4.000 79.390 4.280 ;
        RECT 80.230 4.000 81.230 4.280 ;
        RECT 82.070 4.000 83.530 4.280 ;
      LAYER met3 ;
        RECT 4.400 90.760 81.000 91.625 ;
        RECT 4.000 88.080 81.000 90.760 ;
        RECT 4.000 86.680 80.600 88.080 ;
        RECT 4.000 75.840 81.000 86.680 ;
        RECT 4.400 74.440 81.000 75.840 ;
        RECT 4.000 62.920 81.000 74.440 ;
        RECT 4.000 61.520 80.600 62.920 ;
        RECT 4.000 58.840 81.000 61.520 ;
        RECT 4.400 57.440 81.000 58.840 ;
        RECT 4.000 42.520 81.000 57.440 ;
        RECT 4.400 41.120 81.000 42.520 ;
        RECT 4.000 37.760 81.000 41.120 ;
        RECT 4.000 36.360 80.600 37.760 ;
        RECT 4.000 25.520 81.000 36.360 ;
        RECT 4.400 24.120 81.000 25.520 ;
        RECT 4.000 13.280 81.000 24.120 ;
        RECT 4.000 11.880 80.600 13.280 ;
        RECT 4.000 9.200 81.000 11.880 ;
        RECT 4.400 7.800 81.000 9.200 ;
        RECT 4.000 4.255 81.000 7.800 ;
      LAYER met4 ;
        RECT 31.375 10.640 67.950 87.280 ;
  END
END cby_0__1_
END LIBRARY

