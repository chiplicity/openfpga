VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 137.600 3.590 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 3.440 140.000 4.040 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.920 140.000 11.520 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 137.600 17.390 140.000 ;
    END
  END address[6]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.040 140.000 34.640 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 42.200 140.000 42.800 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.680 140.000 50.280 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 137.600 31.190 140.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 137.600 52.350 140.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 57.840 140.000 58.440 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.320 140.000 65.920 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 137.600 73.510 140.000 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 73.480 140.000 74.080 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 88.440 140.000 89.040 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 96.600 140.000 97.200 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 137.600 101.110 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.080 140.000 104.680 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 119.720 140.000 120.320 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 137.600 108.470 140.000 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.400 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.400 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.400 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 127.880 140.000 128.480 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 137.600 122.270 140.000 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 137.600 129.170 140.000 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 0.040 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.100 137.320 3.030 137.770 ;
        RECT 3.870 137.320 9.930 137.770 ;
        RECT 10.770 137.320 16.830 137.770 ;
        RECT 17.670 137.320 23.730 137.770 ;
        RECT 24.570 137.320 30.630 137.770 ;
        RECT 31.470 137.320 37.990 137.770 ;
        RECT 38.830 137.320 44.890 137.770 ;
        RECT 45.730 137.320 51.790 137.770 ;
        RECT 52.630 137.320 58.690 137.770 ;
        RECT 59.530 137.320 65.590 137.770 ;
        RECT 66.430 137.320 72.950 137.770 ;
        RECT 73.790 137.320 79.850 137.770 ;
        RECT 80.690 137.320 86.750 137.770 ;
        RECT 87.590 137.320 93.650 137.770 ;
        RECT 94.490 137.320 100.550 137.770 ;
        RECT 101.390 137.320 107.910 137.770 ;
        RECT 108.750 137.320 114.810 137.770 ;
        RECT 115.650 137.320 121.710 137.770 ;
        RECT 122.550 137.320 128.610 137.770 ;
        RECT 129.450 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.370 137.770 ;
        RECT 0.100 2.680 138.370 137.320 ;
        RECT 0.100 0.010 2.110 2.680 ;
        RECT 2.950 0.010 6.710 2.680 ;
        RECT 7.550 0.010 11.310 2.680 ;
        RECT 12.150 0.010 16.370 2.680 ;
        RECT 17.210 0.010 20.970 2.680 ;
        RECT 21.810 0.010 26.030 2.680 ;
        RECT 26.870 0.010 30.630 2.680 ;
        RECT 31.470 0.010 35.690 2.680 ;
        RECT 36.530 0.010 40.290 2.680 ;
        RECT 41.130 0.010 45.350 2.680 ;
        RECT 46.190 0.010 49.950 2.680 ;
        RECT 50.790 0.010 55.010 2.680 ;
        RECT 55.850 0.010 59.610 2.680 ;
        RECT 60.450 0.010 64.670 2.680 ;
        RECT 65.510 0.010 69.270 2.680 ;
        RECT 70.110 0.010 74.330 2.680 ;
        RECT 75.170 0.010 78.930 2.680 ;
        RECT 79.770 0.010 83.990 2.680 ;
        RECT 84.830 0.010 88.590 2.680 ;
        RECT 89.430 0.010 93.650 2.680 ;
        RECT 94.490 0.010 98.250 2.680 ;
        RECT 99.090 0.010 103.310 2.680 ;
        RECT 104.150 0.010 107.910 2.680 ;
        RECT 108.750 0.010 112.970 2.680 ;
        RECT 113.810 0.010 117.570 2.680 ;
        RECT 118.410 0.010 122.630 2.680 ;
        RECT 123.470 0.010 127.230 2.680 ;
        RECT 128.070 0.010 132.290 2.680 ;
        RECT 133.130 0.010 136.890 2.680 ;
        RECT 137.730 0.010 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 134.960 137.200 135.360 ;
        RECT 0.310 128.880 138.650 134.960 ;
        RECT 0.310 127.520 137.200 128.880 ;
        RECT 2.800 127.480 137.200 127.520 ;
        RECT 2.800 126.120 138.650 127.480 ;
        RECT 0.310 120.720 138.650 126.120 ;
        RECT 0.310 119.320 137.200 120.720 ;
        RECT 0.310 118.680 138.650 119.320 ;
        RECT 2.800 117.280 138.650 118.680 ;
        RECT 0.310 113.240 138.650 117.280 ;
        RECT 0.310 111.840 137.200 113.240 ;
        RECT 0.310 109.840 138.650 111.840 ;
        RECT 2.800 108.440 138.650 109.840 ;
        RECT 0.310 105.080 138.650 108.440 ;
        RECT 0.310 103.680 137.200 105.080 ;
        RECT 0.310 101.000 138.650 103.680 ;
        RECT 2.800 99.600 138.650 101.000 ;
        RECT 0.310 97.600 138.650 99.600 ;
        RECT 0.310 96.200 137.200 97.600 ;
        RECT 0.310 92.160 138.650 96.200 ;
        RECT 2.800 90.760 138.650 92.160 ;
        RECT 0.310 89.440 138.650 90.760 ;
        RECT 0.310 88.040 137.200 89.440 ;
        RECT 0.310 83.320 138.650 88.040 ;
        RECT 2.800 81.960 138.650 83.320 ;
        RECT 2.800 81.920 137.200 81.960 ;
        RECT 0.310 80.560 137.200 81.920 ;
        RECT 0.310 75.160 138.650 80.560 ;
        RECT 2.800 74.480 138.650 75.160 ;
        RECT 2.800 73.760 137.200 74.480 ;
        RECT 0.310 73.080 137.200 73.760 ;
        RECT 0.310 66.320 138.650 73.080 ;
        RECT 2.800 64.920 137.200 66.320 ;
        RECT 0.310 58.840 138.650 64.920 ;
        RECT 0.310 57.480 137.200 58.840 ;
        RECT 2.800 57.440 137.200 57.480 ;
        RECT 2.800 56.080 138.650 57.440 ;
        RECT 0.310 50.680 138.650 56.080 ;
        RECT 0.310 49.280 137.200 50.680 ;
        RECT 0.310 48.640 138.650 49.280 ;
        RECT 2.800 47.240 138.650 48.640 ;
        RECT 0.310 43.200 138.650 47.240 ;
        RECT 0.310 41.800 137.200 43.200 ;
        RECT 0.310 39.800 138.650 41.800 ;
        RECT 2.800 38.400 138.650 39.800 ;
        RECT 0.310 35.040 138.650 38.400 ;
        RECT 0.310 33.640 137.200 35.040 ;
        RECT 0.310 30.960 138.650 33.640 ;
        RECT 2.800 29.560 138.650 30.960 ;
        RECT 0.310 27.560 138.650 29.560 ;
        RECT 0.310 26.160 137.200 27.560 ;
        RECT 0.310 22.120 138.650 26.160 ;
        RECT 2.800 20.720 138.650 22.120 ;
        RECT 0.310 19.400 138.650 20.720 ;
        RECT 0.310 18.000 137.200 19.400 ;
        RECT 0.310 13.280 138.650 18.000 ;
        RECT 2.800 11.920 138.650 13.280 ;
        RECT 2.800 11.880 137.200 11.920 ;
        RECT 0.310 10.520 137.200 11.880 ;
        RECT 0.310 5.120 138.650 10.520 ;
        RECT 2.800 4.440 138.650 5.120 ;
        RECT 2.800 3.720 137.200 4.440 ;
        RECT 0.310 3.040 137.200 3.720 ;
        RECT 0.310 0.175 138.650 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.240 27.655 128.080 ;
        RECT 30.055 10.240 50.985 128.080 ;
        RECT 53.385 10.240 138.625 128.080 ;
        RECT 0.295 0.175 138.625 10.240 ;
  END
END sb_1__0_
END LIBRARY

